
module oc8051_gm_top(clk, rst, word_in, xram_data_in, p0_in, p1_in, p2_in, p3_in, property_invalid_rom_pc, property_invalid_dec_rom_pc, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp, property_invalid_xram_addr, property_invalid_xram_data_out);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire [7:0] _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire [7:0] _35795_;
  wire _35796_;
  wire [7:0] _35797_;
  wire _35798_;
  wire [7:0] _35799_;
  wire _35800_;
  wire [7:0] _35801_;
  wire _35802_;
  wire [7:0] _35803_;
  wire _35804_;
  wire [7:0] _35805_;
  wire _35806_;
  wire [7:0] _35807_;
  wire _35808_;
  wire [7:0] _35809_;
  wire _35810_;
  wire [7:0] _35811_;
  wire _35812_;
  wire [7:0] _35813_;
  wire _35814_;
  wire [7:0] _35815_;
  wire _35816_;
  wire [7:0] _35817_;
  wire _35818_;
  wire [7:0] _35819_;
  wire _35820_;
  wire [7:0] _35821_;
  wire _35822_;
  wire [7:0] _35823_;
  wire _35824_;
  wire [7:0] _35825_;
  wire _35826_;
  wire [7:0] _35827_;
  wire [7:0] _35828_;
  wire [7:0] _35829_;
  wire [7:0] _35830_;
  wire [7:0] _35831_;
  wire [7:0] _35832_;
  wire [7:0] _35833_;
  wire [7:0] _35834_;
  wire [7:0] _35835_;
  wire [7:0] _35836_;
  wire [7:0] _35837_;
  wire [7:0] _35838_;
  wire [7:0] _35839_;
  wire [7:0] _35840_;
  wire [7:0] _35841_;
  wire [15:0] _35842_;
  wire [7:0] _35843_;
  wire [7:0] _35844_;
  wire [7:0] _35845_;
  wire [7:0] _35846_;
  wire [7:0] _35847_;
  wire [7:0] _35848_;
  wire [7:0] _35849_;
  wire [7:0] _35850_;
  wire [7:0] _35851_;
  wire [7:0] _35852_;
  wire [15:0] _35853_;
  wire [7:0] _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire [7:0] _35983_;
  wire [7:0] _35984_;
  wire [7:0] _35985_;
  wire [2:0] _35986_;
  wire [2:0] _35987_;
  wire [1:0] _35988_;
  wire [7:0] _35989_;
  wire _35990_;
  wire [1:0] _35991_;
  wire [1:0] _35992_;
  wire [2:0] _35993_;
  wire [2:0] _35994_;
  wire [1:0] _35995_;
  wire [3:0] _35996_;
  wire [1:0] _35997_;
  wire _35998_;
  wire _35999_;
  wire [15:0] _36000_;
  wire [15:0] _36001_;
  wire _36002_;
  wire _36003_;
  wire [4:0] _36004_;
  wire [7:0] _36005_;
  wire [7:0] _36006_;
  wire [7:0] _36007_;
  wire _36008_;
  wire _36009_;
  wire [7:0] _36010_;
  wire [15:0] _36011_;
  wire [15:0] _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire [7:0] _36016_;
  wire [2:0] _36017_;
  wire [7:0] _36018_;
  wire [7:0] _36019_;
  wire _36020_;
  wire [7:0] _36021_;
  wire _36022_;
  wire _36023_;
  wire [3:0] _36024_;
  wire [31:0] _36025_;
  wire [31:0] _36026_;
  wire [7:0] _36027_;
  wire _36028_;
  wire _36029_;
  wire [15:0] _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire [15:0] _36034_;
  wire _36035_;
  wire _36036_;
  wire [7:0] _36037_;
  wire _36038_;
  wire [2:0] _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire [7:0] _36134_;
  wire _36135_;
  wire _36136_;
  wire [7:0] _36137_;
  wire _36138_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IE_gm_next;
  wire [7:0] IP_gm;
  wire [7:0] IP_gm_next;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PCON_gm_next;
  wire [15:0] PC_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SBUF_gm_next;
  wire [7:0] SCON_gm;
  wire [7:0] SCON_gm_next;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TCON_gm_next;
  wire [7:0] TH0_gm;
  wire [7:0] TH0_gm_next;
  wire [7:0] TH1_gm;
  wire [7:0] TH1_gm_next;
  wire [7:0] TL0_gm;
  wire [7:0] TL0_gm_next;
  wire [7:0] TL1_gm;
  wire [7:0] TL1_gm_next;
  wire [7:0] TMOD_gm;
  wire [7:0] TMOD_gm_next;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e0 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e2 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e3 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IE_next ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IP_next ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [7:0] \oc8051_golden_model_1.PCON_next ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SBUF_next ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SCON_next ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TCON_next ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH0_next ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TH1_next ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL0_next ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TL1_next ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire [7:0] \oc8051_golden_model_1.TMOD_next ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_e0 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_e2 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_e3 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_f0 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_f2 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_f3 ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_IN ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_f0 ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_f2 ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_f3 ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [6:0] \oc8051_golden_model_1.n1002 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire \oc8051_golden_model_1.n1004 ;
  wire \oc8051_golden_model_1.n1005 ;
  wire \oc8051_golden_model_1.n1006 ;
  wire \oc8051_golden_model_1.n1007 ;
  wire \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire [7:0] \oc8051_golden_model_1.n1018 ;
  wire [7:0] \oc8051_golden_model_1.n1025 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1028 ;
  wire \oc8051_golden_model_1.n1029 ;
  wire \oc8051_golden_model_1.n1030 ;
  wire \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1040 ;
  wire [7:0] \oc8051_golden_model_1.n1041 ;
  wire \oc8051_golden_model_1.n1057 ;
  wire [7:0] \oc8051_golden_model_1.n1058 ;
  wire [3:0] \oc8051_golden_model_1.n1139 ;
  wire [3:0] \oc8051_golden_model_1.n1141 ;
  wire [3:0] \oc8051_golden_model_1.n1143 ;
  wire [3:0] \oc8051_golden_model_1.n1144 ;
  wire [3:0] \oc8051_golden_model_1.n1145 ;
  wire [3:0] \oc8051_golden_model_1.n1146 ;
  wire [3:0] \oc8051_golden_model_1.n1147 ;
  wire [3:0] \oc8051_golden_model_1.n1148 ;
  wire [3:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1195 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire [8:0] \oc8051_golden_model_1.n1239 ;
  wire [7:0] \oc8051_golden_model_1.n1240 ;
  wire \oc8051_golden_model_1.n1241 ;
  wire [2:0] \oc8051_golden_model_1.n1242 ;
  wire \oc8051_golden_model_1.n1243 ;
  wire [1:0] \oc8051_golden_model_1.n1244 ;
  wire [7:0] \oc8051_golden_model_1.n1245 ;
  wire [6:0] \oc8051_golden_model_1.n1246 ;
  wire \oc8051_golden_model_1.n1247 ;
  wire \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1251 ;
  wire \oc8051_golden_model_1.n1252 ;
  wire \oc8051_golden_model_1.n1253 ;
  wire \oc8051_golden_model_1.n1254 ;
  wire \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1278 ;
  wire [7:0] \oc8051_golden_model_1.n1279 ;
  wire [15:0] \oc8051_golden_model_1.n1310 ;
  wire [7:0] \oc8051_golden_model_1.n1312 ;
  wire \oc8051_golden_model_1.n1313 ;
  wire \oc8051_golden_model_1.n1314 ;
  wire \oc8051_golden_model_1.n1315 ;
  wire \oc8051_golden_model_1.n1316 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire \oc8051_golden_model_1.n1318 ;
  wire \oc8051_golden_model_1.n1319 ;
  wire \oc8051_golden_model_1.n1320 ;
  wire \oc8051_golden_model_1.n1327 ;
  wire [7:0] \oc8051_golden_model_1.n1328 ;
  wire [8:0] \oc8051_golden_model_1.n1330 ;
  wire [8:0] \oc8051_golden_model_1.n1334 ;
  wire \oc8051_golden_model_1.n1335 ;
  wire [3:0] \oc8051_golden_model_1.n1336 ;
  wire [4:0] \oc8051_golden_model_1.n1337 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire [8:0] \oc8051_golden_model_1.n1343 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire [7:0] \oc8051_golden_model_1.n1352 ;
  wire [6:0] \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [7:0] \oc8051_golden_model_1.n1369 ;
  wire [8:0] \oc8051_golden_model_1.n1392 ;
  wire \oc8051_golden_model_1.n1393 ;
  wire [4:0] \oc8051_golden_model_1.n1398 ;
  wire \oc8051_golden_model_1.n1399 ;
  wire \oc8051_golden_model_1.n1407 ;
  wire [7:0] \oc8051_golden_model_1.n1408 ;
  wire [6:0] \oc8051_golden_model_1.n1409 ;
  wire \oc8051_golden_model_1.n1424 ;
  wire [7:0] \oc8051_golden_model_1.n1425 ;
  wire [8:0] \oc8051_golden_model_1.n1427 ;
  wire [8:0] \oc8051_golden_model_1.n1429 ;
  wire \oc8051_golden_model_1.n1430 ;
  wire [3:0] \oc8051_golden_model_1.n1431 ;
  wire [4:0] \oc8051_golden_model_1.n1432 ;
  wire [4:0] \oc8051_golden_model_1.n1434 ;
  wire \oc8051_golden_model_1.n1435 ;
  wire [8:0] \oc8051_golden_model_1.n1436 ;
  wire \oc8051_golden_model_1.n1443 ;
  wire [7:0] \oc8051_golden_model_1.n1444 ;
  wire [6:0] \oc8051_golden_model_1.n1445 ;
  wire \oc8051_golden_model_1.n1460 ;
  wire [7:0] \oc8051_golden_model_1.n1461 ;
  wire [8:0] \oc8051_golden_model_1.n1463 ;
  wire \oc8051_golden_model_1.n1464 ;
  wire \oc8051_golden_model_1.n1471 ;
  wire [7:0] \oc8051_golden_model_1.n1472 ;
  wire [6:0] \oc8051_golden_model_1.n1473 ;
  wire [7:0] \oc8051_golden_model_1.n1474 ;
  wire [8:0] \oc8051_golden_model_1.n1476 ;
  wire [8:0] \oc8051_golden_model_1.n1478 ;
  wire \oc8051_golden_model_1.n1479 ;
  wire [4:0] \oc8051_golden_model_1.n1480 ;
  wire [4:0] \oc8051_golden_model_1.n1482 ;
  wire \oc8051_golden_model_1.n1483 ;
  wire [8:0] \oc8051_golden_model_1.n1484 ;
  wire \oc8051_golden_model_1.n1491 ;
  wire [7:0] \oc8051_golden_model_1.n1492 ;
  wire [6:0] \oc8051_golden_model_1.n1493 ;
  wire \oc8051_golden_model_1.n1508 ;
  wire [7:0] \oc8051_golden_model_1.n1509 ;
  wire [4:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [7:0] \oc8051_golden_model_1.n1513 ;
  wire [6:0] \oc8051_golden_model_1.n1514 ;
  wire [7:0] \oc8051_golden_model_1.n1515 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1518 ;
  wire \oc8051_golden_model_1.n1525 ;
  wire [7:0] \oc8051_golden_model_1.n1526 ;
  wire [6:0] \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [8:0] \oc8051_golden_model_1.n1531 ;
  wire [8:0] \oc8051_golden_model_1.n1532 ;
  wire [7:0] \oc8051_golden_model_1.n1533 ;
  wire [7:0] \oc8051_golden_model_1.n1534 ;
  wire [6:0] \oc8051_golden_model_1.n1535 ;
  wire \oc8051_golden_model_1.n1536 ;
  wire \oc8051_golden_model_1.n1537 ;
  wire \oc8051_golden_model_1.n1538 ;
  wire \oc8051_golden_model_1.n1539 ;
  wire \oc8051_golden_model_1.n1540 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire \oc8051_golden_model_1.n1542 ;
  wire \oc8051_golden_model_1.n1543 ;
  wire \oc8051_golden_model_1.n1550 ;
  wire [7:0] \oc8051_golden_model_1.n1551 ;
  wire [7:0] \oc8051_golden_model_1.n1552 ;
  wire [8:0] \oc8051_golden_model_1.n1555 ;
  wire [8:0] \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [4:0] \oc8051_golden_model_1.n1559 ;
  wire [4:0] \oc8051_golden_model_1.n1561 ;
  wire \oc8051_golden_model_1.n1562 ;
  wire \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1586 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire \oc8051_golden_model_1.n1592 ;
  wire [4:0] \oc8051_golden_model_1.n1594 ;
  wire \oc8051_golden_model_1.n1595 ;
  wire \oc8051_golden_model_1.n1602 ;
  wire [7:0] \oc8051_golden_model_1.n1603 ;
  wire [6:0] \oc8051_golden_model_1.n1604 ;
  wire \oc8051_golden_model_1.n1619 ;
  wire [7:0] \oc8051_golden_model_1.n1620 ;
  wire [8:0] \oc8051_golden_model_1.n1624 ;
  wire \oc8051_golden_model_1.n1625 ;
  wire [4:0] \oc8051_golden_model_1.n1627 ;
  wire \oc8051_golden_model_1.n1628 ;
  wire \oc8051_golden_model_1.n1635 ;
  wire [7:0] \oc8051_golden_model_1.n1636 ;
  wire [6:0] \oc8051_golden_model_1.n1637 ;
  wire \oc8051_golden_model_1.n1652 ;
  wire [7:0] \oc8051_golden_model_1.n1653 ;
  wire [8:0] \oc8051_golden_model_1.n1657 ;
  wire \oc8051_golden_model_1.n1658 ;
  wire [4:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire \oc8051_golden_model_1.n1668 ;
  wire [7:0] \oc8051_golden_model_1.n1669 ;
  wire [6:0] \oc8051_golden_model_1.n1670 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire [7:0] \oc8051_golden_model_1.n1686 ;
  wire [7:0] \oc8051_golden_model_1.n1700 ;
  wire [6:0] \oc8051_golden_model_1.n1701 ;
  wire [7:0] \oc8051_golden_model_1.n1702 ;
  wire \oc8051_golden_model_1.n1746 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire \oc8051_golden_model_1.n1763 ;
  wire [7:0] \oc8051_golden_model_1.n1764 ;
  wire \oc8051_golden_model_1.n1780 ;
  wire [7:0] \oc8051_golden_model_1.n1781 ;
  wire \oc8051_golden_model_1.n1797 ;
  wire [7:0] \oc8051_golden_model_1.n1798 ;
  wire [7:0] \oc8051_golden_model_1.n1810 ;
  wire [6:0] \oc8051_golden_model_1.n1811 ;
  wire [7:0] \oc8051_golden_model_1.n1812 ;
  wire \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1857 ;
  wire \oc8051_golden_model_1.n1873 ;
  wire [7:0] \oc8051_golden_model_1.n1874 ;
  wire \oc8051_golden_model_1.n1890 ;
  wire [7:0] \oc8051_golden_model_1.n1891 ;
  wire \oc8051_golden_model_1.n1907 ;
  wire [7:0] \oc8051_golden_model_1.n1908 ;
  wire \oc8051_golden_model_1.n1983 ;
  wire [7:0] \oc8051_golden_model_1.n1984 ;
  wire \oc8051_golden_model_1.n2000 ;
  wire [7:0] \oc8051_golden_model_1.n2001 ;
  wire \oc8051_golden_model_1.n2017 ;
  wire [7:0] \oc8051_golden_model_1.n2018 ;
  wire \oc8051_golden_model_1.n2034 ;
  wire [7:0] \oc8051_golden_model_1.n2035 ;
  wire \oc8051_golden_model_1.n2039 ;
  wire [6:0] \oc8051_golden_model_1.n2040 ;
  wire [7:0] \oc8051_golden_model_1.n2041 ;
  wire [6:0] \oc8051_golden_model_1.n2042 ;
  wire [7:0] \oc8051_golden_model_1.n2043 ;
  wire \oc8051_golden_model_1.n2058 ;
  wire [7:0] \oc8051_golden_model_1.n2059 ;
  wire \oc8051_golden_model_1.n2087 ;
  wire [7:0] \oc8051_golden_model_1.n2088 ;
  wire [6:0] \oc8051_golden_model_1.n2089 ;
  wire [7:0] \oc8051_golden_model_1.n2090 ;
  wire [3:0] \oc8051_golden_model_1.n2097 ;
  wire \oc8051_golden_model_1.n2098 ;
  wire [7:0] \oc8051_golden_model_1.n2099 ;
  wire [6:0] \oc8051_golden_model_1.n2100 ;
  wire \oc8051_golden_model_1.n2115 ;
  wire [7:0] \oc8051_golden_model_1.n2116 ;
  wire [7:0] \oc8051_golden_model_1.n2273 ;
  wire \oc8051_golden_model_1.n2276 ;
  wire \oc8051_golden_model_1.n2278 ;
  wire \oc8051_golden_model_1.n2284 ;
  wire [7:0] \oc8051_golden_model_1.n2285 ;
  wire [6:0] \oc8051_golden_model_1.n2286 ;
  wire \oc8051_golden_model_1.n2301 ;
  wire [7:0] \oc8051_golden_model_1.n2302 ;
  wire \oc8051_golden_model_1.n2306 ;
  wire \oc8051_golden_model_1.n2308 ;
  wire \oc8051_golden_model_1.n2314 ;
  wire [7:0] \oc8051_golden_model_1.n2315 ;
  wire [6:0] \oc8051_golden_model_1.n2316 ;
  wire \oc8051_golden_model_1.n2331 ;
  wire [7:0] \oc8051_golden_model_1.n2332 ;
  wire \oc8051_golden_model_1.n2336 ;
  wire \oc8051_golden_model_1.n2338 ;
  wire \oc8051_golden_model_1.n2344 ;
  wire [7:0] \oc8051_golden_model_1.n2345 ;
  wire [6:0] \oc8051_golden_model_1.n2346 ;
  wire \oc8051_golden_model_1.n2361 ;
  wire [7:0] \oc8051_golden_model_1.n2362 ;
  wire \oc8051_golden_model_1.n2366 ;
  wire \oc8051_golden_model_1.n2368 ;
  wire \oc8051_golden_model_1.n2374 ;
  wire [7:0] \oc8051_golden_model_1.n2375 ;
  wire [6:0] \oc8051_golden_model_1.n2376 ;
  wire \oc8051_golden_model_1.n2391 ;
  wire [7:0] \oc8051_golden_model_1.n2392 ;
  wire \oc8051_golden_model_1.n2394 ;
  wire [7:0] \oc8051_golden_model_1.n2395 ;
  wire [6:0] \oc8051_golden_model_1.n2396 ;
  wire [7:0] \oc8051_golden_model_1.n2397 ;
  wire [7:0] \oc8051_golden_model_1.n2398 ;
  wire [6:0] \oc8051_golden_model_1.n2399 ;
  wire [7:0] \oc8051_golden_model_1.n2400 ;
  wire [15:0] \oc8051_golden_model_1.n2404 ;
  wire \oc8051_golden_model_1.n2410 ;
  wire [7:0] \oc8051_golden_model_1.n2411 ;
  wire [6:0] \oc8051_golden_model_1.n2412 ;
  wire \oc8051_golden_model_1.n2427 ;
  wire [7:0] \oc8051_golden_model_1.n2428 ;
  wire \oc8051_golden_model_1.n2430 ;
  wire [7:0] \oc8051_golden_model_1.n2431 ;
  wire [6:0] \oc8051_golden_model_1.n2432 ;
  wire [7:0] \oc8051_golden_model_1.n2433 ;
  wire \oc8051_golden_model_1.n2461 ;
  wire [7:0] \oc8051_golden_model_1.n2462 ;
  wire [6:0] \oc8051_golden_model_1.n2463 ;
  wire [7:0] \oc8051_golden_model_1.n2464 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire [6:0] \oc8051_golden_model_1.n2471 ;
  wire [7:0] \oc8051_golden_model_1.n2472 ;
  wire \oc8051_golden_model_1.n2477 ;
  wire [7:0] \oc8051_golden_model_1.n2478 ;
  wire [6:0] \oc8051_golden_model_1.n2479 ;
  wire [7:0] \oc8051_golden_model_1.n2480 ;
  wire \oc8051_golden_model_1.n2485 ;
  wire [7:0] \oc8051_golden_model_1.n2486 ;
  wire [6:0] \oc8051_golden_model_1.n2487 ;
  wire [7:0] \oc8051_golden_model_1.n2488 ;
  wire \oc8051_golden_model_1.n2493 ;
  wire [7:0] \oc8051_golden_model_1.n2494 ;
  wire [6:0] \oc8051_golden_model_1.n2495 ;
  wire [7:0] \oc8051_golden_model_1.n2496 ;
  wire [7:0] \oc8051_golden_model_1.n2517 ;
  wire [6:0] \oc8051_golden_model_1.n2518 ;
  wire [7:0] \oc8051_golden_model_1.n2519 ;
  wire [3:0] \oc8051_golden_model_1.n2520 ;
  wire [7:0] \oc8051_golden_model_1.n2521 ;
  wire \oc8051_golden_model_1.n2522 ;
  wire \oc8051_golden_model_1.n2523 ;
  wire \oc8051_golden_model_1.n2524 ;
  wire \oc8051_golden_model_1.n2525 ;
  wire \oc8051_golden_model_1.n2526 ;
  wire \oc8051_golden_model_1.n2527 ;
  wire \oc8051_golden_model_1.n2528 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire [7:0] \oc8051_golden_model_1.n2537 ;
  wire [7:0] \oc8051_golden_model_1.n2546 ;
  wire [6:0] \oc8051_golden_model_1.n2547 ;
  wire \oc8051_golden_model_1.n2562 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire \oc8051_golden_model_1.n2564 ;
  wire \oc8051_golden_model_1.n2565 ;
  wire \oc8051_golden_model_1.n2566 ;
  wire \oc8051_golden_model_1.n2567 ;
  wire \oc8051_golden_model_1.n2568 ;
  wire \oc8051_golden_model_1.n2569 ;
  wire \oc8051_golden_model_1.n2570 ;
  wire \oc8051_golden_model_1.n2571 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2581 ;
  wire \oc8051_golden_model_1.n2582 ;
  wire \oc8051_golden_model_1.n2583 ;
  wire \oc8051_golden_model_1.n2584 ;
  wire \oc8051_golden_model_1.n2585 ;
  wire \oc8051_golden_model_1.n2586 ;
  wire \oc8051_golden_model_1.n2587 ;
  wire \oc8051_golden_model_1.n2594 ;
  wire [7:0] \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2625 ;
  wire [6:0] \oc8051_golden_model_1.n2626 ;
  wire [7:0] \oc8051_golden_model_1.n2627 ;
  wire \oc8051_golden_model_1.n2646 ;
  wire [7:0] \oc8051_golden_model_1.n2647 ;
  wire [6:0] \oc8051_golden_model_1.n2648 ;
  wire \oc8051_golden_model_1.n2663 ;
  wire [7:0] \oc8051_golden_model_1.n2664 ;
  wire [7:0] \oc8051_golden_model_1.n2668 ;
  wire [3:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2670 ;
  wire \oc8051_golden_model_1.n2671 ;
  wire \oc8051_golden_model_1.n2672 ;
  wire \oc8051_golden_model_1.n2673 ;
  wire \oc8051_golden_model_1.n2674 ;
  wire \oc8051_golden_model_1.n2675 ;
  wire \oc8051_golden_model_1.n2676 ;
  wire \oc8051_golden_model_1.n2677 ;
  wire \oc8051_golden_model_1.n2678 ;
  wire \oc8051_golden_model_1.n2685 ;
  wire [7:0] \oc8051_golden_model_1.n2686 ;
  wire \oc8051_golden_model_1.n2690 ;
  wire \oc8051_golden_model_1.n2691 ;
  wire \oc8051_golden_model_1.n2692 ;
  wire \oc8051_golden_model_1.n2693 ;
  wire \oc8051_golden_model_1.n2694 ;
  wire \oc8051_golden_model_1.n2695 ;
  wire \oc8051_golden_model_1.n2696 ;
  wire \oc8051_golden_model_1.n2697 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire [7:0] \oc8051_golden_model_1.n2705 ;
  wire [15:0] \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2721 ;
  wire [7:0] \oc8051_golden_model_1.n2722 ;
  wire [7:0] \oc8051_golden_model_1.n2723 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire [7:0] \oc8051_golden_model_1.n2740 ;
  wire [7:0] \oc8051_golden_model_1.n2741 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_i ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_i ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire \oc8051_top_1.wbd_ack_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_i ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc_impl;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dec_rom_pc;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  wire property_invalid_psw_1_r;
  output property_invalid_rom_pc;
  output property_invalid_sp;
  wire property_invalid_sp_1_r;
  output property_invalid_xram_addr;
  output property_invalid_xram_data_out;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire wbd_ack_i;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_i;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  wire [15:0] xram_addr_gm;
  input [7:0] xram_data_in;
  wire [7:0] xram_data_in_model;
  wire [7:0] xram_data_in_reg;
  wire [7:0] xram_data_out_gm;
  not (_35796_, rst);
  not (_15249_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_15260_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15271_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15260_);
  and (_15282_, _15271_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_15293_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15260_);
  and (_15304_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _15260_);
  nor (_15314_, _15304_, _15293_);
  and (_15325_, _15314_, _15282_);
  nor (_15336_, _15325_, _15249_);
  and (_15347_, _15249_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15358_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_15369_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _15358_);
  nor (_15380_, _15369_, _15347_);
  not (_15391_, _15380_);
  and (_15401_, _15391_, _15325_);
  or (_15412_, _15401_, _15336_);
  and (_24509_, _15412_, _35796_);
  nor (_15433_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15444_, _15433_);
  and (_15455_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_15466_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_15477_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_15488_, _15477_);
  not (_15498_, _15369_);
  nor (_15509_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_15520_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_15531_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _15520_);
  nor (_15542_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_15553_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_15564_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _15553_);
  nor (_15575_, _15564_, _15542_);
  nor (_15585_, _15575_, _15531_);
  not (_15596_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_15607_, _15531_, _15596_);
  nor (_15618_, _15607_, _15585_);
  and (_15629_, _15618_, _15509_);
  not (_15640_, _15629_);
  and (_15651_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15662_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_15673_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15683_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _15673_);
  and (_15694_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_15705_, _15694_, _15662_);
  and (_15716_, _15705_, _15640_);
  nor (_15727_, _15716_, _15498_);
  not (_15738_, _15347_);
  nor (_15749_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_15760_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _15553_);
  nor (_15770_, _15760_, _15749_);
  nor (_15781_, _15770_, _15531_);
  not (_15792_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_15803_, _15531_, _15792_);
  nor (_15814_, _15803_, _15781_);
  and (_15825_, _15814_, _15509_);
  not (_15836_, _15825_);
  and (_15847_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_15858_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_15868_, _15858_, _15847_);
  and (_15879_, _15868_, _15836_);
  nor (_15890_, _15879_, _15738_);
  nor (_15901_, _15890_, _15727_);
  nor (_15912_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_15923_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _15553_);
  nor (_15934_, _15923_, _15912_);
  nor (_15945_, _15934_, _15531_);
  not (_15955_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_15966_, _15531_, _15955_);
  nor (_15977_, _15966_, _15945_);
  and (_15988_, _15977_, _15509_);
  not (_15999_, _15988_);
  and (_16010_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_16021_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_16032_, _16021_, _16010_);
  and (_16042_, _16032_, _15999_);
  nor (_16053_, _16042_, _15391_);
  nor (_16064_, _16053_, _15433_);
  and (_16075_, _16064_, _15901_);
  nor (_16086_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_16097_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _15553_);
  nor (_16108_, _16097_, _16086_);
  nor (_16119_, _16108_, _15531_);
  not (_16130_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_16140_, _15531_, _16130_);
  nor (_16151_, _16140_, _16119_);
  and (_16162_, _16151_, _15509_);
  not (_16173_, _16162_);
  and (_16184_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_16195_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16206_, _16195_, _16184_);
  and (_16217_, _16206_, _16173_);
  and (_16227_, _16217_, _15433_);
  nor (_16238_, _16227_, _16075_);
  not (_16249_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16260_, _16249_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16271_, _16260_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16282_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_16293_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16304_, _16293_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16314_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_16325_, _16314_, _16282_);
  nor (_16336_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16347_, _16336_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16358_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_16369_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16380_, _16260_, _16369_);
  and (_16391_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_16402_, _16391_, _16358_);
  and (_16412_, _16402_, _16325_);
  and (_16423_, _16336_, _16249_);
  and (_16445_, _16423_, _16151_);
  and (_16446_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16457_, _16446_, _16369_);
  and (_16468_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_16479_, _16446_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16490_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_16500_, _16490_, _16468_);
  not (_16511_, _16500_);
  nor (_16522_, _16511_, _16445_);
  and (_16533_, _16522_, _16412_);
  not (_16544_, _16533_);
  and (_16555_, _16544_, _16238_);
  not (_16566_, _16555_);
  nor (_16577_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_16588_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _15553_);
  nor (_16589_, _16588_, _16577_);
  nor (_16595_, _16589_, _15531_);
  not (_16606_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_16617_, _15531_, _16606_);
  nor (_16628_, _16617_, _16595_);
  and (_16639_, _16628_, _15509_);
  not (_16650_, _16639_);
  and (_16661_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_16672_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_16683_, _16672_, _16661_);
  and (_16693_, _16683_, _16650_);
  nor (_16704_, _16693_, _15498_);
  nor (_16715_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_16726_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _15553_);
  nor (_16737_, _16726_, _16715_);
  nor (_16748_, _16737_, _15531_);
  not (_16759_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_16770_, _15531_, _16759_);
  nor (_16781_, _16770_, _16748_);
  and (_16792_, _16781_, _15509_);
  not (_16803_, _16792_);
  and (_16813_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_16824_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_16835_, _16824_, _16813_);
  and (_16846_, _16835_, _16803_);
  nor (_16857_, _16846_, _15738_);
  nor (_16868_, _16857_, _16704_);
  nor (_16879_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_16890_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _15553_);
  nor (_16901_, _16890_, _16879_);
  nor (_16912_, _16901_, _15531_);
  not (_16922_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_16933_, _15531_, _16922_);
  nor (_16944_, _16933_, _16912_);
  and (_16955_, _16944_, _15509_);
  not (_16966_, _16955_);
  and (_16977_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_16988_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_16999_, _16988_, _16977_);
  and (_17010_, _16999_, _16966_);
  nor (_17021_, _17010_, _15391_);
  nor (_17031_, _17021_, _15433_);
  and (_17042_, _17031_, _16868_);
  nor (_17053_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_17064_, _15553_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_17075_, _17064_, _17053_);
  nor (_17086_, _17075_, _15531_);
  not (_17097_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_17108_, _15531_, _17097_);
  nor (_17119_, _17108_, _17086_);
  and (_17130_, _17119_, _15509_);
  not (_17150_, _17130_);
  and (_17151_, _15651_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_17172_, _15683_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_17173_, _17172_, _17151_);
  and (_17184_, _17173_, _17150_);
  and (_17195_, _17184_, _15433_);
  or (_17206_, _17195_, _17042_);
  and (_17217_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_17228_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_17239_, _17228_, _17217_);
  and (_17249_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_17260_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_17271_, _17260_, _17249_);
  and (_17282_, _17271_, _17239_);
  and (_17293_, _17119_, _16423_);
  and (_17304_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_17315_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_17326_, _17315_, _17304_);
  not (_17337_, _17326_);
  nor (_17348_, _17337_, _17293_);
  and (_17358_, _17348_, _17282_);
  nor (_17369_, _17358_, _17206_);
  and (_17380_, _17369_, _16566_);
  not (_17391_, _17380_);
  and (_17402_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_17413_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_17424_, _17413_, _17402_);
  and (_17435_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_17446_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_17456_, _17446_, _17435_);
  and (_17467_, _17456_, _17424_);
  and (_17478_, _16781_, _16423_);
  and (_17489_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_17500_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17511_, _17500_, _17489_);
  not (_17522_, _17511_);
  nor (_17533_, _17522_, _17478_);
  and (_17544_, _17533_, _17467_);
  nor (_17555_, _17544_, _17206_);
  and (_17565_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_17576_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_17587_, _17576_, _17565_);
  and (_17598_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_17609_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_17620_, _17609_, _17598_);
  and (_17631_, _17620_, _17587_);
  and (_17642_, _16423_, _15814_);
  and (_17653_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_17664_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_17674_, _17664_, _17653_);
  not (_17685_, _17674_);
  nor (_17696_, _17685_, _17642_);
  and (_17707_, _17696_, _17631_);
  not (_17718_, _17707_);
  and (_17729_, _17718_, _16238_);
  and (_17740_, _17555_, _17729_);
  and (_17751_, _16544_, _17740_);
  nor (_17762_, _16555_, _17740_);
  nor (_17773_, _17762_, _17751_);
  and (_17783_, _17773_, _17555_);
  and (_17794_, _17369_, _16555_);
  nor (_17805_, _16533_, _17206_);
  not (_17816_, _17358_);
  and (_17827_, _17816_, _16238_);
  nor (_17838_, _17827_, _17805_);
  nor (_17849_, _17838_, _17794_);
  and (_17860_, _17849_, _17783_);
  nor (_17871_, _17849_, _17783_);
  nor (_17882_, _17871_, _17860_);
  and (_17892_, _17882_, _17751_);
  nor (_17903_, _17892_, _17860_);
  nor (_17914_, _17903_, _17391_);
  nor (_17925_, _17206_, _17707_);
  and (_17936_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_17947_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_17958_, _17947_, _17936_);
  and (_17969_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_17980_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_17990_, _17980_, _17969_);
  and (_18001_, _17990_, _17958_);
  and (_18012_, _16628_, _16423_);
  and (_18023_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_18034_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_18045_, _18034_, _18023_);
  not (_18056_, _18045_);
  nor (_18067_, _18056_, _18012_);
  and (_18078_, _18067_, _18001_);
  not (_18089_, _18078_);
  and (_18099_, _18089_, _16238_);
  and (_18110_, _18099_, _17925_);
  not (_18121_, _17544_);
  and (_18132_, _18121_, _16238_);
  nor (_18143_, _18132_, _17925_);
  nor (_18154_, _18143_, _17740_);
  and (_18165_, _18154_, _18110_);
  nor (_18176_, _16555_, _17555_);
  nor (_18187_, _18176_, _17783_);
  and (_18198_, _18187_, _18165_);
  nor (_18208_, _17882_, _17751_);
  nor (_18219_, _18208_, _17892_);
  and (_18230_, _18219_, _18198_);
  nor (_18241_, _18219_, _18198_);
  nor (_18252_, _18241_, _18230_);
  not (_18263_, _18252_);
  and (_18274_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_18285_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_18296_, _18285_, _18274_);
  and (_18307_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_18317_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_18328_, _18317_, _18307_);
  and (_18339_, _18328_, _18296_);
  and (_18350_, _16944_, _16423_);
  and (_18361_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_18372_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_18383_, _18372_, _18361_);
  not (_18394_, _18383_);
  nor (_18405_, _18394_, _18350_);
  and (_18416_, _18405_, _18339_);
  nor (_18426_, _18416_, _17206_);
  and (_18437_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_18448_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_18459_, _18448_, _18437_);
  and (_18470_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_18481_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  nor (_18492_, _18481_, _18470_);
  and (_18503_, _18492_, _18459_);
  and (_18514_, _16423_, _15618_);
  and (_18524_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_18535_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_18546_, _18535_, _18524_);
  not (_18557_, _18546_);
  nor (_18568_, _18557_, _18514_);
  and (_18579_, _18568_, _18503_);
  not (_18590_, _18579_);
  and (_18601_, _18590_, _16238_);
  and (_18612_, _18601_, _18426_);
  not (_18623_, _18416_);
  and (_18633_, _18623_, _16238_);
  not (_18644_, _18633_);
  nor (_18655_, _18579_, _17206_);
  and (_18666_, _18655_, _18644_);
  and (_18677_, _18666_, _18099_);
  nor (_18688_, _18677_, _18612_);
  nor (_18699_, _18078_, _17206_);
  nor (_18710_, _18699_, _17729_);
  nor (_18721_, _18710_, _18110_);
  not (_18732_, _18721_);
  nor (_18742_, _18732_, _18688_);
  nor (_18753_, _18154_, _18110_);
  nor (_18764_, _18753_, _18165_);
  and (_18775_, _18764_, _18742_);
  nor (_18786_, _18187_, _18165_);
  nor (_18797_, _18786_, _18198_);
  and (_18808_, _18797_, _18775_);
  and (_18819_, _16271_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_18830_, _16304_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_18841_, _18830_, _18819_);
  and (_18851_, _16380_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_18862_, _16347_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_18873_, _18862_, _18851_);
  and (_18884_, _18873_, _18841_);
  and (_18895_, _16423_, _15977_);
  and (_18906_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_18917_, _16479_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_18928_, _18917_, _18906_);
  not (_18939_, _18928_);
  nor (_18949_, _18939_, _18895_);
  and (_18960_, _18949_, _18884_);
  nor (_18971_, _18960_, _17206_);
  and (_18982_, _18971_, _18633_);
  nor (_18993_, _18601_, _18426_);
  nor (_19004_, _18993_, _18612_);
  and (_19015_, _19004_, _18982_);
  nor (_19026_, _18666_, _18099_);
  nor (_19037_, _19026_, _18677_);
  and (_19048_, _19037_, _19015_);
  and (_19058_, _18732_, _18688_);
  nor (_19069_, _19058_, _18742_);
  and (_19080_, _19069_, _19048_);
  nor (_19091_, _18764_, _18742_);
  nor (_19102_, _19091_, _18775_);
  and (_19113_, _19102_, _19080_);
  nor (_19124_, _18797_, _18775_);
  nor (_19135_, _19124_, _18808_);
  and (_19146_, _19135_, _19113_);
  nor (_19157_, _19146_, _18808_);
  nor (_19167_, _19157_, _18263_);
  nor (_19178_, _19167_, _18230_);
  and (_19189_, _17903_, _17391_);
  nor (_19200_, _19189_, _17914_);
  not (_19211_, _19200_);
  nor (_19222_, _19211_, _19178_);
  or (_19233_, _19222_, _17794_);
  nor (_19244_, _19233_, _17914_);
  nor (_19255_, _19244_, _15488_);
  and (_19266_, _19244_, _15488_);
  nor (_19276_, _19266_, _19255_);
  not (_19287_, _19276_);
  and (_19298_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_19309_, _19211_, _19178_);
  nor (_19320_, _19309_, _19222_);
  and (_19331_, _19320_, _19298_);
  and (_19342_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_19353_, _19157_, _18263_);
  nor (_19364_, _19353_, _19167_);
  and (_19375_, _19364_, _19342_);
  nor (_19385_, _19364_, _19342_);
  nor (_19396_, _19385_, _19375_);
  not (_19407_, _19396_);
  and (_19418_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_19429_, _19135_, _19113_);
  nor (_19440_, _19429_, _19146_);
  and (_19451_, _19440_, _19418_);
  nor (_19462_, _19440_, _19418_);
  nor (_19473_, _19462_, _19451_);
  not (_19484_, _19473_);
  and (_19494_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_19505_, _19102_, _19080_);
  nor (_19516_, _19505_, _19113_);
  and (_19527_, _19516_, _19494_);
  nor (_19538_, _19516_, _19494_);
  nor (_19549_, _19538_, _19527_);
  not (_19560_, _19549_);
  and (_19571_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_19582_, _19069_, _19048_);
  nor (_19593_, _19582_, _19080_);
  and (_19603_, _19593_, _19571_);
  and (_19614_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_19625_, _19037_, _19015_);
  nor (_19636_, _19625_, _19048_);
  and (_19647_, _19636_, _19614_);
  and (_19658_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_19669_, _19004_, _18982_);
  nor (_19680_, _19669_, _19015_);
  and (_19691_, _19680_, _19658_);
  nor (_19702_, _19636_, _19614_);
  nor (_19713_, _19702_, _19647_);
  and (_19724_, _19713_, _19691_);
  nor (_19735_, _19724_, _19647_);
  not (_19746_, _19735_);
  nor (_19757_, _19593_, _19571_);
  nor (_19768_, _19757_, _19603_);
  and (_19779_, _19768_, _19746_);
  nor (_19790_, _19779_, _19603_);
  nor (_19801_, _19790_, _19560_);
  nor (_19812_, _19801_, _19527_);
  nor (_19823_, _19812_, _19484_);
  nor (_19834_, _19823_, _19451_);
  nor (_19845_, _19834_, _19407_);
  nor (_19856_, _19845_, _19375_);
  nor (_19867_, _19320_, _19298_);
  nor (_19877_, _19867_, _19331_);
  not (_19888_, _19877_);
  nor (_19899_, _19888_, _19856_);
  nor (_19910_, _19899_, _19331_);
  nor (_19921_, _19910_, _19287_);
  nor (_19932_, _19921_, _19255_);
  not (_19943_, _19932_);
  and (_19954_, _19943_, _15466_);
  and (_19965_, _19954_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_19976_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_19987_, _19976_, _19965_);
  and (_19998_, _19987_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_20009_, _19998_, _15455_);
  and (_20020_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20031_, _20020_, _20009_);
  and (_20042_, _20009_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20053_, _20042_, _20031_);
  and (_26705_, _20053_, _35796_);
  nor (_20074_, _15325_, _15358_);
  and (_20085_, _15325_, _15358_);
  or (_20096_, _20085_, _20074_);
  and (_02556_, _20096_, _35796_);
  not (_20117_, _18960_);
  and (_20128_, _20117_, _16238_);
  and (_02757_, _20128_, _35796_);
  nor (_20149_, _18971_, _18633_);
  nor (_20160_, _20149_, _18982_);
  and (_02961_, _20160_, _35796_);
  nor (_20181_, _19680_, _19658_);
  nor (_20192_, _20181_, _19691_);
  and (_03172_, _20192_, _35796_);
  nor (_20213_, _19713_, _19691_);
  nor (_20224_, _20213_, _19724_);
  and (_03373_, _20224_, _35796_);
  nor (_20245_, _19768_, _19746_);
  nor (_20256_, _20245_, _19779_);
  and (_03574_, _20256_, _35796_);
  and (_20276_, _19790_, _19560_);
  nor (_20287_, _20276_, _19801_);
  and (_03775_, _20287_, _35796_);
  and (_20308_, _19812_, _19484_);
  nor (_20319_, _20308_, _19823_);
  and (_03976_, _20319_, _35796_);
  and (_20340_, _19834_, _19407_);
  nor (_20351_, _20340_, _19845_);
  and (_04177_, _20351_, _35796_);
  and (_20372_, _19888_, _19856_);
  nor (_20383_, _20372_, _19899_);
  and (_04278_, _20383_, _35796_);
  and (_20404_, _19910_, _19287_);
  nor (_20415_, _20404_, _19921_);
  and (_04379_, _20415_, _35796_);
  nor (_20436_, _19943_, _15466_);
  nor (_20447_, _20436_, _19954_);
  and (_04480_, _20447_, _35796_);
  and (_20468_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_20479_, _20468_, _19954_);
  nor (_20490_, _20479_, _19965_);
  and (_04581_, _20490_, _35796_);
  nor (_20511_, _19976_, _19965_);
  nor (_20522_, _20511_, _19987_);
  and (_04682_, _20522_, _35796_);
  and (_20543_, _15444_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_20554_, _20543_, _19987_);
  nor (_20565_, _20554_, _19998_);
  and (_04783_, _20565_, _35796_);
  nor (_20586_, _19998_, _15455_);
  nor (_20597_, _20586_, _20009_);
  and (_04884_, _20597_, _35796_);
  and (_20618_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15260_);
  nor (_20629_, _20618_, _15271_);
  not (_20639_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_20650_, _15293_, _20639_);
  and (_20661_, _20650_, _20629_);
  and (_20672_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_20683_, _20672_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20694_, _20672_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20705_, _20694_, _20683_);
  and (_00915_, _20705_, _35796_);
  and (_00945_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _35796_);
  not (_20736_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_20747_, _17010_, _20736_);
  and (_20758_, _16693_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20769_, _20758_, _20747_);
  nor (_20780_, _20769_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20791_, _16846_, _20736_);
  and (_20802_, _17184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_20813_, _20802_, _20791_);
  and (_20824_, _20813_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20835_, _20824_, _20780_);
  nor (_20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20857_, _20846_, _17358_);
  nor (_20868_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_20879_, _20868_, _20857_);
  not (_20890_, _20879_);
  and (_20901_, _16042_, _20736_);
  and (_20912_, _15716_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20923_, _20912_, _20901_);
  nor (_20934_, _20923_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20945_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20956_, _15879_, _20736_);
  and (_20967_, _16217_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20978_, _20967_, _20956_);
  nor (_20989_, _20978_, _20945_);
  nor (_20999_, _20989_, _20934_);
  nor (_21010_, _20999_, _20890_);
  and (_21021_, _20999_, _20890_);
  nor (_21032_, _21021_, _21010_);
  nor (_21043_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_21054_, _20846_, _16533_);
  nor (_21065_, _21054_, _21043_);
  not (_21076_, _21065_);
  nor (_21087_, _17010_, _20736_);
  nor (_21098_, _21087_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21109_, _16693_, _20736_);
  and (_21120_, _16846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21131_, _21120_, _21109_);
  nor (_21142_, _21131_, _20945_);
  nor (_21153_, _21142_, _21098_);
  nor (_21164_, _21153_, _21076_);
  and (_21175_, _21153_, _21076_);
  nor (_21186_, _21175_, _21164_);
  not (_21197_, _21186_);
  and (_21208_, _20846_, _17544_);
  nor (_21219_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor (_21230_, _21219_, _21208_);
  not (_21241_, _21230_);
  nor (_21252_, _16042_, _20736_);
  nor (_21263_, _21252_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21274_, _15716_, _20736_);
  and (_21285_, _15879_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21296_, _21285_, _21274_);
  nor (_21307_, _21296_, _20945_);
  nor (_21318_, _21307_, _21263_);
  nor (_21329_, _21318_, _21241_);
  and (_21340_, _21318_, _21241_);
  and (_21351_, _20769_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21372_, _21351_);
  and (_21384_, _20846_, _17707_);
  nor (_21396_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  nor (_21408_, _21396_, _21384_);
  and (_21420_, _21408_, _21372_);
  and (_21432_, _20923_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21433_, _21432_);
  and (_21444_, _20846_, _18078_);
  nor (_21455_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_21466_, _21455_, _21444_);
  and (_21477_, _21466_, _21433_);
  nor (_21488_, _21466_, _21433_);
  nor (_21499_, _21488_, _21477_);
  not (_21510_, _21499_);
  and (_21521_, _21087_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21532_, _21521_);
  and (_21543_, _20846_, _18579_);
  nor (_21554_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_21565_, _21554_, _21543_);
  and (_21576_, _21565_, _21532_);
  and (_21587_, _21252_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21598_, _21587_);
  nor (_21609_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_21620_, _20846_, _18416_);
  nor (_21631_, _21620_, _21609_);
  nor (_21642_, _21631_, _21598_);
  not (_21653_, _21642_);
  nor (_21664_, _21565_, _21532_);
  nor (_21675_, _21664_, _21576_);
  and (_21686_, _21675_, _21653_);
  nor (_21697_, _21686_, _21576_);
  nor (_21708_, _21697_, _21510_);
  nor (_21719_, _21708_, _21477_);
  nor (_21730_, _21408_, _21372_);
  nor (_21740_, _21730_, _21420_);
  not (_21751_, _21740_);
  nor (_21762_, _21751_, _21719_);
  nor (_21773_, _21762_, _21420_);
  nor (_21784_, _21773_, _21340_);
  nor (_21795_, _21784_, _21329_);
  nor (_21806_, _21795_, _21197_);
  nor (_21817_, _21806_, _21164_);
  not (_21828_, _21817_);
  and (_21839_, _21828_, _21032_);
  or (_21850_, _21839_, _21010_);
  and (_21861_, _17184_, _16217_);
  or (_21872_, _21861_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_21883_, _21131_);
  and (_21894_, _20813_, _21883_);
  nor (_21905_, _21296_, _20978_);
  and (_21916_, _21905_, _21894_);
  or (_21927_, _21916_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21948_, _21927_, _21872_);
  and (_21949_, _21948_, _21850_);
  and (_21960_, _21949_, _20835_);
  nor (_21971_, _21828_, _21032_);
  or (_21982_, _21971_, _21839_);
  and (_21993_, _21982_, _21960_);
  nor (_22004_, _21960_, _20879_);
  nor (_22015_, _22004_, _21993_);
  not (_22026_, _22015_);
  and (_22037_, _22015_, _20835_);
  not (_22048_, _20999_);
  nor (_22059_, _21960_, _21076_);
  and (_22070_, _21795_, _21197_);
  nor (_22081_, _22070_, _21806_);
  and (_22091_, _22081_, _21960_);
  or (_22102_, _22091_, _22059_);
  and (_22113_, _22102_, _22048_);
  nor (_22124_, _22102_, _22048_);
  nor (_22135_, _22124_, _22113_);
  not (_22146_, _22135_);
  not (_22157_, _21153_);
  nor (_22168_, _21960_, _21241_);
  nor (_22179_, _21340_, _21329_);
  nor (_22190_, _22179_, _21773_);
  and (_22212_, _22179_, _21773_);
  or (_22213_, _22212_, _22190_);
  and (_22224_, _22213_, _21960_);
  or (_22235_, _22224_, _22168_);
  and (_22246_, _22235_, _22157_);
  nor (_22257_, _22235_, _22157_);
  not (_22268_, _21318_);
  and (_22279_, _21751_, _21719_);
  or (_22290_, _22279_, _21762_);
  and (_22301_, _22290_, _21960_);
  nor (_22312_, _21960_, _21408_);
  nor (_22323_, _22312_, _22301_);
  and (_22334_, _22323_, _22268_);
  and (_22345_, _21697_, _21510_);
  nor (_22356_, _22345_, _21708_);
  not (_22367_, _22356_);
  and (_22378_, _22367_, _21960_);
  nor (_22389_, _21960_, _21466_);
  nor (_22400_, _22389_, _22378_);
  and (_22411_, _22400_, _21372_);
  nor (_22422_, _22400_, _21372_);
  nor (_22433_, _22422_, _22411_);
  not (_22444_, _22433_);
  nor (_22455_, _21675_, _21653_);
  nor (_22465_, _22455_, _21686_);
  not (_22476_, _22465_);
  and (_22487_, _22476_, _21960_);
  nor (_22498_, _21960_, _21565_);
  nor (_22509_, _22498_, _22487_);
  and (_22520_, _22509_, _21433_);
  and (_22531_, _21960_, _21587_);
  nor (_22542_, _22531_, _21631_);
  and (_22553_, _22531_, _21631_);
  nor (_22564_, _22553_, _22542_);
  and (_22575_, _22564_, _21532_);
  nor (_22586_, _22564_, _21532_);
  nor (_22597_, _22586_, _22575_);
  and (_22608_, _20846_, _18960_);
  nor (_22619_, _20846_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_22630_, _22619_, _22608_);
  nor (_22641_, _22630_, _21598_);
  not (_22652_, _22641_);
  and (_22663_, _22652_, _22597_);
  nor (_22674_, _22663_, _22575_);
  nor (_22685_, _22509_, _21433_);
  nor (_22696_, _22685_, _22520_);
  not (_22707_, _22696_);
  nor (_22718_, _22707_, _22674_);
  nor (_22729_, _22718_, _22520_);
  nor (_22740_, _22729_, _22444_);
  nor (_22751_, _22740_, _22411_);
  nor (_22762_, _22323_, _22268_);
  nor (_22773_, _22762_, _22334_);
  not (_22784_, _22773_);
  nor (_22794_, _22784_, _22751_);
  nor (_22805_, _22794_, _22334_);
  nor (_22816_, _22805_, _22257_);
  nor (_22827_, _22816_, _22246_);
  nor (_22838_, _22827_, _22146_);
  or (_22849_, _22838_, _22113_);
  or (_22860_, _22849_, _22037_);
  and (_22871_, _22860_, _21948_);
  nor (_22892_, _22871_, _22026_);
  and (_22893_, _22037_, _21948_);
  and (_22904_, _22893_, _22849_);
  or (_22925_, _22904_, _22892_);
  and (_00965_, _22925_, _35796_);
  or (_22936_, _22015_, _20835_);
  and (_22957_, _22936_, _22871_);
  and (_02918_, _22957_, _35796_);
  and (_02929_, _21960_, _35796_);
  and (_02950_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _35796_);
  and (_02972_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _35796_);
  and (_02993_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _35796_);
  or (_23018_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23019_, _20672_, rst);
  and (_03004_, _23019_, _23018_);
  and (_23050_, _22957_, _21587_);
  or (_23051_, _23050_, _22630_);
  nand (_23062_, _23050_, _22630_);
  and (_23083_, _23062_, _23051_);
  and (_03015_, _23083_, _35796_);
  nor (_23094_, _22652_, _22597_);
  or (_23105_, _23094_, _22663_);
  nand (_23116_, _23105_, _22957_);
  or (_23126_, _22957_, _22564_);
  and (_23137_, _23126_, _23116_);
  and (_03026_, _23137_, _35796_);
  and (_23158_, _22707_, _22674_);
  or (_23169_, _23158_, _22718_);
  nand (_23180_, _23169_, _22957_);
  or (_23191_, _22957_, _22509_);
  and (_23202_, _23191_, _23180_);
  and (_03037_, _23202_, _35796_);
  and (_23223_, _22729_, _22444_);
  or (_23234_, _23223_, _22740_);
  nand (_23245_, _23234_, _22957_);
  or (_23256_, _22957_, _22400_);
  and (_23267_, _23256_, _23245_);
  and (_03048_, _23267_, _35796_);
  and (_23288_, _22784_, _22751_);
  or (_23299_, _23288_, _22794_);
  nand (_23310_, _23299_, _22957_);
  or (_23321_, _22957_, _22323_);
  and (_23332_, _23321_, _23310_);
  and (_03059_, _23332_, _35796_);
  or (_23353_, _22257_, _22246_);
  and (_23364_, _23353_, _22805_);
  nor (_23375_, _23353_, _22805_);
  or (_23386_, _23375_, _23364_);
  nand (_23397_, _23386_, _22957_);
  or (_23408_, _22957_, _22235_);
  and (_23419_, _23408_, _23397_);
  and (_03070_, _23419_, _35796_);
  and (_23440_, _22827_, _22146_);
  or (_23450_, _23440_, _22838_);
  nand (_23461_, _23450_, _22957_);
  or (_23472_, _22957_, _22102_);
  and (_23483_, _23472_, _23461_);
  and (_03081_, _23483_, _35796_);
  not (_23504_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23515_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15260_);
  and (_23526_, _23515_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_23537_, _23526_, _23504_);
  not (_23548_, _23537_);
  not (_23559_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_23570_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23581_, _23570_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_23592_, _23581_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_23603_, _23592_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_23614_, _23603_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_23625_, _23614_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_23636_, _23625_, _23559_);
  and (_23647_, _23625_, _23559_);
  nor (_23658_, _23647_, _23636_);
  nor (_23669_, _23658_, _23548_);
  not (_23680_, _23669_);
  not (_23691_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23702_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15260_);
  and (_23713_, _23702_, _23504_);
  and (_23724_, _23713_, _23691_);
  and (_23735_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_23746_, _23735_);
  and (_23757_, _23526_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_23767_, _23757_);
  not (_23778_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_23789_, _23515_, _23778_);
  and (_23800_, _23789_, _23504_);
  and (_23811_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_23822_, _23789_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23833_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_23844_, _23833_, _23811_);
  and (_23855_, _23844_, _23767_);
  and (_23866_, _23855_, _23746_);
  and (_23877_, _23866_, _23680_);
  not (_23888_, _23625_);
  nor (_23899_, _23614_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_23910_, _23899_, _23548_);
  and (_23921_, _23910_, _23888_);
  not (_23932_, _23921_);
  and (_23943_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_23954_, _23943_, _23757_);
  and (_23965_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_23976_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_23987_, _23976_, _23965_);
  and (_23998_, _23987_, _23954_);
  and (_24009_, _23998_, _23932_);
  nor (_24020_, _24009_, _23877_);
  and (_24031_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_24042_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_24053_, _24042_, _24031_);
  not (_24074_, _23592_);
  nor (_24086_, _23581_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_24098_, _24086_, _23548_);
  and (_24110_, _24098_, _24074_);
  or (_24122_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24134_, _24122_, _15260_);
  nor (_24146_, _24134_, _23515_);
  and (_24147_, _24146_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_24158_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_24169_, _24158_, _24147_);
  not (_24180_, _24169_);
  nor (_24191_, _24180_, _24110_);
  and (_24202_, _24191_, _24053_);
  not (_24213_, _24202_);
  and (_24224_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_24235_, _24224_);
  and (_24246_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_24257_, _24246_, _23757_);
  and (_24268_, _24257_, _24235_);
  nor (_24279_, _23592_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_24290_, _24279_);
  nor (_24301_, _23603_, _23548_);
  and (_24312_, _24301_, _24290_);
  and (_24323_, _24146_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_24334_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_24345_, _24334_, _24323_);
  not (_24356_, _24345_);
  nor (_24367_, _24356_, _24312_);
  and (_24378_, _24367_, _24268_);
  nor (_24389_, _24378_, _24213_);
  nor (_24399_, _23603_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_24410_, _24399_);
  nor (_24421_, _23614_, _23548_);
  and (_24432_, _24421_, _24410_);
  not (_24443_, _24432_);
  and (_24454_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_24465_, _24454_, _23757_);
  and (_24476_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_24487_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_24498_, _24487_, _24476_);
  and (_24510_, _24498_, _24465_);
  and (_24521_, _24510_, _24443_);
  not (_24532_, _24521_);
  and (_24543_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_24554_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_24565_, _24554_, _24543_);
  and (_24576_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_24587_, _24576_);
  not (_24598_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24609_, _23537_, _24598_);
  and (_24620_, _24146_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24631_, _24620_, _24609_);
  and (_24642_, _24631_, _24587_);
  and (_24653_, _24642_, _24565_);
  nor (_24664_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24675_, _24664_, _23570_);
  and (_24686_, _24675_, _23537_);
  and (_24697_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_24707_, _24697_, _24686_);
  and (_24718_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_24729_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_24740_, _24146_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_24751_, _24740_, _24729_);
  nor (_24762_, _24751_, _24718_);
  and (_24773_, _24762_, _24707_);
  nor (_24784_, _23570_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24795_, _24784_, _23581_);
  and (_24806_, _24795_, _23537_);
  and (_24817_, _23724_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24828_, _24817_, _24806_);
  and (_24839_, _23822_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24850_, _23800_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_24861_, _24146_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24872_, _24861_, _24850_);
  nor (_24883_, _24872_, _24839_);
  and (_24894_, _24883_, _24828_);
  and (_24905_, _24894_, _24773_);
  and (_24916_, _24905_, _24653_);
  and (_24927_, _24916_, _24532_);
  and (_24938_, _24927_, _24389_);
  nand (_24949_, _24938_, _24020_);
  and (_24960_, _22925_, _20661_);
  not (_24971_, _24960_);
  and (_24982_, _20053_, _15325_);
  not (_25003_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_25004_, _20618_, _25003_);
  and (_25015_, _25004_, _15314_);
  nor (_25026_, _16533_, _16217_);
  and (_25047_, _16533_, _16217_);
  nor (_25048_, _25047_, _25026_);
  not (_25059_, _25048_);
  nor (_25080_, _17544_, _16846_);
  and (_25081_, _17544_, _16846_);
  nor (_25092_, _25081_, _25080_);
  nor (_25103_, _17707_, _15879_);
  and (_25114_, _25103_, _25092_);
  nor (_25135_, _25114_, _25080_);
  nor (_25136_, _25135_, _25059_);
  and (_25147_, _17707_, _15879_);
  nor (_25158_, _25147_, _25103_);
  nor (_25169_, _18078_, _16693_);
  and (_25180_, _18078_, _16693_);
  nor (_25191_, _25180_, _25169_);
  nor (_25202_, _18579_, _15716_);
  and (_25213_, _18579_, _15716_);
  nor (_25224_, _25213_, _25202_);
  not (_25235_, _25224_);
  nor (_25246_, _18416_, _17010_);
  nor (_25267_, _18960_, _16042_);
  and (_25268_, _18416_, _17010_);
  nor (_25279_, _25268_, _25246_);
  and (_25290_, _25279_, _25267_);
  nor (_25301_, _25290_, _25246_);
  nor (_25312_, _25301_, _25235_);
  nor (_25323_, _25312_, _25202_);
  nor (_25334_, _25323_, _25191_);
  and (_25345_, _25323_, _25191_);
  nor (_25356_, _25345_, _25334_);
  not (_25367_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_25378_, _15531_, _25367_);
  not (_25389_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_25400_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25411_, _25400_, _17075_);
  nor (_25422_, _25411_, _25389_);
  nor (_25443_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25444_, _25443_, _15770_);
  not (_25455_, _25444_);
  not (_25466_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25477_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25466_);
  and (_25488_, _25477_, _16737_);
  not (_25499_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_25510_, _25499_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25521_, _25510_, _16108_);
  nor (_25532_, _25521_, _25488_);
  and (_25543_, _25532_, _25455_);
  and (_25554_, _25543_, _25422_);
  and (_25565_, _25400_, _16589_);
  nor (_25576_, _25565_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_25587_, _25510_, _15575_);
  not (_25598_, _25587_);
  and (_25609_, _25477_, _16901_);
  and (_25620_, _25443_, _15934_);
  nor (_25641_, _25620_, _25609_);
  and (_25642_, _25641_, _25598_);
  and (_25653_, _25642_, _25576_);
  nor (_25664_, _25653_, _25554_);
  nor (_25675_, _25664_, _15531_);
  nor (_25686_, _25675_, _25378_);
  and (_25697_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_25708_, _25697_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_25719_, _25708_);
  and (_25730_, _25719_, _25686_);
  and (_25741_, _25719_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_25752_, _25741_, _25730_);
  and (_25763_, _18960_, _16042_);
  nor (_25774_, _25763_, _25267_);
  not (_25785_, _25774_);
  nor (_25796_, _25785_, _25752_);
  and (_25807_, _25796_, _25279_);
  and (_25818_, _25301_, _25235_);
  nor (_25829_, _25818_, _25312_);
  and (_25840_, _25829_, _25807_);
  not (_25851_, _25840_);
  nor (_25862_, _25851_, _25356_);
  nor (_25873_, _25323_, _25180_);
  or (_25884_, _25873_, _25169_);
  or (_25895_, _25884_, _25862_);
  and (_25906_, _25895_, _25158_);
  and (_25917_, _25906_, _25092_);
  and (_25928_, _25135_, _25059_);
  nor (_25939_, _25928_, _25136_);
  and (_25950_, _25939_, _25917_);
  or (_25961_, _25950_, _25136_);
  nor (_25972_, _25961_, _25026_);
  nor (_25993_, _17358_, _17184_);
  and (_25994_, _17358_, _17184_);
  nor (_26005_, _25994_, _25993_);
  and (_26016_, _26005_, _25972_);
  nor (_26027_, _26005_, _25972_);
  or (_26038_, _26027_, _26016_);
  and (_26049_, _26038_, _25015_);
  not (_26060_, _26049_);
  not (_26071_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_26082_, _15271_, _26071_);
  and (_26103_, _26082_, _15314_);
  not (_26104_, _26103_);
  not (_26115_, _16217_);
  nor (_26126_, _16533_, _26115_);
  not (_26137_, _16846_);
  nor (_26148_, _17544_, _26137_);
  not (_26159_, _15879_);
  and (_26170_, _17707_, _26159_);
  nor (_26181_, _26170_, _25092_);
  nor (_26192_, _26181_, _26148_);
  nor (_26203_, _26192_, _25048_);
  nor (_26214_, _26203_, _26126_);
  and (_26224_, _26192_, _25048_);
  nor (_26235_, _26224_, _26203_);
  not (_26246_, _26235_);
  and (_26257_, _26170_, _25092_);
  nor (_26268_, _26257_, _26181_);
  not (_26279_, _26268_);
  not (_26290_, _25158_);
  not (_26301_, _16042_);
  and (_26312_, _18960_, _26301_);
  nor (_26323_, _26312_, _25279_);
  not (_26333_, _17010_);
  nor (_26344_, _18416_, _26333_);
  nor (_26355_, _26344_, _26323_);
  nor (_26366_, _26355_, _25224_);
  not (_26377_, _15716_);
  nor (_26388_, _18579_, _26377_);
  nor (_26399_, _26388_, _26366_);
  nor (_26410_, _26399_, _25191_);
  and (_26421_, _26399_, _25191_);
  nor (_26432_, _26421_, _26410_);
  not (_26443_, _26432_);
  and (_26454_, _26355_, _25224_);
  nor (_26465_, _26454_, _26366_);
  not (_26476_, _26465_);
  and (_26487_, _26312_, _25279_);
  nor (_26498_, _26487_, _26323_);
  not (_26509_, _26498_);
  nor (_26520_, _25774_, _25752_);
  and (_26531_, _26520_, _26509_);
  and (_26552_, _26531_, _26476_);
  and (_26553_, _26552_, _26443_);
  not (_26564_, _16693_);
  or (_26574_, _18078_, _26564_);
  and (_26585_, _18078_, _26564_);
  or (_26596_, _26399_, _26585_);
  and (_26607_, _26596_, _26574_);
  or (_26618_, _26607_, _26553_);
  and (_26629_, _26618_, _26290_);
  and (_26640_, _26629_, _26279_);
  and (_26651_, _26640_, _26246_);
  nor (_26662_, _26651_, _26214_);
  nor (_26673_, _26662_, _26005_);
  and (_26683_, _26662_, _26005_);
  nor (_26694_, _26683_, _26673_);
  nor (_26706_, _26694_, _26104_);
  and (_26717_, _15304_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_26728_, _26717_, _26082_);
  nor (_26739_, _18960_, _18416_);
  and (_26750_, _26739_, _18590_);
  and (_26761_, _26750_, _18089_);
  and (_26772_, _26761_, _17718_);
  and (_26783_, _26772_, _18121_);
  and (_26793_, _26783_, _16544_);
  and (_26804_, _26793_, _25752_);
  not (_26815_, _25752_);
  and (_26826_, _16533_, _17544_);
  and (_26847_, _18960_, _18416_);
  and (_26848_, _26847_, _18579_);
  and (_26859_, _26848_, _18078_);
  and (_26870_, _26859_, _17707_);
  and (_26881_, _26870_, _26826_);
  and (_26892_, _26881_, _26815_);
  nor (_26902_, _26892_, _26804_);
  and (_26913_, _26902_, _17358_);
  nor (_26924_, _26902_, _17358_);
  nor (_26935_, _26924_, _26913_);
  and (_26956_, _26935_, _26728_);
  not (_26957_, _17184_);
  nor (_26968_, _25752_, _26957_);
  not (_26979_, _26968_);
  and (_26990_, _25752_, _17358_);
  and (_27001_, _26717_, _15282_);
  not (_27012_, _27001_);
  nor (_27023_, _27012_, _26990_);
  and (_27034_, _27023_, _26979_);
  nor (_27045_, _27034_, _26956_);
  and (_27056_, _25004_, _20650_);
  not (_27067_, _27056_);
  and (_27078_, _18579_, _18416_);
  nor (_27079_, _27078_, _18078_);
  and (_27080_, _27079_, _27056_);
  and (_27089_, _27080_, _17718_);
  nor (_27100_, _27089_, _18121_);
  and (_27111_, _27100_, _16533_);
  nor (_27122_, _26826_, _17358_);
  nor (_27133_, _27122_, _27080_);
  and (_27154_, _27133_, _25752_);
  nor (_27155_, _27154_, _27111_);
  and (_27165_, _27155_, _17358_);
  nor (_27176_, _27155_, _17358_);
  nor (_27187_, _27176_, _27165_);
  nor (_27198_, _27187_, _27067_);
  not (_27209_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27220_, _15304_, _27209_);
  and (_27231_, _27220_, _25004_);
  not (_27242_, _27231_);
  nor (_27253_, _27242_, _25994_);
  and (_27264_, _27220_, _20629_);
  and (_27275_, _27264_, _26005_);
  nor (_27286_, _27275_, _27253_);
  and (_27296_, _26717_, _20629_);
  not (_27307_, _27296_);
  nor (_27318_, _27307_, _18960_);
  and (_27329_, _27220_, _15271_);
  not (_27340_, _27329_);
  nor (_27351_, _27340_, _16533_);
  nor (_27362_, _27351_, _27318_);
  and (_27373_, _26717_, _25004_);
  not (_27384_, _27373_);
  nor (_27395_, _27384_, _25752_);
  and (_27415_, _20650_, _15282_);
  and (_27416_, _27415_, _25993_);
  and (_27427_, _26082_, _20650_);
  and (_27438_, _27427_, _17358_);
  nor (_27449_, _27438_, _27416_);
  and (_27460_, _20629_, _15314_);
  not (_27471_, _27460_);
  nor (_27482_, _27471_, _17358_);
  not (_27493_, _27482_);
  nand (_27504_, _27493_, _27449_);
  nor (_27515_, _27504_, _27395_);
  and (_27526_, _27515_, _27362_);
  and (_27536_, _27526_, _27286_);
  not (_27547_, _27536_);
  nor (_27558_, _27547_, _27198_);
  and (_27569_, _27558_, _27045_);
  not (_27580_, _27569_);
  nor (_27591_, _27580_, _26706_);
  and (_27602_, _27591_, _26060_);
  not (_27613_, _27602_);
  nor (_27624_, _27613_, _24982_);
  and (_27635_, _27624_, _24971_);
  not (_27646_, _27635_);
  or (_27657_, _27646_, _24949_);
  not (_27668_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_27678_, \oc8051_top_1.oc8051_decoder1.wr , _15260_);
  not (_27699_, _27678_);
  nor (_27700_, _27699_, _23713_);
  and (_27711_, _27700_, _27668_);
  not (_27722_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_27733_, _24949_, _27722_);
  and (_27744_, _27733_, _27711_);
  and (_27755_, _27744_, _27657_);
  nor (_27766_, _27700_, _27722_);
  not (_27777_, _25015_);
  nor (_27788_, _25994_, _25972_);
  nor (_27799_, _27788_, _25993_);
  nor (_27809_, _27799_, _27777_);
  not (_27820_, _27809_);
  and (_27831_, _17358_, _26957_);
  nor (_27842_, _27831_, _26673_);
  nor (_27853_, _27842_, _26104_);
  and (_27864_, _25752_, _16533_);
  and (_27875_, _27864_, _27100_);
  nor (_27886_, _27875_, _26990_);
  nor (_27897_, _25752_, _17358_);
  not (_27908_, _27897_);
  nor (_27919_, _27908_, _27111_);
  nor (_27930_, _27919_, _27067_);
  and (_27941_, _27930_, _27886_);
  or (_27945_, _27941_, _27080_);
  nor (_27946_, _25741_, _25686_);
  not (_27947_, _27264_);
  nor (_27948_, _27947_, _25730_);
  not (_27953_, _27948_);
  nor (_27964_, _27307_, _25686_);
  nor (_27975_, _27964_, _27231_);
  and (_27986_, _27975_, _27953_);
  nor (_27997_, _27986_, _27946_);
  not (_28008_, _27997_);
  nor (_28019_, _27471_, _25752_);
  nor (_28030_, _27384_, _18960_);
  and (_28041_, _27220_, _15282_);
  not (_28052_, _28041_);
  nor (_28062_, _28052_, _17358_);
  nor (_28073_, _28062_, _28030_);
  not (_28094_, _28073_);
  nor (_28095_, _28094_, _28019_);
  and (_28105_, _27427_, _25752_);
  and (_28116_, _25708_, _25686_);
  and (_28127_, _27220_, _26082_);
  and (_28137_, _27415_, _25686_);
  nor (_28147_, _28137_, _28127_);
  nor (_28158_, _28147_, _28116_);
  nor (_28169_, _28158_, _28105_);
  and (_28179_, _28169_, _28095_);
  and (_28190_, _28179_, _28008_);
  not (_28201_, _28190_);
  nor (_28211_, _28201_, _27945_);
  not (_28222_, _28211_);
  nor (_28233_, _28222_, _27853_);
  and (_28243_, _28233_, _27820_);
  nor (_28254_, _24521_, _24009_);
  not (_28274_, _23877_);
  and (_28275_, _24389_, _28274_);
  and (_28285_, _28275_, _28254_);
  not (_28296_, _24653_);
  nor (_28306_, _24894_, _24773_);
  and (_28316_, _28306_, _28296_);
  and (_28327_, _28316_, _28285_);
  nand (_28337_, _28327_, _28243_);
  and (_28347_, _27700_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_28358_, _28327_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_28368_, _28358_, _28347_);
  and (_28378_, _28368_, _28337_);
  or (_28388_, _28378_, _27766_);
  or (_28399_, _28388_, _27755_);
  and (_06574_, _28399_, _35796_);
  and (_28419_, _23083_, _20661_);
  not (_28430_, _28419_);
  and (_28440_, _20383_, _15325_);
  and (_28451_, _25785_, _25752_);
  nor (_28461_, _28451_, _25796_);
  nor (_28472_, _26103_, _25015_);
  not (_28483_, _28472_);
  and (_28493_, _28483_, _28461_);
  not (_28503_, _28493_);
  nor (_28514_, _28052_, _25752_);
  not (_28525_, _28514_);
  nor (_28534_, _27947_, _25267_);
  nor (_28542_, _28534_, _27231_);
  or (_28549_, _28542_, _25763_);
  and (_28557_, _27415_, _25267_);
  and (_28565_, _27427_, _18960_);
  nor (_28572_, _28565_, _28557_);
  nor (_28580_, _27012_, _16042_);
  and (_28588_, _26728_, _18960_);
  nor (_28595_, _28588_, _28580_);
  and (_28596_, _26717_, _25003_);
  not (_28597_, _28596_);
  nor (_28600_, _28597_, _18416_);
  not (_28608_, _28600_);
  and (_28617_, _28127_, _17816_);
  nor (_28626_, _27460_, _27056_);
  nor (_28637_, _28626_, _18960_);
  nor (_28648_, _28637_, _28617_);
  and (_28659_, _28648_, _28608_);
  and (_28669_, _28659_, _28595_);
  and (_28680_, _28669_, _28572_);
  and (_28691_, _28680_, _28549_);
  and (_28699_, _28691_, _28525_);
  and (_28706_, _28699_, _28503_);
  not (_28727_, _28706_);
  nor (_28728_, _28727_, _28440_);
  and (_28739_, _28728_, _28430_);
  not (_28750_, _28739_);
  or (_28761_, _28750_, _24949_);
  not (_28772_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_28783_, _24949_, _28772_);
  and (_28794_, _28783_, _27711_);
  and (_28805_, _28794_, _28761_);
  nor (_28816_, _27700_, _28772_);
  not (_28827_, _28243_);
  or (_28838_, _28827_, _24949_);
  and (_28849_, _28783_, _28347_);
  and (_28860_, _28849_, _28838_);
  or (_28871_, _28860_, _28816_);
  or (_28882_, _28871_, _28805_);
  and (_08805_, _28882_, _35796_);
  and (_28903_, _20415_, _15325_);
  not (_28914_, _28903_);
  and (_28925_, _23137_, _20661_);
  nor (_28936_, _27012_, _17010_);
  nor (_28947_, _26847_, _26739_);
  not (_28958_, _28947_);
  nor (_28969_, _28958_, _25752_);
  and (_28980_, _28958_, _25752_);
  nor (_28991_, _28980_, _28969_);
  and (_29002_, _28991_, _26728_);
  nor (_29013_, _29002_, _28936_);
  nor (_29024_, _27471_, _18416_);
  nor (_29035_, _28597_, _18579_);
  nor (_29046_, _27340_, _18960_);
  or (_29057_, _29046_, _29035_);
  nor (_29068_, _29057_, _29024_);
  and (_29079_, _27415_, _25246_);
  and (_29090_, _27427_, _18416_);
  nor (_29101_, _29090_, _29079_);
  and (_29112_, _29101_, _29068_);
  nor (_29122_, _27079_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_29133_, _29122_, _18623_);
  nor (_29144_, _29122_, _18623_);
  nor (_29154_, _29144_, _29133_);
  nor (_29165_, _29154_, _27067_);
  and (_29176_, _27264_, _25279_);
  nor (_29186_, _27242_, _25268_);
  or (_29197_, _29186_, _29176_);
  nor (_29208_, _29197_, _29165_);
  and (_29218_, _29208_, _29112_);
  and (_29229_, _29218_, _29013_);
  nor (_29240_, _25279_, _25267_);
  or (_29251_, _29240_, _25290_);
  and (_29272_, _29251_, _25796_);
  nor (_29273_, _29251_, _25796_);
  or (_29284_, _29273_, _29272_);
  and (_29294_, _29284_, _25015_);
  nor (_29305_, _26520_, _26509_);
  nor (_29316_, _29305_, _26531_);
  nor (_29326_, _29316_, _26104_);
  nor (_29337_, _29326_, _29294_);
  and (_29348_, _29337_, _29229_);
  not (_29358_, _29348_);
  nor (_29369_, _29358_, _28925_);
  and (_29380_, _29369_, _28914_);
  not (_29390_, _29380_);
  or (_29401_, _29390_, _24949_);
  not (_29412_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_29423_, _24949_, _29412_);
  and (_29433_, _29423_, _27711_);
  and (_29444_, _29433_, _29401_);
  nor (_29455_, _27700_, _29412_);
  and (_29466_, _24905_, _28296_);
  and (_29477_, _29466_, _28285_);
  or (_29488_, _29477_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_29499_, _29488_, _28347_);
  nand (_29510_, _29477_, _28243_);
  and (_29531_, _29510_, _29499_);
  or (_29532_, _29531_, _29455_);
  or (_29543_, _29532_, _29444_);
  and (_08816_, _29543_, _35796_);
  and (_29564_, _20447_, _15325_);
  not (_29575_, _29564_);
  and (_29586_, _23202_, _20661_);
  nor (_29597_, _27012_, _15716_);
  nor (_29608_, _26847_, _25752_);
  nor (_29619_, _26739_, _26815_);
  nor (_29630_, _29619_, _29608_);
  and (_29641_, _29630_, _18590_);
  nor (_29652_, _29630_, _18590_);
  nor (_29663_, _29652_, _29641_);
  and (_29674_, _29663_, _26728_);
  nor (_29685_, _29674_, _29597_);
  nor (_29696_, _26531_, _26476_);
  nor (_29707_, _29696_, _26552_);
  nor (_29718_, _29707_, _26104_);
  not (_29729_, _29718_);
  nor (_29740_, _28597_, _18078_);
  and (_29751_, _27415_, _25202_);
  and (_29762_, _27427_, _18579_);
  nor (_29773_, _29762_, _29751_);
  nor (_29784_, _27242_, _25213_);
  and (_29795_, _27264_, _25224_);
  nor (_29806_, _29795_, _29784_);
  nor (_29817_, _27340_, _18416_);
  nor (_29838_, _27471_, _18579_);
  nor (_29839_, _29838_, _29817_);
  and (_29850_, _29839_, _29806_);
  nand (_29861_, _29850_, _29773_);
  nor (_29872_, _29861_, _29740_);
  and (_29883_, _29872_, _29729_);
  nor (_29894_, _25829_, _25807_);
  nor (_29905_, _29894_, _27777_);
  and (_29916_, _29905_, _25851_);
  nor (_29927_, _29144_, _18579_);
  and (_29938_, _27078_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_29949_, _29938_, _29927_);
  nor (_29960_, _29949_, _27067_);
  nor (_29971_, _29960_, _29916_);
  and (_29982_, _29971_, _29883_);
  and (_29992_, _29982_, _29685_);
  not (_30003_, _29992_);
  nor (_30014_, _30003_, _29586_);
  and (_30024_, _30014_, _29575_);
  not (_30035_, _30024_);
  or (_30046_, _30035_, _24949_);
  not (_30056_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_30067_, _24949_, _30056_);
  and (_30078_, _30067_, _27711_);
  and (_30088_, _30078_, _30046_);
  nor (_30099_, _27700_, _30056_);
  nand (_30110_, _28285_, _24894_);
  nor (_30121_, _24773_, _24653_);
  or (_30131_, _30121_, _30110_);
  and (_30142_, _30131_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_30163_, _24773_);
  and (_30164_, _24894_, _30163_);
  and (_30175_, _30164_, _24653_);
  and (_30186_, _30175_, _28827_);
  and (_30192_, _24905_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_30193_, _30192_, _30186_);
  and (_30194_, _30193_, _28285_);
  or (_30195_, _30194_, _30142_);
  and (_30196_, _30195_, _28347_);
  or (_30197_, _30196_, _30099_);
  or (_30198_, _30197_, _30088_);
  and (_08827_, _30198_, _35796_);
  and (_30199_, _23267_, _20661_);
  not (_30200_, _30199_);
  and (_30201_, _20490_, _15325_);
  nor (_30202_, _26552_, _26443_);
  nor (_30203_, _30202_, _26553_);
  nor (_30204_, _30203_, _26104_);
  not (_30205_, _30204_);
  and (_30206_, _25851_, _25356_);
  or (_30207_, _30206_, _27777_);
  nor (_30208_, _30207_, _25862_);
  not (_30209_, _30208_);
  nor (_30210_, _27012_, _16693_);
  and (_30211_, _26750_, _25752_);
  and (_30212_, _26848_, _26815_);
  nor (_30213_, _30212_, _30211_);
  nor (_30214_, _30213_, _18078_);
  not (_30215_, _26728_);
  and (_30216_, _30213_, _18078_);
  or (_30217_, _30216_, _30215_);
  nor (_30218_, _30217_, _30214_);
  nor (_30219_, _30218_, _30210_);
  and (_30220_, _27264_, _25191_);
  nor (_30221_, _27242_, _25180_);
  or (_30222_, _30221_, _30220_);
  not (_30223_, _30222_);
  not (_30224_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30225_, _27078_, _30224_);
  nor (_30226_, _30225_, _18089_);
  or (_30227_, _30226_, _27067_);
  nor (_30228_, _30227_, _27079_);
  nor (_30229_, _28597_, _17707_);
  not (_30230_, _30229_);
  nor (_30231_, _27471_, _18078_);
  nor (_30232_, _27340_, _18579_);
  nor (_30233_, _30232_, _30231_);
  and (_30234_, _30233_, _30230_);
  and (_30235_, _27415_, _25169_);
  and (_30236_, _27427_, _18078_);
  nor (_30237_, _30236_, _30235_);
  and (_30238_, _30237_, _30234_);
  not (_30239_, _30238_);
  nor (_30240_, _30239_, _30228_);
  and (_30241_, _30240_, _30223_);
  and (_30242_, _30241_, _30219_);
  and (_30243_, _30242_, _30209_);
  and (_30244_, _30243_, _30205_);
  not (_30245_, _30244_);
  nor (_30246_, _30245_, _30201_);
  and (_30247_, _30246_, _30200_);
  not (_30248_, _30247_);
  or (_30249_, _30248_, _24949_);
  not (_30250_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_30251_, _24949_, _30250_);
  and (_30252_, _30251_, _27711_);
  and (_30253_, _30252_, _30249_);
  nor (_30254_, _27700_, _30250_);
  and (_30255_, _30110_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_30256_, _30121_, _24894_);
  not (_30257_, _30256_);
  nor (_30258_, _30257_, _28243_);
  not (_30259_, _24894_);
  or (_30260_, _30121_, _30259_);
  nor (_30261_, _30260_, _30250_);
  or (_30262_, _30261_, _30258_);
  and (_30263_, _30262_, _28285_);
  or (_30264_, _30263_, _30255_);
  and (_30265_, _30264_, _28347_);
  or (_30266_, _30265_, _30254_);
  or (_30267_, _30266_, _30253_);
  and (_08838_, _30267_, _35796_);
  and (_30268_, _23332_, _20661_);
  not (_30269_, _30268_);
  and (_30270_, _20522_, _15325_);
  nor (_30271_, _26618_, _25158_);
  and (_30272_, _26618_, _25158_);
  nor (_30273_, _30272_, _30271_);
  and (_30274_, _30273_, _26103_);
  not (_30275_, _30274_);
  not (_30276_, _25906_);
  nor (_30277_, _25895_, _25158_);
  nor (_30278_, _30277_, _27777_);
  and (_30279_, _30278_, _30276_);
  nor (_30280_, _25752_, _15879_);
  and (_30281_, _25752_, _17718_);
  nor (_30282_, _30281_, _30280_);
  nor (_30283_, _30282_, _27012_);
  and (_30284_, _26761_, _25752_);
  and (_30285_, _26859_, _26815_);
  nor (_30286_, _30285_, _30284_);
  and (_30287_, _30286_, _17707_);
  nor (_30288_, _30286_, _17707_);
  nor (_30289_, _30288_, _30287_);
  and (_30290_, _30289_, _26728_);
  nor (_30291_, _30290_, _30283_);
  nor (_30292_, _27080_, _17718_);
  not (_30293_, _30292_);
  nor (_30294_, _27089_, _27067_);
  and (_30295_, _30294_, _30293_);
  not (_30296_, _30295_);
  and (_30297_, _27264_, _25158_);
  nor (_30298_, _27242_, _25147_);
  not (_30299_, _30298_);
  and (_30300_, _27415_, _25103_);
  and (_30301_, _27427_, _17707_);
  nor (_30302_, _30301_, _30300_);
  nand (_30303_, _30302_, _30299_);
  nor (_30304_, _30303_, _30297_);
  nor (_30305_, _27340_, _18078_);
  not (_30306_, _30305_);
  nor (_30307_, _27471_, _17707_);
  nor (_30308_, _28597_, _17544_);
  nor (_30309_, _30308_, _30307_);
  and (_30310_, _30309_, _30306_);
  and (_30311_, _30310_, _30304_);
  and (_30312_, _30311_, _30296_);
  and (_30313_, _30312_, _30291_);
  not (_30314_, _30313_);
  nor (_30315_, _30314_, _30279_);
  and (_30316_, _30315_, _30275_);
  not (_30317_, _30316_);
  nor (_30318_, _30317_, _30270_);
  and (_30319_, _30318_, _30269_);
  not (_30320_, _30319_);
  or (_30321_, _30320_, _24949_);
  not (_30322_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_30323_, _24949_, _30322_);
  and (_30324_, _30323_, _27711_);
  and (_30325_, _30324_, _30321_);
  nor (_30326_, _27700_, _30322_);
  not (_30327_, _28285_);
  and (_30328_, _24773_, _24653_);
  and (_30329_, _30328_, _30259_);
  nor (_30330_, _30328_, _30259_);
  nor (_30331_, _30330_, _30329_);
  or (_30332_, _30331_, _30327_);
  and (_30333_, _30332_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_30334_, _30329_);
  nor (_30335_, _30334_, _28243_);
  and (_30336_, _30330_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_30337_, _30336_, _30335_);
  and (_30338_, _30337_, _28285_);
  or (_30339_, _30338_, _30333_);
  and (_30340_, _30339_, _28347_);
  or (_30341_, _30340_, _30326_);
  or (_30342_, _30341_, _30325_);
  and (_08849_, _30342_, _35796_);
  and (_30343_, _23419_, _20661_);
  not (_30344_, _30343_);
  and (_30345_, _20565_, _15325_);
  nor (_30346_, _26629_, _26279_);
  nor (_30347_, _30346_, _26640_);
  nor (_30348_, _30347_, _26104_);
  not (_30349_, _30348_);
  nor (_30350_, _25103_, _25092_);
  or (_30351_, _30350_, _25114_);
  and (_30352_, _30351_, _30276_);
  not (_30353_, _30352_);
  nor (_30354_, _27777_, _25917_);
  and (_30355_, _30354_, _30353_);
  nor (_30356_, _25752_, _16846_);
  and (_30357_, _25752_, _18121_);
  nor (_30358_, _30357_, _30356_);
  nor (_30359_, _30358_, _27012_);
  and (_30360_, _26772_, _25752_);
  and (_30361_, _26870_, _26815_);
  nor (_30362_, _30361_, _30360_);
  nor (_30363_, _30362_, _17544_);
  not (_30364_, _30363_);
  and (_30365_, _30362_, _17544_);
  nor (_30366_, _30365_, _30215_);
  and (_30367_, _30366_, _30364_);
  nor (_30368_, _30367_, _30359_);
  not (_30369_, _27154_);
  and (_30370_, _30369_, _27100_);
  nor (_30371_, _27154_, _27089_);
  nor (_30372_, _30371_, _17544_);
  nor (_30373_, _30372_, _30370_);
  nor (_30374_, _30373_, _27067_);
  and (_30375_, _27264_, _25092_);
  and (_30376_, _27415_, _25080_);
  nor (_30377_, _27242_, _25081_);
  and (_30378_, _27427_, _17544_);
  or (_30379_, _30378_, _30377_);
  or (_30380_, _30379_, _30376_);
  nor (_30381_, _30380_, _30375_);
  nor (_30382_, _27471_, _17544_);
  nor (_30383_, _27340_, _17707_);
  nor (_30384_, _28597_, _16533_);
  or (_30385_, _30384_, _30383_);
  nor (_30386_, _30385_, _30382_);
  and (_30387_, _30386_, _30381_);
  not (_30388_, _30387_);
  nor (_30389_, _30388_, _30374_);
  and (_30390_, _30389_, _30368_);
  not (_30391_, _30390_);
  nor (_30392_, _30391_, _30355_);
  and (_30393_, _30392_, _30349_);
  not (_30394_, _30393_);
  nor (_30395_, _30394_, _30345_);
  and (_30396_, _30395_, _30344_);
  not (_30397_, _30396_);
  or (_30398_, _30397_, _24949_);
  not (_30399_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_30400_, _24949_, _30399_);
  and (_30401_, _30400_, _27711_);
  and (_30402_, _30401_, _30398_);
  nor (_30403_, _27700_, _30399_);
  and (_30404_, _30259_, _24773_);
  nor (_30405_, _30404_, _30164_);
  or (_30406_, _30405_, _30327_);
  and (_30407_, _30406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_30408_, _24773_, _28296_);
  and (_30409_, _30408_, _30259_);
  not (_30410_, _30409_);
  nor (_30411_, _30410_, _28243_);
  or (_30412_, _30329_, _30164_);
  and (_30413_, _30412_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_30414_, _30413_, _30411_);
  and (_30415_, _30414_, _28285_);
  or (_30416_, _30415_, _30407_);
  and (_30417_, _30416_, _28347_);
  or (_30418_, _30417_, _30403_);
  or (_30419_, _30418_, _30402_);
  and (_08860_, _30419_, _35796_);
  and (_30420_, _23483_, _20661_);
  not (_30421_, _30420_);
  and (_30422_, _20597_, _15325_);
  nor (_30423_, _25939_, _25917_);
  not (_30424_, _30423_);
  nor (_30425_, _27777_, _25950_);
  and (_30426_, _30425_, _30424_);
  not (_30427_, _30426_);
  nor (_30428_, _26640_, _26246_);
  nor (_30429_, _30428_, _26651_);
  nor (_30430_, _30429_, _26104_);
  nor (_30431_, _25752_, _26115_);
  or (_30432_, _30431_, _27012_);
  nor (_30433_, _30432_, _27864_);
  or (_30434_, _25752_, _17544_);
  or (_30435_, _30361_, _26783_);
  and (_30436_, _30435_, _30434_);
  nor (_30437_, _30436_, _16544_);
  and (_30438_, _30436_, _16544_);
  or (_30439_, _30438_, _30215_);
  nor (_30440_, _30439_, _30437_);
  nor (_30441_, _30440_, _30433_);
  nor (_30442_, _30370_, _16533_);
  and (_30443_, _30370_, _16533_);
  nor (_30444_, _30443_, _30442_);
  nor (_30445_, _30444_, _27067_);
  and (_30446_, _27264_, _25048_);
  and (_30447_, _27415_, _25026_);
  nor (_30448_, _27242_, _25047_);
  and (_30449_, _27427_, _16533_);
  or (_30450_, _30449_, _30448_);
  or (_30451_, _30450_, _30447_);
  nor (_30452_, _30451_, _30446_);
  nor (_30453_, _27471_, _16533_);
  not (_30454_, _30453_);
  nor (_30455_, _28597_, _17358_);
  nor (_30456_, _27340_, _17544_);
  nor (_30457_, _30456_, _30455_);
  and (_30458_, _30457_, _30454_);
  and (_30459_, _30458_, _30452_);
  not (_30460_, _30459_);
  nor (_30461_, _30460_, _30445_);
  and (_30462_, _30461_, _30441_);
  not (_30463_, _30462_);
  nor (_30464_, _30463_, _30430_);
  and (_30465_, _30464_, _30427_);
  not (_30466_, _30465_);
  nor (_30467_, _30466_, _30422_);
  and (_30468_, _30467_, _30421_);
  not (_30469_, _30468_);
  or (_30470_, _30469_, _24949_);
  not (_30471_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_30472_, _24949_, _30471_);
  and (_30473_, _30472_, _27711_);
  and (_30474_, _30473_, _30470_);
  nor (_30475_, _27700_, _30471_);
  not (_30476_, _28316_);
  nand (_30477_, _30476_, _28285_);
  and (_30478_, _30477_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_30479_, _28306_, _24653_);
  and (_30480_, _30479_, _28827_);
  nor (_30481_, _28306_, _30471_);
  or (_30482_, _30481_, _30480_);
  and (_30483_, _30482_, _28285_);
  or (_30484_, _30483_, _30478_);
  and (_30485_, _30484_, _28347_);
  or (_30486_, _30485_, _30475_);
  or (_30487_, _30486_, _30474_);
  and (_08871_, _30487_, _35796_);
  and (_30488_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30489_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_30490_, _30489_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_30491_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_30492_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_30493_, _30492_, _30491_);
  and (_30494_, _30489_, _15260_);
  and (_30495_, _30494_, _30493_);
  and (_30496_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_30497_, _30496_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_30498_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_30499_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_30500_, _30499_, _30498_);
  and (_30501_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not (_30502_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_30503_, _30502_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30504_, _30503_, _30498_);
  and (_30505_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_30506_, _30505_, _30501_);
  and (_30507_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30508_, _30507_, _30498_);
  and (_30509_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_30510_, _30502_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30511_, _30510_, _30498_);
  and (_30512_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_30513_, _30512_, _30509_);
  and (_30514_, _30499_, _30498_);
  and (_30515_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_30516_, _30499_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_30517_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_30518_, _30517_, _30515_);
  and (_30519_, _30518_, _30513_);
  and (_30520_, _30519_, _30506_);
  and (_30521_, _30520_, _30497_);
  not (_30522_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30523_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _30522_);
  or (_30524_, _30523_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30525_, _30524_, _30521_);
  and (_30526_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_30527_, _30526_, _30525_);
  and (_30528_, _30527_, _30495_);
  not (_30529_, _30495_);
  and (_30530_, _30493_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_30531_, _30530_, _30529_);
  nor (_30532_, _30531_, _30528_);
  and (_30533_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_30534_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_30535_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_30536_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_30537_, _30536_, _30535_);
  and (_30538_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_30539_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_30540_, _30539_, _30538_);
  and (_30541_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_30542_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_30543_, _30542_, _30541_);
  and (_30544_, _30543_, _30540_);
  and (_30545_, _30544_, _30537_);
  nor (_30546_, _30545_, _30496_);
  and (_30547_, _30546_, _30522_);
  nor (_30548_, _30547_, _30534_);
  nor (_30549_, _30548_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30550_, _30549_, _30533_);
  nor (_30551_, _30550_, _30529_);
  and (_30552_, _30493_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_30553_, _30552_, _30529_);
  nor (_30554_, _30553_, _30551_);
  not (_30555_, _30554_);
  and (_30556_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30557_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_30558_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_30559_, _30558_, _30557_);
  and (_30560_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_30561_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_30562_, _30561_, _30560_);
  and (_30563_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_30564_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_30565_, _30564_, _30563_);
  and (_30566_, _30565_, _30562_);
  and (_30567_, _30566_, _30559_);
  nor (_30568_, _30567_, _30496_);
  nor (_30569_, _30568_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30570_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _30522_);
  nor (_30571_, _30570_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_30572_, _30571_);
  nor (_30573_, _30572_, _30569_);
  nor (_30574_, _30573_, _30556_);
  nor (_30575_, _30574_, _30529_);
  and (_30576_, _30493_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_30577_, _30576_, _30529_);
  nor (_30578_, _30577_, _30575_);
  and (_30579_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30580_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_30581_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_30582_, _30581_, _30580_);
  and (_30583_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_30584_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_30585_, _30584_, _30583_);
  and (_30586_, _30585_, _30582_);
  and (_30587_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_30588_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_30589_, _30588_, _30587_);
  and (_30590_, _30589_, _30586_);
  nor (_30591_, _30590_, _30496_);
  nor (_30592_, _30591_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30593_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _30522_);
  nor (_30594_, _30593_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_30595_, _30594_);
  nor (_30596_, _30595_, _30592_);
  nor (_30597_, _30596_, _30579_);
  nor (_30598_, _30597_, _30529_);
  and (_30599_, _30493_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_30600_, _30599_, _30529_);
  nor (_30601_, _30600_, _30598_);
  not (_30602_, _30601_);
  and (_30603_, _30602_, _30578_);
  and (_30604_, _30603_, _30555_);
  and (_30605_, _30604_, _30532_);
  and (_30606_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30607_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_30608_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_30609_, _30608_, _30607_);
  and (_30610_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_30611_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_30612_, _30611_, _30610_);
  and (_30613_, _30612_, _30609_);
  and (_30614_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_30615_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_30616_, _30615_, _30614_);
  and (_30617_, _30616_, _30613_);
  nor (_30618_, _30617_, _30496_);
  nor (_30619_, _30618_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30620_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _30522_);
  nor (_30621_, _30620_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_30622_, _30621_);
  nor (_30623_, _30622_, _30619_);
  nor (_30624_, _30623_, _30606_);
  nor (_30625_, _30624_, _30529_);
  and (_30626_, _30493_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_30627_, _30626_, _30529_);
  nor (_30628_, _30627_, _30625_);
  not (_30629_, _30628_);
  and (_30630_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30631_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_30632_, _30496_);
  and (_30633_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_30634_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_30635_, _30634_, _30633_);
  and (_30636_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_30637_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_30638_, _30637_, _30636_);
  and (_30639_, _30638_, _30635_);
  and (_30640_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_30641_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_30642_, _30641_, _30640_);
  and (_30643_, _30642_, _30639_);
  and (_30644_, _30643_, _30632_);
  nor (_30645_, _30644_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30646_, _30645_, _30631_);
  nor (_30647_, _30646_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30649_, _30647_, _30630_);
  nor (_30650_, _30649_, _30529_);
  and (_30652_, _30493_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_30653_, _30652_, _30529_);
  nor (_30655_, _30653_, _30650_);
  not (_30656_, _30655_);
  and (_30658_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30659_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_30660_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_30661_, _30660_, _30659_);
  and (_30662_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_30663_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_30664_, _30663_, _30662_);
  and (_30665_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_30666_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_30667_, _30666_, _30665_);
  and (_30668_, _30667_, _30664_);
  and (_30669_, _30668_, _30661_);
  nor (_30670_, _30669_, _30496_);
  nor (_30671_, _30670_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30672_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _30522_);
  nor (_30673_, _30672_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_30674_, _30673_);
  nor (_30675_, _30674_, _30671_);
  nor (_30676_, _30675_, _30658_);
  nor (_30677_, _30676_, _30529_);
  and (_30678_, _30493_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_30679_, _30678_, _30529_);
  nor (_30680_, _30679_, _30677_);
  and (_30681_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30682_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_30683_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_30684_, _30683_, _30682_);
  and (_30685_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_30686_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_30687_, _30686_, _30685_);
  and (_30688_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_30689_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_30690_, _30689_, _30688_);
  and (_30691_, _30690_, _30687_);
  and (_30692_, _30691_, _30684_);
  nor (_30693_, _30692_, _30496_);
  nor (_30694_, _30693_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30695_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _30522_);
  nor (_30696_, _30695_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_30697_, _30696_);
  nor (_30698_, _30697_, _30694_);
  nor (_30699_, _30698_, _30681_);
  nor (_30700_, _30699_, _30529_);
  and (_30701_, _30493_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_30702_, _30701_, _30529_);
  nor (_30703_, _30702_, _30700_);
  and (_30704_, _30703_, _30680_);
  and (_30705_, _30704_, _30656_);
  and (_30706_, _30705_, _30629_);
  and (_30707_, _30706_, _30605_);
  not (_30708_, _30706_);
  not (_30709_, _30532_);
  not (_30710_, _30578_);
  nor (_30711_, _30554_, _30710_);
  and (_30712_, _30601_, _30711_);
  and (_30713_, _30712_, _30709_);
  nor (_30714_, _30601_, _30578_);
  and (_30715_, _30714_, _30554_);
  and (_30716_, _30715_, _30709_);
  nor (_30717_, _30716_, _30713_);
  nor (_30718_, _30717_, _30708_);
  nor (_30719_, _30718_, _30707_);
  and (_30720_, _30712_, _30532_);
  not (_30721_, _30680_);
  and (_30722_, _30703_, _30721_);
  and (_30723_, _30655_, _30628_);
  and (_30724_, _30723_, _30722_);
  and (_30725_, _30724_, _30720_);
  and (_30726_, _30724_, _30605_);
  nor (_30727_, _30726_, _30725_);
  and (_30728_, _30727_, _30719_);
  nor (_30729_, _30728_, _30490_);
  not (_30730_, _30729_);
  not (_30731_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_30732_, _15260_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_30733_, _30732_, _30731_);
  and (_30734_, _30554_, _30710_);
  and (_30735_, _30723_, _30704_);
  and (_30736_, _30735_, _30734_);
  and (_30737_, _30736_, _30733_);
  and (_30738_, _30726_, _15260_);
  and (_30739_, _30725_, _15260_);
  nor (_30740_, _30739_, _30738_);
  nor (_30741_, _30740_, _30489_);
  nor (_30742_, _30741_, _30737_);
  and (_30743_, _30742_, _30730_);
  nor (_30744_, _30743_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30745_, _30744_, _30488_);
  and (_30746_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30747_, _30705_, _30628_);
  and (_30748_, _30747_, _30713_);
  and (_30749_, _30655_, _30629_);
  and (_30750_, _30749_, _30722_);
  and (_30751_, _30750_, _30720_);
  nor (_30752_, _30751_, _30748_);
  and (_30753_, _30554_, _30578_);
  and (_30754_, _30753_, _30602_);
  and (_30755_, _30754_, _30747_);
  not (_30756_, _30703_);
  and (_30757_, _30605_, _30756_);
  nor (_30758_, _30757_, _30755_);
  and (_30759_, _30758_, _30752_);
  and (_30760_, _30720_, _30747_);
  and (_30761_, _30734_, _30601_);
  and (_30762_, _30761_, _30709_);
  and (_30763_, _30762_, _30705_);
  nor (_30764_, _30763_, _30760_);
  and (_30765_, _30601_, _30710_);
  and (_30766_, _30765_, _30555_);
  and (_30767_, _30766_, _30532_);
  and (_30768_, _30767_, _30750_);
  and (_30769_, _30734_, _30532_);
  and (_30770_, _30769_, _30602_);
  and (_30771_, _30770_, _30750_);
  nor (_30772_, _30771_, _30768_);
  and (_30773_, _30772_, _30764_);
  and (_30774_, _30773_, _30759_);
  and (_30775_, _30735_, _30754_);
  and (_30776_, _30775_, _30532_);
  not (_30777_, _30735_);
  and (_30778_, _30754_, _30709_);
  and (_30779_, _30753_, _30601_);
  and (_30780_, _30779_, _30709_);
  nor (_30781_, _30780_, _30778_);
  nor (_30782_, _30781_, _30777_);
  nor (_30783_, _30782_, _30776_);
  and (_30784_, _30714_, _30555_);
  and (_30785_, _30784_, _30532_);
  and (_30786_, _30785_, _30750_);
  not (_30787_, _30786_);
  and (_30788_, _30779_, _30532_);
  and (_30789_, _30788_, _30750_);
  nor (_30790_, _30680_, _30655_);
  and (_30791_, _30790_, _30703_);
  and (_30792_, _30791_, _30532_);
  and (_30793_, _30792_, _30604_);
  nor (_30794_, _30793_, _30789_);
  and (_30795_, _30794_, _30787_);
  and (_30796_, _30795_, _30783_);
  and (_30797_, _30796_, _30774_);
  and (_30798_, _30766_, _30709_);
  and (_30799_, _30798_, _30750_);
  and (_30800_, _30780_, _30750_);
  nor (_30801_, _30800_, _30799_);
  and (_30802_, _30761_, _30532_);
  and (_30803_, _30802_, _30750_);
  and (_30804_, _30735_, _30604_);
  nor (_30805_, _30804_, _30803_);
  and (_30806_, _30805_, _30801_);
  and (_30807_, _30604_, _30709_);
  and (_30808_, _30807_, _30747_);
  and (_30809_, _30767_, _30747_);
  nor (_30810_, _30809_, _30808_);
  and (_30811_, _30716_, _30747_);
  and (_30812_, _30802_, _30705_);
  nor (_30813_, _30812_, _30811_);
  and (_30814_, _30813_, _30810_);
  and (_30815_, _30814_, _30806_);
  and (_30816_, _30735_, _30766_);
  and (_30817_, _30770_, _30705_);
  nor (_30818_, _30817_, _30816_);
  not (_30819_, _30818_);
  and (_30820_, _30711_, _30709_);
  and (_30821_, _30820_, _30750_);
  nor (_30822_, _30821_, _30819_);
  not (_30823_, _30750_);
  nor (_30824_, _30762_, _30754_);
  nor (_30825_, _30824_, _30823_);
  and (_30826_, _30798_, _30747_);
  and (_30827_, _30605_, _30747_);
  nor (_30828_, _30827_, _30826_);
  not (_30829_, _30828_);
  nor (_30830_, _30829_, _30825_);
  and (_30831_, _30830_, _30822_);
  and (_30832_, _30831_, _30815_);
  and (_30833_, _30832_, _30797_);
  nor (_30834_, _30833_, _30490_);
  and (_30835_, _30732_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_30836_, _30835_, _30755_);
  not (_30837_, _30836_);
  nor (_30838_, _30601_, _30709_);
  and (_30839_, _30838_, _30753_);
  and (_30840_, _30735_, _30839_);
  and (_30841_, _30780_, _30735_);
  nor (_30842_, _30841_, _30840_);
  not (_30843_, _30733_);
  nor (_30844_, _30843_, _30842_);
  nor (_30845_, _30844_, _30737_);
  and (_30846_, _30845_, _30837_);
  not (_30847_, _30846_);
  nor (_30848_, _30847_, _30834_);
  nor (_30849_, _30848_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30850_, _30849_, _30746_);
  and (_30851_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30852_, _30703_, _30709_);
  and (_30853_, _30852_, _30790_);
  and (_30854_, _30853_, _30604_);
  and (_30855_, _30791_, _30779_);
  nor (_30856_, _30855_, _30854_);
  and (_30857_, _30791_, _30720_);
  nor (_30858_, _30857_, _30755_);
  and (_30859_, _30858_, _30856_);
  and (_30860_, _30791_, _30766_);
  and (_30861_, _30853_, _30712_);
  nor (_30862_, _30861_, _30860_);
  not (_30863_, _30862_);
  not (_30864_, _30791_);
  nor (_30865_, _30824_, _30864_);
  nor (_30866_, _30865_, _30863_);
  and (_30867_, _30866_, _30859_);
  and (_30868_, _30791_, _30770_);
  not (_30869_, _30868_);
  and (_30870_, _30798_, _30735_);
  not (_30871_, _30792_);
  nor (_30872_, _30784_, _30761_);
  nor (_30873_, _30872_, _30871_);
  nor (_30874_, _30873_, _30870_);
  and (_30875_, _30874_, _30869_);
  and (_30876_, _30875_, _30719_);
  and (_30877_, _30876_, _30867_);
  nor (_30878_, _30877_, _30490_);
  and (_30879_, _30755_, _30732_);
  and (_30880_, _30879_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_30881_, _30733_, _30715_);
  and (_30882_, _30881_, _30735_);
  or (_30883_, _30882_, _30880_);
  nor (_30884_, _30883_, _30878_);
  nor (_30885_, _30884_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30886_, _30885_, _30851_);
  nor (_30887_, _30886_, _30850_);
  and (_30888_, _30887_, _30745_);
  and (_09422_, _30888_, _35796_);
  and (_30889_, _24521_, _24378_);
  not (_30890_, _24009_);
  nor (_30891_, _30890_, _23877_);
  and (_30892_, _30891_, _30889_);
  and (_30893_, _30892_, _24202_);
  and (_30894_, _30893_, _29466_);
  and (_30895_, _30894_, _27700_);
  and (_30896_, _30895_, _27668_);
  or (_30897_, _20661_, _15325_);
  and (_30898_, _25004_, _20639_);
  or (_30899_, _27329_, _27460_);
  or (_30900_, _30899_, _30898_);
  or (_30901_, _30900_, _30897_);
  nor (_30902_, _30901_, _28596_);
  nor (_30903_, _30902_, _17358_);
  not (_30904_, _30903_);
  and (_30905_, _30904_, _27449_);
  and (_30906_, _30905_, _27286_);
  and (_30907_, _30906_, _27045_);
  not (_30908_, _30907_);
  and (_30909_, _30908_, _30896_);
  and (_30910_, _27711_, _24202_);
  and (_30911_, _30892_, _29466_);
  and (_30912_, _30911_, _30910_);
  not (_30913_, _30912_);
  and (_30914_, _30913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_30915_, _30902_, _16533_);
  not (_30916_, _30915_);
  and (_30917_, _30916_, _30452_);
  and (_30918_, _30917_, _30441_);
  nor (_30919_, _30918_, _30913_);
  nor (_30920_, _30919_, _30914_);
  and (_30921_, _30913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_30922_, _30902_, _17544_);
  not (_30923_, _30922_);
  and (_30924_, _30923_, _30381_);
  and (_30925_, _30924_, _30368_);
  nor (_30926_, _30925_, _30913_);
  nor (_30927_, _30926_, _30921_);
  and (_30928_, _30913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_30929_, _30902_, _17707_);
  not (_30930_, _30929_);
  and (_30931_, _30930_, _30304_);
  and (_30932_, _30931_, _30291_);
  nor (_30933_, _30932_, _30913_);
  nor (_30934_, _30933_, _30928_);
  and (_30935_, _30913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_30936_, _30902_, _18078_);
  nor (_30937_, _30936_, _30222_);
  and (_30938_, _30937_, _30237_);
  and (_30939_, _30938_, _30219_);
  nor (_30940_, _30939_, _30913_);
  nor (_30941_, _30940_, _30935_);
  and (_30942_, _30913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_30943_, _30902_, _18579_);
  not (_30944_, _30943_);
  and (_30945_, _30944_, _29773_);
  and (_30946_, _30945_, _29806_);
  and (_30947_, _30946_, _29685_);
  nor (_30948_, _30947_, _30913_);
  nor (_30949_, _30948_, _30942_);
  and (_30950_, _30913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_30951_, _30902_, _18416_);
  nor (_30952_, _30951_, _29197_);
  and (_30953_, _30952_, _29101_);
  and (_30954_, _30953_, _29013_);
  nor (_30955_, _30954_, _30913_);
  nor (_30956_, _30955_, _30950_);
  nor (_30957_, _30912_, _24598_);
  nor (_30958_, _30902_, _18960_);
  not (_30959_, _30958_);
  and (_30960_, _30959_, _28595_);
  and (_30961_, _30960_, _28572_);
  and (_30962_, _30961_, _28549_);
  not (_30963_, _30962_);
  and (_30964_, _30963_, _30912_);
  nor (_30965_, _30964_, _30957_);
  and (_30966_, _30965_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_30967_, _30966_, _30956_);
  and (_30968_, _30967_, _30949_);
  and (_30969_, _30968_, _30941_);
  and (_30970_, _30969_, _30934_);
  and (_30971_, _30970_, _30927_);
  and (_30972_, _30971_, _30920_);
  nor (_30973_, _30912_, _23559_);
  and (_30974_, _30973_, _30972_);
  nor (_30975_, _30973_, _30972_);
  nor (_30976_, _30975_, _30974_);
  and (_30977_, _30976_, _23548_);
  nor (_30978_, _30977_, _23669_);
  nor (_30979_, _30978_, _30912_);
  nor (_30980_, _30979_, _30909_);
  nor (_09443_, _30980_, rst);
  not (_30981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_30982_, _30965_, _30981_);
  nor (_30983_, _30965_, _30981_);
  nor (_30984_, _30983_, _30982_);
  and (_30985_, _30984_, _23548_);
  nor (_30986_, _30985_, _24609_);
  nor (_30987_, _30986_, _30912_);
  nor (_30988_, _30987_, _30964_);
  nand (_10555_, _30988_, _35796_);
  nor (_30989_, _30966_, _30956_);
  nor (_30990_, _30989_, _30967_);
  nor (_30991_, _30990_, _23537_);
  nor (_30992_, _30991_, _24686_);
  nor (_30993_, _30992_, _30912_);
  nor (_30994_, _30993_, _30955_);
  nand (_10566_, _30994_, _35796_);
  nor (_30995_, _30967_, _30949_);
  nor (_30996_, _30995_, _30968_);
  nor (_30997_, _30996_, _23537_);
  nor (_30998_, _30997_, _24806_);
  nor (_30999_, _30998_, _30912_);
  nor (_31000_, _30999_, _30948_);
  nand (_10577_, _31000_, _35796_);
  nor (_31001_, _30968_, _30941_);
  nor (_31002_, _31001_, _30969_);
  nor (_31003_, _31002_, _23537_);
  nor (_31004_, _31003_, _24110_);
  nor (_31005_, _31004_, _30912_);
  nor (_31006_, _31005_, _30940_);
  nor (_10588_, _31006_, rst);
  nor (_31007_, _30969_, _30934_);
  nor (_31008_, _31007_, _30970_);
  nor (_31009_, _31008_, _23537_);
  nor (_31010_, _31009_, _24312_);
  nor (_31011_, _31010_, _30912_);
  nor (_31012_, _31011_, _30933_);
  nor (_10599_, _31012_, rst);
  nor (_31013_, _30970_, _30927_);
  nor (_31014_, _31013_, _30971_);
  nor (_31015_, _31014_, _23537_);
  nor (_31016_, _31015_, _24432_);
  nor (_31017_, _31016_, _30912_);
  nor (_31018_, _31017_, _30926_);
  nor (_10610_, _31018_, rst);
  nor (_31019_, _30971_, _30920_);
  nor (_31020_, _31019_, _30972_);
  nor (_31021_, _31020_, _23537_);
  nor (_31022_, _31021_, _23921_);
  nor (_31023_, _31022_, _30912_);
  nor (_31024_, _31023_, _30919_);
  nor (_10621_, _31024_, rst);
  and (_31025_, _30910_, _30256_);
  nand (_31026_, _31025_, _30892_);
  nor (_31027_, _31026_, _27635_);
  and (_31028_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15260_);
  and (_31029_, _31028_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_31030_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_31031_, _31030_, _31029_);
  or (_31032_, _31031_, _31027_);
  nor (_31033_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_31034_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_31035_, _31034_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31036_, _31035_, _31033_);
  nor (_31037_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_31038_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_31039_, _31038_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31040_, _31039_, _31037_);
  nor (_31041_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_31042_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_31043_, _31042_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31044_, _31043_, _31041_);
  not (_31045_, _31044_);
  nor (_31046_, _31045_, _27799_);
  nor (_31047_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_31048_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_31049_, _31048_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31050_, _31049_, _31047_);
  and (_31051_, _31050_, _31046_);
  nor (_31052_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_31053_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_31054_, _31053_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31055_, _31054_, _31052_);
  and (_31056_, _31055_, _31051_);
  and (_31057_, _31056_, _31040_);
  nor (_31058_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_31059_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_31060_, _31059_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31061_, _31060_, _31058_);
  and (_31062_, _31061_, _31057_);
  and (_31063_, _31062_, _31036_);
  nor (_31064_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_31065_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_31066_, _31065_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31067_, _31066_, _31064_);
  and (_31068_, _31067_, _31063_);
  nor (_31069_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_31070_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_31071_, _31070_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_31072_, _31071_, _31069_);
  or (_31073_, _31072_, _31068_);
  nand (_31074_, _31072_, _31068_);
  and (_31075_, _31074_, _25015_);
  and (_31076_, _31075_, _31073_);
  not (_31077_, _31076_);
  and (_31078_, _20351_, _15325_);
  nor (_31079_, _17358_, _16042_);
  and (_31080_, _31079_, _26793_);
  and (_31081_, _31080_, _26333_);
  and (_31082_, _31081_, _26377_);
  and (_31083_, _31082_, _26564_);
  nor (_31084_, _31083_, _26815_);
  and (_31085_, _25752_, _15879_);
  nor (_31086_, _31085_, _31084_);
  and (_31087_, _26881_, _17358_);
  and (_31088_, _16693_, _15716_);
  and (_31089_, _17010_, _16042_);
  and (_31090_, _31089_, _31088_);
  and (_31091_, _31090_, _31087_);
  and (_31092_, _16846_, _15879_);
  and (_31093_, _31092_, _31091_);
  nor (_31094_, _31093_, _25752_);
  and (_31095_, _25752_, _16846_);
  nor (_31096_, _31095_, _31094_);
  and (_31097_, _31096_, _31086_);
  nor (_31098_, _25752_, _16217_);
  and (_31099_, _25752_, _16217_);
  nor (_31100_, _31099_, _31098_);
  and (_31101_, _31100_, _31097_);
  and (_31102_, _31101_, _26957_);
  nor (_31103_, _31101_, _26957_);
  nor (_31104_, _31103_, _31102_);
  and (_31105_, _31104_, _26728_);
  and (_31106_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_31107_, _25752_, _26957_);
  nor (_31108_, _31107_, _27897_);
  nor (_31109_, _31108_, _27012_);
  nor (_31110_, _28052_, _18078_);
  nor (_31111_, _27471_, _17184_);
  or (_31112_, _31111_, _31110_);
  or (_31113_, _31112_, _31109_);
  nor (_31114_, _31113_, _31106_);
  not (_31115_, _31114_);
  nor (_31116_, _31115_, _31105_);
  not (_31117_, _31116_);
  nor (_31118_, _31117_, _31078_);
  and (_31119_, _31118_, _31077_);
  nand (_31120_, _31119_, _31029_);
  and (_31121_, _31120_, _35796_);
  and (_12457_, _31121_, _31032_);
  and (_31122_, _30910_, _30175_);
  and (_31123_, _31122_, _30892_);
  nor (_31124_, _31123_, _31029_);
  not (_31125_, _31124_);
  nand (_31126_, _31125_, _27635_);
  not (_31127_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_31128_, _31124_, _31127_);
  and (_31129_, _31128_, _35796_);
  and (_12477_, _31129_, _31126_);
  nor (_31130_, _31026_, _28739_);
  and (_31131_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_31132_, _31131_, _31029_);
  or (_31133_, _31132_, _31130_);
  and (_31134_, _22957_, _20661_);
  not (_31135_, _31134_);
  and (_31136_, _31045_, _27799_);
  nor (_31137_, _31136_, _31046_);
  and (_31138_, _31137_, _25015_);
  nor (_31139_, _27897_, _26990_);
  not (_31140_, _31139_);
  nor (_31141_, _31140_, _26902_);
  nor (_31142_, _31141_, _26301_);
  and (_31143_, _31141_, _26301_);
  nor (_31144_, _31143_, _31142_);
  and (_31145_, _31144_, _26728_);
  nor (_31146_, _27471_, _16042_);
  and (_31147_, _20128_, _15325_);
  nor (_31148_, _28052_, _17707_);
  nor (_31149_, _27012_, _18960_);
  or (_31150_, _31149_, _31148_);
  or (_31151_, _31150_, _31147_);
  nor (_31152_, _31151_, _31146_);
  not (_31153_, _31152_);
  nor (_31154_, _31153_, _31145_);
  not (_31155_, _31154_);
  nor (_31156_, _31155_, _31138_);
  and (_31157_, _31156_, _31135_);
  nand (_31158_, _31157_, _31029_);
  and (_31159_, _31158_, _35796_);
  and (_13391_, _31159_, _31133_);
  nor (_31160_, _31026_, _29380_);
  and (_31161_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_31162_, _31161_, _31029_);
  or (_31163_, _31162_, _31160_);
  nor (_31164_, _31050_, _31046_);
  not (_31165_, _31164_);
  nor (_31166_, _31051_, _27777_);
  and (_31167_, _31166_, _31165_);
  not (_31168_, _31167_);
  and (_31169_, _21960_, _20661_);
  and (_31170_, _31080_, _25752_);
  and (_31171_, _31087_, _16042_);
  and (_31172_, _31171_, _26815_);
  nor (_31173_, _31172_, _31170_);
  nor (_31174_, _31173_, _26333_);
  and (_31175_, _31173_, _26333_);
  nor (_31176_, _31175_, _31174_);
  nor (_31177_, _31176_, _30215_);
  nor (_31178_, _27471_, _17010_);
  and (_31179_, _20160_, _15325_);
  nor (_31180_, _28052_, _17544_);
  nor (_31181_, _27012_, _18416_);
  or (_31182_, _31181_, _31180_);
  or (_31183_, _31182_, _31179_);
  nor (_31184_, _31183_, _31178_);
  not (_31185_, _31184_);
  nor (_31186_, _31185_, _31177_);
  not (_31187_, _31186_);
  nor (_31188_, _31187_, _31169_);
  and (_31189_, _31188_, _31168_);
  nand (_31190_, _31189_, _31029_);
  and (_31191_, _31190_, _35796_);
  and (_13402_, _31191_, _31163_);
  nor (_31192_, _31026_, _30024_);
  and (_31193_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_31194_, _31193_, _31029_);
  or (_31195_, _31194_, _31192_);
  nor (_31196_, _31055_, _31051_);
  nor (_31197_, _31196_, _31056_);
  and (_31198_, _31197_, _25015_);
  not (_31199_, _31198_);
  and (_31200_, _31171_, _17010_);
  and (_31201_, _31200_, _26815_);
  and (_31202_, _31081_, _25752_);
  nor (_31203_, _31202_, _31201_);
  and (_31204_, _31203_, _15716_);
  nor (_31205_, _31203_, _15716_);
  nor (_31206_, _31205_, _31204_);
  and (_31207_, _31206_, _26728_);
  not (_31208_, _31207_);
  nor (_31209_, _27012_, _18579_);
  and (_31210_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_31211_, _31210_, _31209_);
  and (_31212_, _20192_, _15325_);
  nor (_31213_, _28052_, _16533_);
  nor (_31214_, _27471_, _15716_);
  or (_31215_, _31214_, _31213_);
  nor (_31216_, _31215_, _31212_);
  and (_31217_, _31216_, _31211_);
  and (_31218_, _31217_, _31208_);
  and (_31219_, _31218_, _31199_);
  nand (_31220_, _31219_, _31029_);
  and (_31221_, _31220_, _35796_);
  and (_13413_, _31221_, _31195_);
  nor (_31222_, _31026_, _30247_);
  and (_31223_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_31224_, _31223_, _31029_);
  or (_31225_, _31224_, _31222_);
  nor (_31226_, _31056_, _31040_);
  nor (_31227_, _31226_, _31057_);
  and (_31228_, _31227_, _25015_);
  not (_31229_, _31228_);
  and (_31230_, _20224_, _15325_);
  nor (_31231_, _31082_, _26564_);
  not (_31232_, _31231_);
  and (_31233_, _31232_, _31084_);
  and (_31234_, _31200_, _15716_);
  nor (_31235_, _31234_, _16693_);
  nor (_31236_, _31235_, _31091_);
  nor (_31237_, _31236_, _25752_);
  nor (_31238_, _31237_, _31233_);
  nor (_31239_, _31238_, _30215_);
  nor (_31240_, _27471_, _16693_);
  nor (_31241_, _27012_, _18078_);
  and (_31242_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_31243_, _31242_, _31241_);
  or (_31244_, _31243_, _28062_);
  nor (_31245_, _31244_, _31240_);
  not (_31246_, _31245_);
  nor (_31247_, _31246_, _31239_);
  not (_31248_, _31247_);
  nor (_31249_, _31248_, _31230_);
  and (_31250_, _31249_, _31229_);
  nand (_31251_, _31250_, _31029_);
  and (_31252_, _31251_, _35796_);
  and (_13424_, _31252_, _31225_);
  nor (_31253_, _31026_, _30319_);
  and (_31254_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_31255_, _31254_, _31029_);
  or (_31256_, _31255_, _31253_);
  nor (_31257_, _31061_, _31057_);
  nor (_31258_, _31257_, _31062_);
  and (_31259_, _31258_, _25015_);
  not (_31260_, _31259_);
  and (_31261_, _20256_, _15325_);
  nor (_31262_, _31091_, _25752_);
  nor (_31263_, _31262_, _31084_);
  nor (_31264_, _31263_, _26159_);
  and (_31265_, _31263_, _26159_);
  nor (_31266_, _31265_, _31264_);
  and (_31267_, _31266_, _26728_);
  and (_31268_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_31269_, _25752_, _17718_);
  or (_31270_, _31269_, _27012_);
  nor (_31271_, _31270_, _31085_);
  nor (_31272_, _28052_, _18960_);
  nor (_31273_, _27471_, _15879_);
  or (_31274_, _31273_, _31272_);
  or (_31275_, _31274_, _31271_);
  nor (_31276_, _31275_, _31268_);
  not (_31277_, _31276_);
  nor (_31278_, _31277_, _31267_);
  not (_31279_, _31278_);
  nor (_31280_, _31279_, _31261_);
  and (_31281_, _31280_, _31260_);
  nand (_31282_, _31281_, _31029_);
  and (_31283_, _31282_, _35796_);
  and (_13435_, _31283_, _31256_);
  nor (_31284_, _31026_, _30396_);
  and (_31285_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_31286_, _31285_, _31029_);
  or (_31287_, _31286_, _31284_);
  nor (_31288_, _31062_, _31036_);
  not (_31289_, _31288_);
  nor (_31290_, _31063_, _27777_);
  and (_31291_, _31290_, _31289_);
  not (_31292_, _31291_);
  and (_31293_, _20287_, _15325_);
  and (_31294_, _31091_, _15879_);
  nor (_31295_, _31294_, _25752_);
  not (_31296_, _31295_);
  and (_31297_, _31296_, _31086_);
  and (_31298_, _31297_, _16846_);
  nor (_31299_, _31297_, _16846_);
  nor (_31300_, _31299_, _31298_);
  nor (_31301_, _31300_, _30215_);
  and (_31302_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_31303_, _25752_, _18121_);
  or (_31304_, _31303_, _27012_);
  nor (_31305_, _31304_, _31095_);
  nor (_31306_, _28052_, _18416_);
  nor (_31307_, _27471_, _16846_);
  or (_31308_, _31307_, _31306_);
  or (_31309_, _31308_, _31305_);
  nor (_31310_, _31309_, _31302_);
  not (_31311_, _31310_);
  nor (_31312_, _31311_, _31301_);
  not (_31313_, _31312_);
  nor (_31314_, _31313_, _31293_);
  and (_31315_, _31314_, _31292_);
  nand (_31316_, _31315_, _31029_);
  and (_31317_, _31316_, _35796_);
  and (_13446_, _31317_, _31287_);
  nor (_31318_, _31026_, _30468_);
  and (_31319_, _31026_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_31320_, _31319_, _31029_);
  or (_31321_, _31320_, _31318_);
  nor (_31322_, _31067_, _31063_);
  nor (_31323_, _31322_, _31068_);
  and (_31324_, _31323_, _25015_);
  not (_31325_, _31324_);
  and (_31326_, _20319_, _15325_);
  and (_31327_, _31097_, _16217_);
  nor (_31328_, _31097_, _16217_);
  nor (_31329_, _31328_, _31327_);
  nor (_31330_, _31329_, _30215_);
  and (_31331_, _20661_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_31332_, _25752_, _16544_);
  or (_31333_, _31332_, _27012_);
  nor (_31334_, _31333_, _31099_);
  nor (_31335_, _28052_, _18579_);
  nor (_31336_, _27471_, _16217_);
  or (_31337_, _31336_, _31335_);
  or (_31338_, _31337_, _31334_);
  nor (_31339_, _31338_, _31331_);
  not (_31340_, _31339_);
  nor (_31341_, _31340_, _31330_);
  not (_31342_, _31341_);
  nor (_31343_, _31342_, _31326_);
  and (_31344_, _31343_, _31325_);
  nand (_31345_, _31344_, _31029_);
  and (_31346_, _31345_, _35796_);
  and (_13457_, _31346_, _31321_);
  nand (_31347_, _31125_, _28739_);
  not (_31348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_31349_, _31124_, _31348_);
  and (_31350_, _31349_, _35796_);
  and (_13468_, _31350_, _31347_);
  nand (_31351_, _31125_, _29380_);
  not (_31352_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_31353_, _31124_, _31352_);
  and (_31354_, _31353_, _35796_);
  and (_13479_, _31354_, _31351_);
  nand (_31355_, _31125_, _30024_);
  not (_31356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_31357_, _31124_, _31356_);
  and (_31358_, _31357_, _35796_);
  and (_13490_, _31358_, _31355_);
  nand (_31359_, _31125_, _30247_);
  or (_31360_, _31125_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_31361_, _31360_, _35796_);
  and (_13501_, _31361_, _31359_);
  nand (_31362_, _31125_, _30319_);
  or (_31363_, _31125_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_31364_, _31363_, _35796_);
  and (_13511_, _31364_, _31362_);
  nand (_31365_, _31125_, _30396_);
  or (_31366_, _31125_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_31367_, _31366_, _35796_);
  and (_13522_, _31367_, _31365_);
  nand (_31368_, _31125_, _30468_);
  or (_31369_, _31125_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_31370_, _31369_, _35796_);
  and (_13533_, _31370_, _31368_);
  and (_31371_, _24521_, _24389_);
  and (_31372_, _31371_, _24020_);
  and (_31373_, _31372_, _28347_);
  nor (_31374_, _30476_, _28243_);
  not (_31375_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_31376_, _28316_, _31375_);
  or (_31377_, _31376_, _31374_);
  and (_31378_, _31377_, _31373_);
  nor (_31379_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_31380_, _31379_);
  nand (_31381_, _31380_, _28243_);
  and (_31382_, _31379_, _31375_);
  nor (_31383_, _31382_, _31373_);
  and (_31384_, _31383_, _31381_);
  and (_31385_, _27711_, _24916_);
  and (_31386_, _31385_, _31372_);
  or (_31387_, _31386_, _31384_);
  or (_31388_, _31387_, _31378_);
  nand (_31389_, _31386_, _30907_);
  and (_31390_, _31389_, _31388_);
  and (_16434_, _31390_, _35796_);
  not (_31391_, _31386_);
  not (_31392_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_31393_, _31373_, _29466_);
  nand (_31394_, _31393_, _31392_);
  and (_31395_, _31394_, _31391_);
  or (_31396_, _31393_, _28827_);
  and (_31397_, _31396_, _31395_);
  nor (_31398_, _31391_, _30954_);
  or (_31399_, _31398_, _31397_);
  and (_21361_, _31399_, _35796_);
  or (_31400_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_31401_, _20415_, _20383_);
  or (_31402_, _31401_, _20447_);
  or (_31403_, _31402_, _20490_);
  or (_31404_, _31403_, _20522_);
  or (_31405_, _31404_, _20565_);
  or (_31406_, _31405_, _20597_);
  or (_31407_, _31406_, _20053_);
  and (_31408_, _31407_, _15325_);
  and (_31409_, _27831_, _26662_);
  not (_31410_, _26662_);
  and (_31411_, _27842_, _31410_);
  or (_31412_, _31411_, _31409_);
  and (_31413_, _31412_, _26103_);
  not (_31414_, _25993_);
  nand (_31415_, _25972_, _31414_);
  nor (_31416_, _27777_, _27788_);
  and (_31417_, _31416_, _31415_);
  and (_31418_, _31092_, _21861_);
  and (_31419_, _31090_, _20661_);
  nand (_31420_, _31419_, _31418_);
  nand (_31421_, _31420_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_31422_, _31421_, _31417_);
  or (_31423_, _31422_, _31413_);
  or (_31424_, _31423_, _31408_);
  and (_31425_, _31424_, _31400_);
  or (_31426_, _31425_, _31373_);
  not (_31427_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_31428_, _30175_, _31427_);
  nand (_31429_, _31428_, _31373_);
  or (_31430_, _31429_, _30186_);
  and (_31431_, _31430_, _31391_);
  and (_31432_, _31431_, _31426_);
  nor (_31433_, _31391_, _30947_);
  or (_31434_, _31433_, _31432_);
  and (_21373_, _31434_, _35796_);
  and (_31435_, _31373_, _30256_);
  nand (_31436_, _31435_, _28243_);
  and (_31437_, _31371_, _30890_);
  and (_31438_, _28347_, _28274_);
  and (_31439_, _31438_, _31437_);
  and (_31440_, _31439_, _30256_);
  or (_31441_, _31440_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_31442_, _31441_, _31391_);
  and (_31443_, _31442_, _31436_);
  nor (_31444_, _31391_, _30939_);
  or (_31445_, _31444_, _31443_);
  and (_21385_, _31445_, _35796_);
  not (_31446_, _31373_);
  or (_31447_, _31446_, _30331_);
  and (_31448_, _31447_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_31449_, _30330_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_31450_, _31449_, _30335_);
  and (_31451_, _31450_, _31373_);
  or (_31452_, _31451_, _31448_);
  and (_31453_, _31452_, _31391_);
  nor (_31454_, _31391_, _30932_);
  or (_31455_, _31454_, _31453_);
  and (_21397_, _31455_, _35796_);
  or (_31456_, _31446_, _30405_);
  and (_31457_, _31456_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_31458_, _31457_, _31386_);
  and (_31459_, _30412_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_31460_, _31459_, _30411_);
  and (_31461_, _31460_, _31373_);
  or (_31462_, _31461_, _31458_);
  nand (_31463_, _31386_, _30925_);
  and (_31464_, _31463_, _31462_);
  and (_21409_, _31464_, _35796_);
  or (_31465_, _30479_, _30224_);
  nand (_31466_, _31465_, _31373_);
  or (_31467_, _31466_, _30480_);
  nand (_31468_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_31469_, _25015_, _25895_);
  and (_31470_, _26618_, _26103_);
  nor (_31471_, _31470_, _31469_);
  nor (_31472_, _31471_, _31468_);
  or (_31473_, _31468_, _27460_);
  and (_31474_, _31473_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_31475_, _31474_, _31373_);
  or (_31476_, _31475_, _31472_);
  and (_31477_, _31476_, _31391_);
  and (_31478_, _31477_, _31467_);
  nor (_31479_, _31391_, _30918_);
  or (_31480_, _31479_, _31478_);
  and (_21421_, _31480_, _35796_);
  not (_31481_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_31482_, _31028_, _31481_);
  and (_31483_, _31482_, _31119_);
  not (_31484_, _31028_);
  and (_31485_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _15260_);
  and (_31486_, _31485_, _31484_);
  not (_31487_, _31486_);
  and (_31488_, _24916_, _24202_);
  and (_31489_, _24532_, _24378_);
  and (_31490_, _31489_, _24020_);
  and (_31491_, _31490_, _31488_);
  nand (_31492_, _31491_, _27711_);
  and (_31493_, _31492_, _31487_);
  nor (_31494_, _31493_, _27635_);
  and (_31495_, _24378_, _24202_);
  and (_31496_, _31495_, _28254_);
  and (_31497_, _31496_, _31438_);
  and (_31498_, _31497_, _28316_);
  and (_31499_, _31498_, _28243_);
  nor (_31500_, _31498_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_31501_, _31500_);
  not (_31502_, _31482_);
  and (_31503_, _31493_, _31502_);
  and (_31504_, _31503_, _31501_);
  not (_31505_, _31504_);
  nor (_31506_, _31505_, _31499_);
  nor (_31507_, _31506_, _31482_);
  not (_31508_, _31507_);
  nor (_31509_, _31508_, _31494_);
  nor (_31510_, _31509_, _31483_);
  and (_22201_, _31510_, _35796_);
  nor (_31511_, _31493_, _28739_);
  and (_31512_, _31497_, _24916_);
  and (_31513_, _31512_, _28243_);
  nor (_31514_, _31512_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not (_31515_, _31514_);
  and (_31516_, _31515_, _31503_);
  not (_31517_, _31516_);
  nor (_31518_, _31517_, _31513_);
  or (_31519_, _31518_, _31511_);
  and (_31520_, _31519_, _31502_);
  nor (_31521_, _31502_, _31157_);
  or (_31522_, _31521_, _31520_);
  and (_24064_, _31522_, _35796_);
  nor (_31523_, _31493_, _29380_);
  and (_31524_, _31497_, _29466_);
  and (_31525_, _31524_, _28243_);
  nor (_31526_, _31524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not (_31527_, _31526_);
  and (_31528_, _31527_, _31503_);
  not (_31529_, _31528_);
  nor (_31530_, _31529_, _31525_);
  or (_31531_, _31530_, _31523_);
  and (_31532_, _31531_, _31502_);
  nor (_31533_, _31502_, _31189_);
  or (_31534_, _31533_, _31532_);
  and (_24075_, _31534_, _35796_);
  nor (_31535_, _31493_, _30024_);
  and (_31536_, _31497_, _30175_);
  and (_31537_, _31536_, _28243_);
  nor (_31538_, _31536_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_31539_, _31538_);
  and (_31540_, _31539_, _31503_);
  not (_31541_, _31540_);
  nor (_31542_, _31541_, _31537_);
  or (_31543_, _31542_, _31535_);
  and (_31544_, _31543_, _31502_);
  nor (_31545_, _31502_, _31219_);
  or (_31546_, _31545_, _31544_);
  and (_24087_, _31546_, _35796_);
  nor (_31547_, _31502_, _31250_);
  nor (_31548_, _31493_, _30248_);
  not (_31549_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_31550_, _31497_, _31549_);
  not (_31551_, _31550_);
  and (_31552_, _31551_, _31493_);
  not (_31553_, _31552_);
  not (_31554_, _31497_);
  nor (_31555_, _30256_, _31549_);
  nor (_31556_, _31555_, _30258_);
  nor (_31557_, _31556_, _31554_);
  nor (_31558_, _31557_, _31553_);
  nor (_31559_, _31558_, _31482_);
  not (_31560_, _31559_);
  nor (_31561_, _31560_, _31548_);
  nor (_31562_, _31561_, _31547_);
  nor (_24099_, _31562_, rst);
  nor (_31563_, _31493_, _30319_);
  and (_31564_, _31497_, _30329_);
  and (_31565_, _31564_, _28243_);
  nor (_31566_, _31564_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_31567_, _31566_);
  and (_31568_, _31567_, _31503_);
  not (_31569_, _31568_);
  nor (_31570_, _31569_, _31565_);
  or (_31571_, _31570_, _31563_);
  and (_31572_, _31571_, _31502_);
  nor (_31573_, _31502_, _31281_);
  or (_31574_, _31573_, _31572_);
  and (_24111_, _31574_, _35796_);
  nor (_31575_, _31493_, _30396_);
  and (_31576_, _31497_, _30409_);
  and (_31577_, _31576_, _28243_);
  nor (_31578_, _31576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_31579_, _31578_);
  and (_31580_, _31579_, _31503_);
  not (_31581_, _31580_);
  nor (_31582_, _31581_, _31577_);
  or (_31583_, _31582_, _31575_);
  and (_31584_, _31583_, _31502_);
  nor (_31585_, _31502_, _31315_);
  or (_31586_, _31585_, _31584_);
  and (_24123_, _31586_, _35796_);
  nor (_31587_, _31493_, _30468_);
  and (_31588_, _31497_, _30479_);
  and (_31589_, _31588_, _28243_);
  nor (_31590_, _31588_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_31591_, _31590_);
  and (_31592_, _31591_, _31503_);
  not (_31593_, _31592_);
  nor (_31594_, _31593_, _31589_);
  or (_31595_, _31594_, _31587_);
  and (_31596_, _31595_, _31502_);
  nor (_31597_, _31502_, _31344_);
  or (_31598_, _31597_, _31596_);
  and (_24135_, _31598_, _35796_);
  and (_31599_, _30893_, _28316_);
  nand (_31600_, _31599_, _28243_);
  or (_31601_, _31599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_31602_, _31601_, _28347_);
  and (_31603_, _31602_, _31600_);
  and (_31604_, _30892_, _31488_);
  nand (_31605_, _31604_, _30907_);
  or (_31606_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_31607_, _31606_, _27711_);
  and (_31608_, _31607_, _31605_);
  not (_31609_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_31610_, _27700_, _31609_);
  or (_31611_, _31610_, rst);
  or (_31612_, _31611_, _31608_);
  or (_30648_, _31612_, _31603_);
  and (_31613_, _31371_, _30891_);
  and (_31614_, _31613_, _28316_);
  nand (_31615_, _31614_, _28243_);
  or (_31616_, _31614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_31617_, _31616_, _28347_);
  and (_31618_, _31617_, _31615_);
  and (_31619_, _31613_, _24916_);
  not (_31620_, _31619_);
  nor (_31621_, _31620_, _30907_);
  not (_31622_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_31623_, _31619_, _31622_);
  or (_31624_, _31623_, _31621_);
  and (_31625_, _31624_, _27711_);
  nor (_31626_, _27700_, _31622_);
  or (_31627_, _31626_, rst);
  or (_31628_, _31627_, _31625_);
  or (_30651_, _31628_, _31618_);
  and (_31629_, _24532_, _24009_);
  and (_31630_, _31629_, _31495_);
  and (_31631_, _31630_, _28274_);
  and (_31632_, _31631_, _28316_);
  nand (_31633_, _31632_, _28243_);
  or (_31634_, _31632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_31635_, _31634_, _28347_);
  and (_31636_, _31635_, _31633_);
  and (_31637_, _31631_, _24916_);
  not (_31638_, _31637_);
  nor (_31639_, _31638_, _30907_);
  not (_31640_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_31641_, _31637_, _31640_);
  or (_31642_, _31641_, _31639_);
  and (_31643_, _31642_, _27711_);
  nor (_31644_, _27700_, _31640_);
  or (_31645_, _31644_, rst);
  or (_31646_, _31645_, _31643_);
  or (_30654_, _31646_, _31636_);
  and (_31647_, _31629_, _28275_);
  not (_31648_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_31649_, _28316_, _31648_);
  or (_31650_, _31649_, _31374_);
  and (_31651_, _31650_, _31647_);
  nor (_31652_, _31647_, _31648_);
  or (_31653_, _31652_, _31651_);
  and (_31654_, _31653_, _28347_);
  and (_31655_, _30891_, _24938_);
  not (_31656_, _31655_);
  nor (_31657_, _31656_, _30907_);
  nor (_31658_, _31655_, _31648_);
  or (_31659_, _31658_, _31657_);
  and (_31660_, _31659_, _27711_);
  nor (_31661_, _27700_, _31648_);
  or (_31662_, _31661_, rst);
  or (_31663_, _31662_, _31660_);
  or (_30657_, _31663_, _31654_);
  or (_31664_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand (_31665_, _31604_, _28243_);
  and (_31666_, _31665_, _28347_);
  nand (_31667_, _31604_, _30962_);
  and (_31668_, _31667_, _27711_);
  or (_31669_, _31668_, _31666_);
  and (_31670_, _31669_, _31664_);
  not (_31671_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_31672_, _27700_, _31671_);
  or (_31673_, _31672_, rst);
  or (_33289_, _31673_, _31670_);
  or (_31674_, _30894_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_31675_, _31674_, _28347_);
  nand (_31676_, _30894_, _28243_);
  and (_31677_, _31676_, _31675_);
  nand (_31678_, _31604_, _30954_);
  or (_31679_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_31680_, _31679_, _27711_);
  and (_31681_, _31680_, _31678_);
  not (_31682_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_31683_, _27700_, _31682_);
  or (_31684_, _31683_, rst);
  or (_31685_, _31684_, _31681_);
  or (_33290_, _31685_, _31677_);
  not (_31686_, _30260_);
  nand (_31687_, _30893_, _31686_);
  and (_31688_, _31687_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_31689_, _24905_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_31690_, _31689_, _30186_);
  and (_31691_, _31690_, _30893_);
  or (_31692_, _31691_, _31688_);
  and (_31693_, _31692_, _28347_);
  nand (_31694_, _31604_, _30947_);
  or (_31695_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_31696_, _31695_, _27711_);
  and (_31697_, _31696_, _31694_);
  not (_31698_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_31699_, _27700_, _31698_);
  or (_31700_, _31699_, rst);
  or (_31701_, _31700_, _31697_);
  or (_33292_, _31701_, _31693_);
  nand (_31702_, _30893_, _24894_);
  and (_31703_, _31702_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_31704_, _31686_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_31705_, _31704_, _30258_);
  and (_31706_, _31705_, _30893_);
  or (_31707_, _31706_, _31703_);
  and (_31708_, _31707_, _28347_);
  nand (_31709_, _31604_, _30939_);
  or (_31710_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_31711_, _31710_, _27711_);
  and (_31712_, _31711_, _31709_);
  not (_31713_, _27700_);
  and (_31714_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_31715_, _31714_, rst);
  or (_31716_, _31715_, _31712_);
  or (_33294_, _31716_, _31708_);
  and (_31717_, _30893_, _30329_);
  nand (_31718_, _31717_, _28243_);
  or (_31719_, _31717_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_31720_, _31719_, _28347_);
  and (_31721_, _31720_, _31718_);
  nand (_31722_, _31604_, _30932_);
  or (_31723_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_31724_, _31723_, _27711_);
  and (_31725_, _31724_, _31722_);
  and (_31726_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_31727_, _31726_, rst);
  or (_31728_, _31727_, _31725_);
  or (_33296_, _31728_, _31721_);
  and (_31729_, _30893_, _30409_);
  nand (_31730_, _31729_, _28243_);
  or (_31731_, _31729_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_31732_, _31731_, _28347_);
  and (_31733_, _31732_, _31730_);
  nand (_31734_, _31604_, _30925_);
  or (_31735_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_31736_, _31735_, _27711_);
  and (_31737_, _31736_, _31734_);
  and (_31738_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_31739_, _31738_, rst);
  or (_31740_, _31739_, _31737_);
  or (_33298_, _31740_, _31733_);
  nand (_31741_, _30893_, _30476_);
  and (_31742_, _31741_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  not (_31743_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_31744_, _28306_, _31743_);
  or (_31745_, _31744_, _30480_);
  and (_31746_, _31745_, _30893_);
  or (_31747_, _31746_, _31742_);
  and (_31748_, _31747_, _28347_);
  nand (_31749_, _31604_, _30918_);
  or (_31750_, _31604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_31751_, _31750_, _27711_);
  and (_31752_, _31751_, _31749_);
  nor (_31753_, _27700_, _31743_);
  or (_31754_, _31753_, rst);
  or (_31755_, _31754_, _31752_);
  or (_33300_, _31755_, _31748_);
  nand (_31756_, _31619_, _28243_);
  or (_31757_, _31619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_31758_, _31757_, _28347_);
  and (_31759_, _31758_, _31756_);
  and (_31760_, _31619_, _30963_);
  not (_31761_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_31762_, _31619_, _31761_);
  or (_31763_, _31762_, _31760_);
  and (_31764_, _31763_, _27711_);
  nor (_31765_, _27700_, _31761_);
  or (_31766_, _31765_, rst);
  or (_31767_, _31766_, _31764_);
  or (_33302_, _31767_, _31759_);
  and (_31768_, _31613_, _29466_);
  nand (_31769_, _31768_, _28243_);
  or (_31770_, _31768_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_31771_, _31770_, _28347_);
  and (_31772_, _31771_, _31769_);
  nor (_31773_, _31620_, _30954_);
  not (_31774_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_31775_, _31619_, _31774_);
  or (_31776_, _31775_, _31773_);
  and (_31777_, _31776_, _27711_);
  nor (_31778_, _27700_, _31774_);
  or (_31779_, _31778_, rst);
  or (_31780_, _31779_, _31777_);
  or (_33303_, _31780_, _31772_);
  and (_31781_, _31613_, _30175_);
  nand (_31782_, _31781_, _28243_);
  or (_31783_, _31781_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_31784_, _31783_, _28347_);
  and (_31785_, _31784_, _31782_);
  nor (_31786_, _31620_, _30947_);
  not (_31787_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_31788_, _31619_, _31787_);
  or (_31789_, _31788_, _31786_);
  and (_31790_, _31789_, _27711_);
  nor (_31791_, _27700_, _31787_);
  or (_31792_, _31791_, rst);
  or (_31793_, _31792_, _31790_);
  or (_33305_, _31793_, _31785_);
  and (_31794_, _31613_, _30256_);
  nand (_31795_, _31794_, _28243_);
  or (_31796_, _31794_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_31797_, _31796_, _28347_);
  and (_31798_, _31797_, _31795_);
  nor (_31799_, _31620_, _30939_);
  and (_31800_, _31620_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_31801_, _31800_, _31799_);
  and (_31802_, _31801_, _27711_);
  and (_31803_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_31804_, _31803_, rst);
  or (_31805_, _31804_, _31802_);
  or (_33307_, _31805_, _31798_);
  and (_31806_, _31613_, _30329_);
  nand (_31807_, _31806_, _28243_);
  or (_31808_, _31806_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_31809_, _31808_, _28347_);
  and (_31810_, _31809_, _31807_);
  nor (_31811_, _31620_, _30932_);
  and (_31812_, _31620_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_31813_, _31812_, _31811_);
  and (_31814_, _31813_, _27711_);
  and (_31815_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_31816_, _31815_, rst);
  or (_31817_, _31816_, _31814_);
  or (_33309_, _31817_, _31810_);
  and (_31818_, _31613_, _30409_);
  nand (_31819_, _31818_, _28243_);
  or (_31820_, _31818_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_31821_, _31820_, _28347_);
  and (_31822_, _31821_, _31819_);
  nor (_31823_, _31620_, _30925_);
  and (_31824_, _31620_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_31825_, _31824_, _31823_);
  and (_31826_, _31825_, _27711_);
  and (_31827_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_31828_, _31827_, rst);
  or (_31829_, _31828_, _31826_);
  or (_33311_, _31829_, _31822_);
  and (_31830_, _31613_, _30479_);
  nand (_31831_, _31830_, _28243_);
  or (_31832_, _31830_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_31833_, _31832_, _28347_);
  and (_31834_, _31833_, _31831_);
  nor (_31835_, _31620_, _30918_);
  not (_31836_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_31837_, _31619_, _31836_);
  or (_31838_, _31837_, _31835_);
  and (_31839_, _31838_, _27711_);
  nor (_31840_, _27700_, _31836_);
  or (_31841_, _31840_, rst);
  or (_31842_, _31841_, _31839_);
  or (_33313_, _31842_, _31834_);
  nand (_31843_, _31637_, _28243_);
  or (_31844_, _31637_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_31845_, _31844_, _28347_);
  and (_31846_, _31845_, _31843_);
  and (_31847_, _31637_, _30963_);
  not (_31848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_31849_, _31637_, _31848_);
  or (_31850_, _31849_, _31847_);
  and (_31851_, _31850_, _27711_);
  nor (_31852_, _27700_, _31848_);
  or (_31853_, _31852_, rst);
  or (_31854_, _31853_, _31851_);
  or (_33314_, _31854_, _31846_);
  and (_31855_, _31631_, _29466_);
  nand (_31856_, _31855_, _28243_);
  or (_31857_, _31855_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_31858_, _31857_, _28347_);
  and (_31859_, _31858_, _31856_);
  nor (_31860_, _31638_, _30954_);
  not (_31861_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_31862_, _31637_, _31861_);
  or (_31863_, _31862_, _31860_);
  and (_31864_, _31863_, _27711_);
  nor (_31865_, _27700_, _31861_);
  or (_31866_, _31865_, rst);
  or (_31867_, _31866_, _31864_);
  or (_33316_, _31867_, _31859_);
  and (_31868_, _31631_, _30175_);
  nand (_31869_, _31868_, _28243_);
  or (_31870_, _31868_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_31871_, _31870_, _28347_);
  and (_31872_, _31871_, _31869_);
  nor (_31873_, _31638_, _30947_);
  not (_31874_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_31875_, _31637_, _31874_);
  or (_31876_, _31875_, _31873_);
  and (_31877_, _31876_, _27711_);
  nor (_31878_, _27700_, _31874_);
  or (_31879_, _31878_, rst);
  or (_31880_, _31879_, _31877_);
  or (_33318_, _31880_, _31872_);
  and (_31881_, _31631_, _30256_);
  nand (_31882_, _31881_, _28243_);
  or (_31883_, _31881_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_31884_, _31883_, _28347_);
  and (_31885_, _31884_, _31882_);
  nor (_31886_, _31638_, _30939_);
  and (_31887_, _31638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_31888_, _31887_, _31886_);
  and (_31889_, _31888_, _27711_);
  and (_31890_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_31891_, _31890_, rst);
  or (_31892_, _31891_, _31889_);
  or (_33320_, _31892_, _31885_);
  and (_31893_, _31631_, _30329_);
  nand (_31894_, _31893_, _28243_);
  or (_31895_, _31893_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_31896_, _31895_, _28347_);
  and (_31897_, _31896_, _31894_);
  nor (_31898_, _31638_, _30932_);
  and (_31899_, _31638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_31900_, _31899_, _31898_);
  and (_31901_, _31900_, _27711_);
  and (_31902_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_31903_, _31902_, rst);
  or (_31904_, _31903_, _31901_);
  or (_33322_, _31904_, _31897_);
  and (_31905_, _31631_, _30409_);
  nand (_31906_, _31905_, _28243_);
  or (_31907_, _31905_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_31908_, _31907_, _28347_);
  and (_31909_, _31908_, _31906_);
  nor (_31910_, _31638_, _30925_);
  and (_31911_, _31638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_31912_, _31911_, _31910_);
  and (_31913_, _31912_, _27711_);
  and (_31914_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_31915_, _31914_, rst);
  or (_31916_, _31915_, _31913_);
  or (_33324_, _31916_, _31909_);
  and (_31917_, _31631_, _30479_);
  nand (_31918_, _31917_, _28243_);
  or (_31919_, _31917_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_31920_, _31919_, _28347_);
  and (_31921_, _31920_, _31918_);
  nor (_31922_, _31638_, _30918_);
  not (_31923_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_31924_, _31637_, _31923_);
  or (_31925_, _31924_, _31922_);
  and (_31926_, _31925_, _27711_);
  nor (_31927_, _27700_, _31923_);
  or (_31928_, _31927_, rst);
  or (_31929_, _31928_, _31926_);
  or (_33325_, _31929_, _31921_);
  nand (_31930_, _28243_, _24916_);
  or (_31931_, _24916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_31932_, _31931_, _31647_);
  and (_31933_, _31932_, _31930_);
  not (_31934_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_31935_, _31647_, _31934_);
  or (_31936_, _31935_, _31933_);
  and (_31937_, _31936_, _28347_);
  nor (_31938_, _31656_, _30962_);
  nor (_31939_, _31655_, _31934_);
  or (_31940_, _31939_, _31938_);
  and (_31941_, _31940_, _27711_);
  nor (_31942_, _27700_, _31934_);
  or (_31943_, _31942_, rst);
  or (_31944_, _31943_, _31941_);
  or (_33327_, _31944_, _31937_);
  nand (_31945_, _29466_, _28243_);
  or (_31946_, _29466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_31947_, _31946_, _31647_);
  and (_31948_, _31947_, _31945_);
  not (_31949_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_31950_, _31647_, _31949_);
  or (_31951_, _31950_, _31948_);
  and (_31952_, _31951_, _28347_);
  nor (_31953_, _31656_, _30954_);
  nor (_31954_, _31655_, _31949_);
  or (_31955_, _31954_, _31953_);
  and (_31956_, _31955_, _27711_);
  nor (_31957_, _27700_, _31949_);
  or (_31958_, _31957_, rst);
  or (_31959_, _31958_, _31956_);
  or (_33329_, _31959_, _31952_);
  not (_31960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_31961_, _30175_, _31960_);
  or (_31962_, _31961_, _30186_);
  and (_31963_, _31962_, _31647_);
  nor (_31964_, _31647_, _31960_);
  or (_31965_, _31964_, _31963_);
  and (_31966_, _31965_, _28347_);
  nor (_31967_, _31656_, _30947_);
  nor (_31968_, _31655_, _31960_);
  or (_31969_, _31968_, _31967_);
  and (_31970_, _31969_, _27711_);
  nor (_31971_, _27700_, _31960_);
  or (_31972_, _31971_, rst);
  or (_31973_, _31972_, _31970_);
  or (_33331_, _31973_, _31966_);
  and (_31974_, _30257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31975_, _31974_, _30258_);
  and (_31976_, _31975_, _31647_);
  not (_31977_, _31647_);
  and (_31978_, _31977_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31979_, _31978_, _31976_);
  and (_31980_, _31979_, _28347_);
  nor (_31981_, _31656_, _30939_);
  and (_31982_, _31656_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31983_, _31982_, _31981_);
  and (_31984_, _31983_, _27711_);
  and (_31985_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31986_, _31985_, rst);
  or (_31987_, _31986_, _31984_);
  or (_33333_, _31987_, _31980_);
  and (_31988_, _30334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31989_, _31988_, _30335_);
  and (_31990_, _31989_, _31647_);
  and (_31991_, _31977_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31992_, _31991_, _31990_);
  and (_31993_, _31992_, _28347_);
  nor (_31994_, _31656_, _30932_);
  and (_31995_, _31656_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31996_, _31995_, _31994_);
  and (_31997_, _31996_, _27711_);
  and (_31998_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31999_, _31998_, rst);
  or (_32000_, _31999_, _31997_);
  or (_33335_, _32000_, _31993_);
  and (_32001_, _30410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_32002_, _32001_, _30411_);
  and (_32003_, _32002_, _31647_);
  and (_32004_, _31977_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_32005_, _32004_, _32003_);
  and (_32006_, _32005_, _28347_);
  nor (_32007_, _31656_, _30925_);
  and (_32008_, _31656_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_32009_, _32008_, _32007_);
  and (_32010_, _32009_, _27711_);
  and (_32011_, _31713_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_32012_, _32011_, rst);
  or (_32013_, _32012_, _32010_);
  or (_33336_, _32013_, _32006_);
  not (_32014_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_32015_, _30479_, _32014_);
  or (_32016_, _32015_, _30480_);
  and (_32017_, _32016_, _31647_);
  nor (_32018_, _31647_, _32014_);
  or (_32019_, _32018_, _32017_);
  and (_32020_, _32019_, _28347_);
  nor (_32021_, _31656_, _30918_);
  nor (_32022_, _31655_, _32014_);
  or (_32023_, _32022_, _32021_);
  and (_32024_, _32023_, _27711_);
  nor (_32025_, _27700_, _32014_);
  or (_32026_, _32025_, rst);
  or (_32027_, _32026_, _32024_);
  or (_33338_, _32027_, _32020_);
  and (_32028_, _27678_, _23855_);
  not (_32029_, _32028_);
  and (_32030_, _23877_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32031_, _32030_, _24213_);
  nor (_32032_, _24653_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_32033_, _32032_, _32031_);
  not (_32034_, _32033_);
  not (_32035_, _30886_);
  and (_32036_, _32035_, _30850_);
  and (_32037_, _32036_, _30745_);
  nor (_32038_, _30628_, _24653_);
  and (_32039_, _30628_, _24653_);
  nor (_32040_, _32039_, _32038_);
  not (_32041_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_32042_, _24905_, _32041_);
  and (_32043_, _32042_, _32028_);
  not (_32044_, _32043_);
  nor (_32045_, _32044_, _32040_);
  not (_32046_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_32047_, _31386_, _32046_);
  nor (_32048_, _32047_, _31444_);
  nor (_32049_, _32048_, _24213_);
  and (_32050_, _32048_, _24213_);
  nor (_32051_, _32050_, _32049_);
  and (_32052_, _32051_, _32045_);
  not (_32053_, _17075_);
  and (_32054_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25389_);
  not (_32055_, _25400_);
  and (_32056_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_32057_, _32056_, _32055_);
  nor (_32058_, _32057_, _32054_);
  nor (_32059_, _32058_, _32053_);
  and (_32060_, _32056_, _25400_);
  and (_32061_, _32060_, _28827_);
  nor (_32062_, _30907_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32063_, _32062_, _32061_);
  nor (_32064_, _32063_, _32059_);
  nor (_32065_, _32030_, _24213_);
  and (_32066_, _32030_, _24009_);
  nor (_32067_, _32066_, _32065_);
  and (_32068_, _32067_, _32048_);
  not (_32069_, _32068_);
  nor (_32070_, _32067_, _32048_);
  nor (_32071_, _32033_, _30628_);
  and (_32072_, _32033_, _30628_);
  nor (_32073_, _32072_, _32071_);
  not (_32074_, _32073_);
  and (_32075_, _32030_, _24532_);
  nor (_32076_, _24894_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_32077_, _32076_, _32075_);
  not (_32078_, _24378_);
  and (_32079_, _32030_, _32078_);
  nor (_32080_, _24773_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_32081_, _32080_, _32079_);
  and (_32082_, _32081_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_32083_, _32082_, _32077_);
  and (_32084_, _32083_, _32074_);
  not (_32085_, _32084_);
  nor (_32086_, _32085_, _32070_);
  and (_32087_, _32086_, _32069_);
  and (_32088_, _32087_, _32064_);
  not (_32089_, _32087_);
  and (_32090_, _32048_, _30629_);
  and (_32091_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_32092_, _32048_, _30629_);
  and (_32093_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_32094_, _32093_, _32091_);
  nor (_32095_, _32048_, _30628_);
  and (_32096_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_32097_, _32048_, _30628_);
  and (_32098_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_32099_, _32098_, _32096_);
  and (_32100_, _32099_, _32094_);
  and (_32101_, _32100_, _32089_);
  nor (_32102_, _32101_, _32088_);
  nor (_32103_, _32102_, _32052_);
  and (_32104_, _32052_, _30907_);
  nor (_32105_, _32104_, _32103_);
  and (_32106_, _32105_, _32037_);
  not (_32107_, _32106_);
  not (_32108_, _30745_);
  nor (_32109_, _32035_, _30850_);
  not (_32110_, _30494_);
  and (_32111_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_32112_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_32113_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_32114_, _32113_, _32112_);
  and (_32115_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_32116_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_32117_, _32116_, _32115_);
  and (_32118_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_32119_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_32120_, _32119_, _32118_);
  and (_32121_, _32120_, _32117_);
  and (_32122_, _32121_, _32114_);
  and (_32123_, _30632_, _30494_);
  not (_32124_, _32123_);
  nor (_32125_, _32124_, _32122_);
  nor (_32126_, _32125_, _32111_);
  not (_32127_, _32126_);
  and (_32128_, _32127_, _32109_);
  nor (_32129_, _32128_, _32108_);
  not (_32130_, _30980_);
  nand (_32131_, _32130_, _30887_);
  and (_32132_, _32131_, _32129_);
  and (_32133_, _32132_, _32107_);
  and (_32134_, _30804_, _30532_);
  nor (_32135_, _32134_, _30811_);
  and (_32136_, _30807_, _30735_);
  nor (_32137_, _32136_, _30760_);
  and (_32138_, _32137_, _30828_);
  and (_32139_, _32138_, _32135_);
  not (_32140_, _30748_);
  and (_32141_, _30810_, _32140_);
  and (_32142_, _32141_, _30783_);
  and (_32143_, _32142_, _32139_);
  nor (_32144_, _32143_, _30490_);
  and (_32145_, _30735_, _30778_);
  nor (_32146_, _30841_, _32145_);
  nor (_32147_, _30843_, _32146_);
  nor (_32148_, _32147_, _32144_);
  not (_32149_, _32148_);
  and (_32150_, _32149_, _32133_);
  not (_32151_, _30939_);
  and (_32152_, _32052_, _32151_);
  and (_32153_, _32054_, _25400_);
  and (_32154_, _32153_, _28827_);
  nor (_32155_, _30939_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32156_, _32054_, _32055_);
  or (_32157_, _32156_, _32056_);
  and (_32158_, _32157_, _16589_);
  or (_32159_, _32158_, _32155_);
  or (_32160_, _32159_, _32154_);
  or (_32161_, _32160_, _32089_);
  not (_32162_, _32052_);
  and (_32163_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_32164_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_32165_, _32164_, _32163_);
  and (_32166_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_32167_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_32168_, _32167_, _32166_);
  or (_32169_, _32168_, _32165_);
  or (_32170_, _32169_, _32087_);
  and (_32171_, _32170_, _32162_);
  and (_32172_, _32171_, _32161_);
  or (_32173_, _32172_, _32152_);
  and (_32174_, _32173_, _32037_);
  not (_32175_, _32174_);
  not (_32176_, _31006_);
  and (_32177_, _32176_, _30888_);
  not (_32178_, _32177_);
  not (_32179_, _32048_);
  and (_32180_, _30745_, _30886_);
  and (_32181_, _32180_, _30850_);
  and (_32182_, _32181_, _32179_);
  and (_32183_, _32109_, _30745_);
  and (_32184_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_32185_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_32186_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_32187_, _32186_, _32185_);
  and (_32188_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_32189_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_32190_, _32189_, _32188_);
  and (_32191_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_32192_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_32193_, _32192_, _32191_);
  and (_32194_, _32193_, _32190_);
  and (_32195_, _32194_, _32187_);
  nor (_32196_, _32195_, _32124_);
  nor (_32197_, _32196_, _32184_);
  not (_32198_, _32197_);
  and (_32199_, _32198_, _32183_);
  nor (_32200_, _32199_, _32182_);
  and (_32201_, _32200_, _32178_);
  and (_32202_, _32201_, _32175_);
  not (_32203_, _32202_);
  and (_32204_, _32203_, _32150_);
  and (_32205_, _32054_, _25443_);
  and (_32206_, _32205_, _28243_);
  not (_32207_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32208_, _30962_, _32207_);
  nor (_32209_, _15934_, _32207_);
  nor (_32210_, _32209_, _32208_);
  nor (_32211_, _32210_, _32205_);
  nor (_32212_, _32211_, _32206_);
  nor (_32213_, _32212_, _32089_);
  and (_32214_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_32215_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_32216_, _32215_, _32214_);
  and (_32217_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_32218_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_32219_, _32218_, _32217_);
  and (_32220_, _32219_, _32216_);
  and (_32221_, _32220_, _32089_);
  nor (_32222_, _32221_, _32213_);
  nor (_32223_, _32222_, _32052_);
  and (_32224_, _32052_, _30962_);
  nor (_32225_, _32224_, _32223_);
  and (_32226_, _32225_, _32037_);
  not (_32227_, _32226_);
  not (_32228_, _30988_);
  and (_32229_, _32228_, _30888_);
  not (_32230_, _32229_);
  and (_32231_, _32181_, _30629_);
  and (_32232_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_32233_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_32234_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_32235_, _32234_, _32233_);
  and (_32236_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_32237_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_32238_, _32237_, _32236_);
  and (_32239_, _32238_, _32235_);
  and (_32240_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_32241_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_32242_, _32241_, _32240_);
  and (_32243_, _32242_, _32239_);
  nor (_32244_, _32243_, _32124_);
  nor (_32245_, _32244_, _32232_);
  not (_32246_, _32245_);
  and (_32247_, _32246_, _32183_);
  nor (_32248_, _32247_, _32231_);
  and (_32249_, _32248_, _32230_);
  and (_32250_, _32249_, _32227_);
  nor (_32251_, _32250_, _32149_);
  nor (_32252_, _32251_, _32204_);
  and (_32253_, _32252_, _32034_);
  nor (_32254_, _32253_, _32029_);
  not (_32255_, _32077_);
  not (_32256_, _32037_);
  nor (_32257_, _32162_, _30925_);
  and (_32258_, _25477_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_32259_, _32258_);
  and (_32260_, _16737_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32261_, _32260_, _32259_);
  and (_32262_, _32056_, _25477_);
  and (_32263_, _32262_, _28827_);
  nor (_32264_, _30925_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32265_, _32264_, _32263_);
  nor (_32266_, _32265_, _32261_);
  and (_32267_, _32266_, _32087_);
  and (_32268_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_32269_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_32270_, _32269_, _32268_);
  and (_32271_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_32272_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_32273_, _32272_, _32271_);
  and (_32274_, _32273_, _32270_);
  and (_32275_, _32274_, _32089_);
  nor (_32276_, _32275_, _32052_);
  not (_32277_, _32276_);
  nor (_32278_, _32277_, _32267_);
  nor (_32279_, _32278_, _32257_);
  nor (_32280_, _32279_, _32256_);
  not (_32281_, _32280_);
  not (_32282_, _31018_);
  and (_32283_, _32282_, _30888_);
  and (_32284_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_32285_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_32286_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_32287_, _32286_, _32285_);
  and (_32288_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_32289_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_32290_, _32289_, _32288_);
  and (_32291_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_32292_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_32293_, _32292_, _32291_);
  and (_32294_, _32293_, _32290_);
  and (_32295_, _32294_, _32287_);
  nor (_32296_, _32295_, _32124_);
  nor (_32297_, _32296_, _32284_);
  not (_32298_, _32297_);
  and (_32299_, _32298_, _32183_);
  not (_32300_, _32109_);
  nor (_32301_, _32036_, _30745_);
  and (_32302_, _32301_, _32300_);
  or (_32303_, _32302_, _32299_);
  nor (_32304_, _32303_, _32283_);
  and (_32305_, _32304_, _32281_);
  not (_32306_, _32305_);
  and (_32307_, _32306_, _32150_);
  nor (_32308_, _32162_, _30947_);
  nand (_32309_, _32054_, _25510_);
  nor (_32310_, _32309_, _28243_);
  nor (_32311_, _30947_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_32312_, _32153_, _32056_);
  nand (_32313_, _32054_, _25466_);
  nand (_32314_, _32313_, _32312_);
  and (_32315_, _32314_, _15575_);
  or (_32316_, _32315_, _32311_);
  or (_32317_, _32316_, _32310_);
  or (_32318_, _32317_, _32089_);
  and (_32319_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_32320_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_32321_, _32320_, _32319_);
  and (_32322_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_32323_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_32324_, _32323_, _32322_);
  or (_32325_, _32324_, _32321_);
  or (_32326_, _32325_, _32087_);
  and (_32327_, _32326_, _32162_);
  and (_32328_, _32327_, _32318_);
  or (_32329_, _32328_, _32308_);
  and (_32330_, _32329_, _32037_);
  not (_32331_, _32330_);
  not (_32332_, _31000_);
  and (_32333_, _32332_, _30888_);
  not (_32334_, _32333_);
  and (_32335_, _32181_, _30721_);
  and (_32336_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_32337_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_32338_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_32339_, _32338_, _32337_);
  and (_32340_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_32341_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_32342_, _32341_, _32340_);
  and (_32343_, _32342_, _32339_);
  and (_32344_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_32345_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_32346_, _32345_, _32344_);
  and (_32347_, _32346_, _32343_);
  nor (_32348_, _32347_, _32124_);
  nor (_32349_, _32348_, _32336_);
  not (_32350_, _32349_);
  and (_32351_, _32350_, _32183_);
  nor (_32352_, _32351_, _32335_);
  and (_32353_, _32352_, _32334_);
  and (_32354_, _32353_, _32331_);
  nor (_32355_, _32354_, _32149_);
  nor (_32356_, _32355_, _32307_);
  and (_32357_, _32356_, _32255_);
  nor (_32358_, _32252_, _32034_);
  nor (_32359_, _32358_, _32357_);
  and (_32360_, _32359_, _32254_);
  not (_32361_, _30932_);
  and (_32362_, _32052_, _32361_);
  nand (_32363_, _32056_, _25443_);
  nor (_32364_, _32363_, _28243_);
  nor (_32365_, _30932_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_32366_, _25443_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_32367_, _15770_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32368_, _32367_, _32366_);
  or (_32369_, _32368_, _32365_);
  or (_32370_, _32369_, _32364_);
  or (_32371_, _32370_, _32089_);
  and (_32372_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_32373_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_32374_, _32373_, _32372_);
  and (_32375_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_32376_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_32377_, _32376_, _32375_);
  or (_32378_, _32377_, _32374_);
  or (_32379_, _32378_, _32087_);
  and (_32380_, _32379_, _32162_);
  and (_32381_, _32380_, _32371_);
  or (_32382_, _32381_, _32362_);
  and (_32383_, _32382_, _32037_);
  not (_32384_, _32383_);
  not (_32385_, _31012_);
  and (_32386_, _32385_, _30888_);
  and (_32387_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_32388_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_32389_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_32390_, _32389_, _32388_);
  and (_32391_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_32392_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_32393_, _32392_, _32391_);
  and (_32394_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_32395_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_32396_, _32395_, _32394_);
  and (_32397_, _32396_, _32393_);
  and (_32398_, _32397_, _32390_);
  nor (_32399_, _32398_, _32124_);
  nor (_32400_, _32399_, _32387_);
  not (_32401_, _32400_);
  and (_32402_, _32401_, _32183_);
  nor (_32403_, _32402_, _32386_);
  and (_32404_, _32108_, _30886_);
  not (_32405_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_32406_, _31386_, _32405_);
  nor (_32407_, _32406_, _31454_);
  not (_32408_, _32407_);
  and (_32409_, _32408_, _32181_);
  or (_32410_, _32409_, _32404_);
  not (_32411_, _32410_);
  and (_32412_, _32411_, _32403_);
  and (_32413_, _32412_, _32384_);
  not (_32414_, _32413_);
  and (_32415_, _32414_, _32150_);
  and (_32416_, _32036_, _32108_);
  not (_32417_, _30994_);
  and (_32418_, _32417_, _30888_);
  nor (_32419_, _32418_, _32416_);
  and (_32420_, _32181_, _30656_);
  not (_32421_, _16901_);
  and (_32422_, _32054_, _25499_);
  not (_32423_, _32422_);
  and (_32424_, _32312_, _32423_);
  nor (_32425_, _32424_, _32421_);
  and (_32426_, _32054_, _25477_);
  and (_32427_, _32426_, _28827_);
  nor (_32428_, _30954_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32429_, _32428_, _32427_);
  nor (_32430_, _32429_, _32425_);
  and (_32431_, _32430_, _32087_);
  and (_32432_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_32433_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_32434_, _32433_, _32432_);
  and (_32435_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_32436_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_32437_, _32436_, _32435_);
  and (_32438_, _32437_, _32434_);
  and (_32439_, _32438_, _32089_);
  nor (_32440_, _32439_, _32431_);
  nor (_32441_, _32440_, _32052_);
  and (_32442_, _32052_, _30954_);
  nor (_32443_, _32442_, _32441_);
  and (_32444_, _32443_, _32037_);
  and (_32445_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_32446_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_32447_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_32448_, _32447_, _32446_);
  and (_32449_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_32450_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_32451_, _32450_, _32449_);
  and (_32452_, _32451_, _32448_);
  and (_32453_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_32454_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_32455_, _32454_, _32453_);
  and (_32456_, _32455_, _32452_);
  nor (_32457_, _32456_, _32124_);
  nor (_32458_, _32457_, _32445_);
  not (_32459_, _32458_);
  and (_32460_, _32459_, _32183_);
  or (_32461_, _32460_, _32444_);
  nor (_32462_, _32461_, _32420_);
  and (_32463_, _32462_, _32419_);
  nor (_32464_, _32463_, _32149_);
  nor (_32465_, _32464_, _32415_);
  nand (_32466_, _32465_, _32081_);
  or (_32467_, _32465_, _32081_);
  and (_32468_, _32467_, _32466_);
  not (_32469_, _32468_);
  nor (_32470_, _32356_, _32255_);
  not (_32471_, _32470_);
  not (_32472_, _32067_);
  nor (_32473_, _32203_, _32150_);
  not (_32474_, _30918_);
  and (_32475_, _32052_, _32474_);
  and (_32476_, _25510_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_32477_, _32476_);
  and (_32478_, _16108_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32479_, _32478_, _32477_);
  and (_32480_, _32056_, _25510_);
  and (_32481_, _32480_, _28827_);
  nor (_32482_, _30918_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32483_, _32482_, _32481_);
  nor (_32484_, _32483_, _32479_);
  and (_32485_, _32484_, _32087_);
  and (_32486_, _32092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_32487_, _32090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_32488_, _32487_, _32486_);
  and (_32489_, _32095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_32490_, _32097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_32491_, _32490_, _32489_);
  and (_32492_, _32491_, _32488_);
  and (_32493_, _32492_, _32089_);
  nor (_32494_, _32493_, _32052_);
  not (_32495_, _32494_);
  nor (_32496_, _32495_, _32485_);
  nor (_32497_, _32496_, _32475_);
  nor (_32498_, _32497_, _32256_);
  not (_32499_, _31024_);
  and (_32500_, _32499_, _30888_);
  and (_32501_, _32110_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_32502_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_32503_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_32504_, _32503_, _32502_);
  and (_32505_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_32506_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_32507_, _32506_, _32505_);
  and (_32508_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_32509_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_32510_, _32509_, _32508_);
  and (_32511_, _32510_, _32507_);
  and (_32512_, _32511_, _32504_);
  nor (_32513_, _32512_, _32124_);
  nor (_32514_, _32513_, _32501_);
  not (_32515_, _32514_);
  and (_32516_, _32515_, _32109_);
  nor (_32517_, _32516_, _32301_);
  not (_32518_, _32517_);
  nor (_32519_, _32518_, _32500_);
  not (_32520_, _32519_);
  nor (_32521_, _32520_, _32498_);
  and (_32522_, _32521_, _32150_);
  nor (_32523_, _32522_, _32473_);
  nor (_32524_, _32523_, _32472_);
  and (_32525_, _32523_, _32472_);
  nor (_32526_, _32525_, _32524_);
  and (_32527_, _32526_, _32471_);
  and (_32528_, _32527_, _32469_);
  and (_32529_, _32528_, _32360_);
  not (_32530_, _32356_);
  and (_32531_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_32532_, _32252_);
  and (_32533_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_32534_, _32533_, _32531_);
  and (_32535_, _32534_, _32465_);
  not (_32536_, _32465_);
  not (_32537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_32538_, _32252_, _32537_);
  and (_32539_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_32540_, _32539_, _32538_);
  and (_32541_, _32540_, _32536_);
  or (_32542_, _32541_, _32535_);
  or (_32543_, _32542_, _32530_);
  not (_32544_, _32523_);
  and (_32545_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_32546_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_32547_, _32546_, _32545_);
  and (_32548_, _32547_, _32465_);
  not (_32549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_32550_, _32252_, _32549_);
  and (_32551_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_32552_, _32551_, _32550_);
  and (_32553_, _32552_, _32536_);
  or (_32554_, _32553_, _32548_);
  or (_32555_, _32554_, _32356_);
  and (_32556_, _32555_, _32544_);
  and (_32557_, _32556_, _32543_);
  or (_32558_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_32559_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_32560_, _32559_, _32558_);
  and (_32561_, _32560_, _32465_);
  or (_32562_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_32563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_32564_, _32252_, _32563_);
  and (_32565_, _32564_, _32562_);
  and (_32566_, _32565_, _32536_);
  or (_32567_, _32566_, _32561_);
  or (_32568_, _32567_, _32530_);
  or (_32569_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_32570_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_32571_, _32570_, _32569_);
  and (_32572_, _32571_, _32465_);
  or (_32573_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_32574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_32575_, _32252_, _32574_);
  and (_32576_, _32575_, _32573_);
  and (_32577_, _32576_, _32536_);
  or (_32578_, _32577_, _32572_);
  or (_32579_, _32578_, _32356_);
  and (_32580_, _32579_, _32523_);
  and (_32581_, _32580_, _32568_);
  or (_32582_, _32581_, _32557_);
  or (_32583_, _32582_, _32529_);
  not (_32584_, _32529_);
  or (_32585_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_32586_, _32585_, _35796_);
  and (_33414_, _32586_, _32583_);
  nor (_32587_, _32081_, _32029_);
  nor (_32588_, _32033_, _32029_);
  and (_32589_, _32588_, _32587_);
  nor (_32590_, _32077_, _32029_);
  and (_32591_, _32067_, _32028_);
  and (_32592_, _32591_, _32590_);
  and (_32593_, _32592_, _32589_);
  nor (_32594_, _32064_, _32029_);
  and (_32595_, _32594_, _32593_);
  not (_32596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_32597_, _32593_, _32596_);
  or (_33424_, _32597_, _32595_);
  nor (_32598_, _32588_, _32587_);
  nor (_32599_, _32591_, _32590_);
  and (_32600_, _32599_, _32028_);
  and (_32601_, _32600_, _32598_);
  and (_32602_, _32212_, _32028_);
  and (_32603_, _32602_, _32601_);
  not (_32604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_32605_, _32601_, _32604_);
  or (_33667_, _32605_, _32603_);
  nor (_32606_, _32430_, _32029_);
  and (_32607_, _32606_, _32601_);
  not (_32608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_32609_, _32601_, _32608_);
  or (_33672_, _32609_, _32607_);
  and (_32610_, _32317_, _32028_);
  and (_32611_, _32610_, _32601_);
  not (_32612_, _32601_);
  and (_32613_, _32612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_33677_, _32613_, _32611_);
  and (_32614_, _32160_, _32028_);
  and (_32615_, _32614_, _32601_);
  and (_32616_, _32612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_33682_, _32616_, _32615_);
  and (_32617_, _32370_, _32028_);
  and (_32618_, _32617_, _32601_);
  and (_32619_, _32612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_33687_, _32619_, _32618_);
  nor (_32620_, _32266_, _32029_);
  and (_32621_, _32620_, _32601_);
  and (_32622_, _32612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_33693_, _32622_, _32621_);
  nor (_32623_, _32484_, _32029_);
  and (_32624_, _32623_, _32601_);
  and (_32625_, _32612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_33698_, _32625_, _32624_);
  and (_32626_, _32601_, _32594_);
  and (_32627_, _32612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_33701_, _32627_, _32626_);
  and (_32628_, _32588_, _32081_);
  and (_32629_, _32628_, _32599_);
  and (_32630_, _32629_, _32602_);
  not (_32631_, _32629_);
  and (_32632_, _32631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_33707_, _32632_, _32630_);
  and (_32633_, _32629_, _32606_);
  and (_32634_, _32631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_33711_, _32634_, _32633_);
  and (_32635_, _32629_, _32610_);
  and (_32636_, _32631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_33714_, _32636_, _32635_);
  and (_32637_, _32629_, _32614_);
  and (_32638_, _32631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_33718_, _32638_, _32637_);
  and (_32639_, _32629_, _32617_);
  not (_32640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_32641_, _32629_, _32640_);
  or (_33721_, _32641_, _32639_);
  and (_32642_, _32629_, _32620_);
  not (_32643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_32644_, _32629_, _32643_);
  or (_33725_, _32644_, _32642_);
  and (_32645_, _32629_, _32623_);
  not (_32646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_32647_, _32629_, _32646_);
  or (_33728_, _32647_, _32645_);
  and (_32648_, _32629_, _32594_);
  and (_32649_, _32631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_33731_, _32649_, _32648_);
  and (_32650_, _32587_, _32033_);
  and (_32651_, _32650_, _32599_);
  and (_32652_, _32651_, _32602_);
  not (_32653_, _32651_);
  and (_32654_, _32653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_33738_, _32654_, _32652_);
  and (_32655_, _32651_, _32606_);
  and (_32656_, _32653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_33741_, _32656_, _32655_);
  and (_32657_, _32651_, _32610_);
  not (_32658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_32659_, _32651_, _32658_);
  or (_33745_, _32659_, _32657_);
  and (_32660_, _32651_, _32614_);
  and (_32661_, _32653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_33748_, _32661_, _32660_);
  and (_32662_, _32651_, _32617_);
  not (_32663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_32664_, _32651_, _32663_);
  or (_33752_, _32664_, _32662_);
  and (_32665_, _32651_, _32620_);
  not (_32666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_32667_, _32651_, _32666_);
  or (_33756_, _32667_, _32665_);
  and (_32668_, _32651_, _32623_);
  not (_32669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_32670_, _32651_, _32669_);
  or (_33759_, _32670_, _32668_);
  and (_32671_, _32651_, _32594_);
  not (_32672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_32673_, _32651_, _32672_);
  or (_33762_, _32673_, _32671_);
  and (_32674_, _32599_, _32589_);
  and (_32675_, _32674_, _32602_);
  not (_32676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_32677_, _32674_, _32676_);
  or (_33767_, _32677_, _32675_);
  and (_32678_, _32674_, _32606_);
  not (_32679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_32680_, _32674_, _32679_);
  or (_33770_, _32680_, _32678_);
  and (_32681_, _32674_, _32610_);
  not (_32682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_32683_, _32674_, _32682_);
  or (_33774_, _32683_, _32681_);
  and (_32684_, _32674_, _32614_);
  not (_32685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_32686_, _32674_, _32685_);
  or (_33777_, _32686_, _32684_);
  and (_32687_, _32674_, _32617_);
  not (_32688_, _32674_);
  and (_32689_, _32688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_33781_, _32689_, _32687_);
  and (_32690_, _32674_, _32620_);
  and (_32691_, _32688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_33784_, _32691_, _32690_);
  and (_32692_, _32674_, _32623_);
  and (_32693_, _32688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_33788_, _32693_, _32692_);
  and (_32694_, _32674_, _32594_);
  nor (_32695_, _32674_, _32537_);
  or (_33791_, _32695_, _32694_);
  and (_32696_, _32590_, _32472_);
  and (_32697_, _32696_, _32598_);
  and (_32698_, _32697_, _32602_);
  not (_32699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_32700_, _32697_, _32699_);
  or (_33797_, _32700_, _32698_);
  and (_32701_, _32697_, _32606_);
  not (_32702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_32703_, _32697_, _32702_);
  or (_36087_, _32703_, _32701_);
  and (_32704_, _32697_, _32610_);
  not (_32705_, _32697_);
  and (_32706_, _32705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_36088_, _32706_, _32704_);
  and (_32707_, _32697_, _32614_);
  and (_32708_, _32705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_36089_, _32708_, _32707_);
  and (_32709_, _32697_, _32617_);
  and (_32710_, _32705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_36090_, _32710_, _32709_);
  and (_32711_, _32697_, _32620_);
  and (_32712_, _32705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_36091_, _32712_, _32711_);
  and (_32713_, _32697_, _32623_);
  not (_32714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_32715_, _32697_, _32714_);
  or (_36092_, _32715_, _32713_);
  and (_32716_, _32697_, _32594_);
  and (_32717_, _32705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_36093_, _32717_, _32716_);
  and (_32718_, _32696_, _32628_);
  and (_32719_, _32718_, _32602_);
  not (_32720_, _32718_);
  and (_32721_, _32720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_36094_, _32721_, _32719_);
  and (_32722_, _32718_, _32606_);
  and (_32723_, _32720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_36095_, _32723_, _32722_);
  and (_32724_, _32718_, _32610_);
  and (_32725_, _32720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_36096_, _32725_, _32724_);
  and (_32726_, _32718_, _32614_);
  and (_32727_, _32720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_36097_, _32727_, _32726_);
  and (_32728_, _32718_, _32617_);
  not (_32729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_32730_, _32718_, _32729_);
  or (_36098_, _32730_, _32728_);
  and (_32731_, _32718_, _32620_);
  not (_32732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_32733_, _32718_, _32732_);
  or (_36099_, _32733_, _32731_);
  and (_32734_, _32718_, _32623_);
  and (_32735_, _32720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_36100_, _32735_, _32734_);
  and (_32736_, _32718_, _32594_);
  and (_32737_, _32720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_36101_, _32737_, _32736_);
  and (_32738_, _32696_, _32650_);
  and (_32739_, _32738_, _32602_);
  not (_32740_, _32738_);
  and (_32741_, _32740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_36102_, _32741_, _32739_);
  and (_32742_, _32738_, _32606_);
  and (_32743_, _32740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_36103_, _32743_, _32742_);
  and (_32744_, _32738_, _32610_);
  not (_32745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_32746_, _32738_, _32745_);
  or (_36104_, _32746_, _32744_);
  and (_32747_, _32738_, _32614_);
  and (_32748_, _32740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_36105_, _32748_, _32747_);
  and (_32749_, _32738_, _32617_);
  not (_32750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_32751_, _32738_, _32750_);
  or (_36106_, _32751_, _32749_);
  and (_32752_, _32738_, _32620_);
  not (_32753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_32754_, _32738_, _32753_);
  or (_36107_, _32754_, _32752_);
  and (_32755_, _32738_, _32623_);
  and (_32756_, _32740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_36108_, _32756_, _32755_);
  and (_32757_, _32738_, _32594_);
  not (_32758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_32759_, _32738_, _32758_);
  or (_36109_, _32759_, _32757_);
  and (_32760_, _32696_, _32589_);
  and (_32761_, _32760_, _32602_);
  not (_32762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_32763_, _32760_, _32762_);
  or (_36110_, _32763_, _32761_);
  and (_32764_, _32760_, _32606_);
  not (_32765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_32766_, _32760_, _32765_);
  or (_36111_, _32766_, _32764_);
  and (_32767_, _32760_, _32610_);
  not (_32768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_32769_, _32760_, _32768_);
  or (_36112_, _32769_, _32767_);
  and (_32770_, _32760_, _32614_);
  not (_32771_, _32760_);
  and (_32772_, _32771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_36113_, _32772_, _32770_);
  and (_32773_, _32760_, _32617_);
  and (_32774_, _32771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_36114_, _32774_, _32773_);
  and (_32775_, _32760_, _32620_);
  and (_32776_, _32771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_36115_, _32776_, _32775_);
  and (_32777_, _32760_, _32623_);
  not (_32778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_32779_, _32760_, _32778_);
  or (_36116_, _32779_, _32777_);
  and (_32780_, _32760_, _32594_);
  nor (_32781_, _32760_, _32549_);
  or (_36117_, _32781_, _32780_);
  and (_32782_, _32591_, _32077_);
  and (_32783_, _32782_, _32598_);
  and (_32784_, _32783_, _32602_);
  not (_32785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_32786_, _32783_, _32785_);
  or (_36118_, _32786_, _32784_);
  and (_32787_, _32783_, _32606_);
  not (_32788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_32789_, _32783_, _32788_);
  or (_36119_, _32789_, _32787_);
  and (_32790_, _32783_, _32610_);
  not (_32791_, _32783_);
  and (_32792_, _32791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_36120_, _32792_, _32790_);
  and (_32793_, _32783_, _32614_);
  and (_32794_, _32791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_36121_, _32794_, _32793_);
  and (_32795_, _32783_, _32617_);
  and (_32796_, _32791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_36122_, _32796_, _32795_);
  and (_32797_, _32783_, _32620_);
  and (_32798_, _32791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_36123_, _32798_, _32797_);
  and (_32799_, _32783_, _32623_);
  not (_32800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_32801_, _32783_, _32800_);
  or (_36124_, _32801_, _32799_);
  and (_32802_, _32783_, _32594_);
  and (_32803_, _32791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_36125_, _32803_, _32802_);
  and (_32804_, _32782_, _32628_);
  and (_32805_, _32804_, _32602_);
  not (_32806_, _32804_);
  and (_32807_, _32806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_36126_, _32807_, _32805_);
  and (_32808_, _32804_, _32606_);
  and (_32809_, _32806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_36127_, _32809_, _32808_);
  and (_32810_, _32804_, _32610_);
  and (_32811_, _32806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_36128_, _32811_, _32810_);
  and (_32812_, _32804_, _32614_);
  not (_32813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_32814_, _32804_, _32813_);
  or (_36129_, _32814_, _32812_);
  and (_32815_, _32804_, _32617_);
  not (_32816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_32817_, _32804_, _32816_);
  or (_36130_, _32817_, _32815_);
  and (_32818_, _32804_, _32620_);
  not (_32819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_32820_, _32804_, _32819_);
  or (_36131_, _32820_, _32818_);
  and (_32821_, _32804_, _32623_);
  and (_32822_, _32806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_36132_, _32822_, _32821_);
  and (_32823_, _32804_, _32594_);
  and (_32824_, _32806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_36133_, _32824_, _32823_);
  and (_32825_, _32782_, _32650_);
  and (_32826_, _32825_, _32602_);
  not (_32827_, _32825_);
  and (_32828_, _32827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_36040_, _32828_, _32826_);
  and (_32829_, _32825_, _32606_);
  and (_32830_, _32827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_36041_, _32830_, _32829_);
  and (_32831_, _32825_, _32610_);
  not (_32832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_32833_, _32825_, _32832_);
  or (_36042_, _32833_, _32831_);
  and (_32834_, _32825_, _32614_);
  not (_32835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_32836_, _32825_, _32835_);
  or (_36043_, _32836_, _32834_);
  and (_32837_, _32825_, _32617_);
  not (_32838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_32839_, _32825_, _32838_);
  or (_36044_, _32839_, _32837_);
  and (_32840_, _32825_, _32620_);
  not (_32841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_32842_, _32825_, _32841_);
  or (_36045_, _32842_, _32840_);
  and (_32843_, _32825_, _32623_);
  not (_32844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_32845_, _32825_, _32844_);
  or (_36046_, _32845_, _32843_);
  and (_32846_, _32825_, _32594_);
  nor (_32847_, _32825_, _32563_);
  or (_36047_, _32847_, _32846_);
  and (_32848_, _32782_, _32589_);
  and (_32849_, _32848_, _32602_);
  not (_32850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_32851_, _32848_, _32850_);
  or (_36048_, _32851_, _32849_);
  and (_32852_, _32848_, _32606_);
  not (_32853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_32854_, _32848_, _32853_);
  or (_36049_, _32854_, _32852_);
  and (_32855_, _32848_, _32610_);
  not (_32856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_32857_, _32848_, _32856_);
  or (_36050_, _32857_, _32855_);
  and (_32858_, _32848_, _32614_);
  not (_32859_, _32848_);
  and (_32860_, _32859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_36051_, _32860_, _32858_);
  and (_32861_, _32848_, _32617_);
  and (_32862_, _32859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_36052_, _32862_, _32861_);
  and (_32863_, _32848_, _32620_);
  and (_32864_, _32859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_36053_, _32864_, _32863_);
  and (_32865_, _32848_, _32623_);
  and (_32866_, _32859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_36054_, _32866_, _32865_);
  and (_32867_, _32848_, _32594_);
  not (_32868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_32869_, _32848_, _32868_);
  or (_36055_, _32869_, _32867_);
  and (_32870_, _32598_, _32592_);
  and (_32871_, _32870_, _32602_);
  not (_32872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_32873_, _32870_, _32872_);
  or (_36056_, _32873_, _32871_);
  and (_32874_, _32870_, _32606_);
  not (_32875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_32876_, _32870_, _32875_);
  or (_36057_, _32876_, _32874_);
  and (_32877_, _32870_, _32610_);
  not (_32878_, _32870_);
  and (_32879_, _32878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_36058_, _32879_, _32877_);
  and (_32880_, _32870_, _32614_);
  and (_32881_, _32878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_36059_, _32881_, _32880_);
  and (_32882_, _32870_, _32617_);
  and (_32883_, _32878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_36060_, _32883_, _32882_);
  and (_32884_, _32870_, _32620_);
  and (_32885_, _32878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_36061_, _32885_, _32884_);
  and (_32886_, _32870_, _32623_);
  and (_32887_, _32878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_36062_, _32887_, _32886_);
  and (_32888_, _32870_, _32594_);
  and (_32889_, _32878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_36063_, _32889_, _32888_);
  and (_32890_, _32628_, _32592_);
  and (_32891_, _32890_, _32602_);
  not (_32892_, _32890_);
  and (_32893_, _32892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_36064_, _32893_, _32891_);
  and (_32894_, _32890_, _32606_);
  and (_32895_, _32892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_36065_, _32895_, _32894_);
  and (_32896_, _32890_, _32610_);
  and (_32897_, _32892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_36066_, _32897_, _32896_);
  and (_32898_, _32890_, _32614_);
  not (_32899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_32900_, _32890_, _32899_);
  or (_36067_, _32900_, _32898_);
  and (_32901_, _32890_, _32617_);
  not (_32902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_32903_, _32890_, _32902_);
  or (_36068_, _32903_, _32901_);
  and (_32904_, _32890_, _32620_);
  not (_32905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_32906_, _32890_, _32905_);
  or (_36069_, _32906_, _32904_);
  and (_32907_, _32890_, _32623_);
  not (_32908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_32909_, _32890_, _32908_);
  or (_36070_, _32909_, _32907_);
  and (_32910_, _32890_, _32594_);
  and (_32911_, _32892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_36071_, _32911_, _32910_);
  and (_32912_, _32650_, _32592_);
  and (_32913_, _32912_, _32602_);
  not (_32914_, _32912_);
  and (_32915_, _32914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_36072_, _32915_, _32913_);
  and (_32916_, _32912_, _32606_);
  and (_32917_, _32914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_36073_, _32917_, _32916_);
  and (_32918_, _32912_, _32610_);
  not (_32919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_32920_, _32912_, _32919_);
  or (_36074_, _32920_, _32918_);
  and (_32921_, _32912_, _32614_);
  not (_32922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_32923_, _32912_, _32922_);
  or (_36075_, _32923_, _32921_);
  and (_32924_, _32912_, _32617_);
  not (_32925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_32926_, _32912_, _32925_);
  or (_36076_, _32926_, _32924_);
  and (_32927_, _32912_, _32620_);
  not (_32928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_32929_, _32912_, _32928_);
  or (_36077_, _32929_, _32927_);
  and (_32930_, _32912_, _32623_);
  not (_32931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_32932_, _32912_, _32931_);
  or (_36078_, _32932_, _32930_);
  and (_32933_, _32912_, _32594_);
  nor (_32934_, _32912_, _32574_);
  or (_36079_, _32934_, _32933_);
  and (_32935_, _32602_, _32593_);
  not (_32936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_32937_, _32593_, _32936_);
  or (_36080_, _32937_, _32935_);
  and (_32938_, _32606_, _32593_);
  not (_32939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_32940_, _32593_, _32939_);
  or (_36081_, _32940_, _32938_);
  and (_32941_, _32610_, _32593_);
  not (_32942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_32943_, _32593_, _32942_);
  or (_36082_, _32943_, _32941_);
  and (_32944_, _32614_, _32593_);
  not (_32945_, _32593_);
  and (_32946_, _32945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_36083_, _32946_, _32944_);
  and (_32947_, _32617_, _32593_);
  and (_32948_, _32945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_36084_, _32948_, _32947_);
  and (_32949_, _32620_, _32593_);
  and (_32950_, _32945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_36085_, _32950_, _32949_);
  and (_32951_, _32623_, _32593_);
  and (_32952_, _32945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_36086_, _32952_, _32951_);
  or (_32953_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_32954_, _32252_, _32604_);
  and (_32955_, _32954_, _32465_);
  and (_32956_, _32955_, _32953_);
  nor (_32957_, _32252_, _32676_);
  and (_32958_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_32959_, _32958_, _32957_);
  and (_32960_, _32959_, _32536_);
  or (_32961_, _32960_, _32956_);
  or (_32962_, _32961_, _32530_);
  or (_32963_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_32964_, _32252_, _32699_);
  and (_32965_, _32964_, _32465_);
  and (_32966_, _32965_, _32963_);
  nor (_32967_, _32252_, _32762_);
  and (_32968_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_32969_, _32968_, _32967_);
  and (_32970_, _32969_, _32536_);
  or (_32971_, _32970_, _32966_);
  or (_32972_, _32971_, _32356_);
  and (_32973_, _32972_, _32544_);
  and (_32974_, _32973_, _32962_);
  nand (_32975_, _32252_, _32785_);
  or (_32976_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_32977_, _32976_, _32975_);
  and (_32978_, _32977_, _32465_);
  and (_32979_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_32980_, _32252_, _32850_);
  or (_32981_, _32980_, _32979_);
  and (_32982_, _32981_, _32536_);
  or (_32983_, _32982_, _32978_);
  or (_32984_, _32983_, _32530_);
  nand (_32985_, _32252_, _32872_);
  or (_32986_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_32987_, _32986_, _32985_);
  and (_32988_, _32987_, _32465_);
  and (_32989_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_32990_, _32252_, _32936_);
  or (_32991_, _32990_, _32989_);
  and (_32992_, _32991_, _32536_);
  or (_32993_, _32992_, _32988_);
  or (_32994_, _32993_, _32356_);
  and (_32995_, _32994_, _32523_);
  and (_32996_, _32995_, _32984_);
  or (_32997_, _32996_, _32974_);
  or (_32998_, _32997_, _32529_);
  or (_32999_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_33000_, _32999_, _35796_);
  and (_36134_[0], _33000_, _32998_);
  or (_33001_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_33002_, _32252_, _32608_);
  and (_33003_, _33002_, _32465_);
  and (_33004_, _33003_, _33001_);
  nor (_33005_, _32252_, _32679_);
  and (_33006_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_33007_, _33006_, _33005_);
  and (_33008_, _33007_, _32536_);
  or (_33009_, _33008_, _33004_);
  or (_33010_, _33009_, _32530_);
  or (_33011_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_33012_, _32252_, _32702_);
  and (_33013_, _33012_, _32465_);
  and (_33014_, _33013_, _33011_);
  nor (_33015_, _32252_, _32765_);
  and (_33016_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_33017_, _33016_, _33015_);
  and (_33018_, _33017_, _32536_);
  or (_33019_, _33018_, _33014_);
  or (_33020_, _33019_, _32356_);
  and (_33021_, _33020_, _32544_);
  and (_33022_, _33021_, _33010_);
  nand (_33023_, _32252_, _32788_);
  or (_33024_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_33025_, _33024_, _33023_);
  and (_33026_, _33025_, _32465_);
  and (_33027_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_33028_, _32252_, _32853_);
  or (_33029_, _33028_, _33027_);
  and (_33030_, _33029_, _32536_);
  or (_33031_, _33030_, _33026_);
  or (_33032_, _33031_, _32530_);
  nand (_33033_, _32252_, _32875_);
  or (_33034_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_33035_, _33034_, _33033_);
  and (_33036_, _33035_, _32465_);
  and (_33037_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_33038_, _32252_, _32939_);
  or (_33039_, _33038_, _33037_);
  and (_33040_, _33039_, _32536_);
  or (_33041_, _33040_, _33036_);
  or (_33042_, _33041_, _32356_);
  and (_33043_, _33042_, _32523_);
  and (_33044_, _33043_, _33032_);
  or (_33045_, _33044_, _33022_);
  or (_33046_, _33045_, _32529_);
  or (_33047_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_33048_, _33047_, _35796_);
  and (_36134_[1], _33048_, _33046_);
  and (_33049_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_33050_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_33051_, _33050_, _33049_);
  and (_33052_, _33051_, _32465_);
  nor (_33053_, _32252_, _32682_);
  and (_33054_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_33055_, _33054_, _33053_);
  and (_33056_, _33055_, _32536_);
  or (_33057_, _33056_, _33052_);
  or (_33058_, _33057_, _32530_);
  and (_33059_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_33060_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_33061_, _33060_, _33059_);
  and (_33062_, _33061_, _32465_);
  nor (_33063_, _32252_, _32768_);
  and (_33064_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_33065_, _33064_, _33063_);
  and (_33066_, _33065_, _32536_);
  or (_33067_, _33066_, _33062_);
  or (_33068_, _33067_, _32356_);
  and (_33069_, _33068_, _32544_);
  and (_33070_, _33069_, _33058_);
  or (_33071_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_33072_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_33073_, _33072_, _33071_);
  and (_33074_, _33073_, _32465_);
  or (_33075_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_33076_, _32252_, _32832_);
  and (_33077_, _33076_, _33075_);
  and (_33078_, _33077_, _32536_);
  or (_33079_, _33078_, _33074_);
  or (_33080_, _33079_, _32530_);
  or (_33081_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_33082_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_33083_, _33082_, _33081_);
  and (_33084_, _33083_, _32465_);
  or (_33085_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_33086_, _32252_, _32919_);
  and (_33087_, _33086_, _33085_);
  and (_33088_, _33087_, _32536_);
  or (_33089_, _33088_, _33084_);
  or (_33090_, _33089_, _32356_);
  and (_33091_, _33090_, _32523_);
  and (_33092_, _33091_, _33080_);
  or (_33093_, _33092_, _33070_);
  or (_33094_, _33093_, _32529_);
  or (_33095_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_33096_, _33095_, _35796_);
  and (_36134_[2], _33096_, _33094_);
  or (_33097_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_33098_, _32252_, _32922_);
  and (_33099_, _33098_, _33097_);
  or (_33100_, _33099_, _32465_);
  and (_33101_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_33102_, _32252_, _32899_);
  or (_33103_, _33102_, _33101_);
  or (_33104_, _33103_, _32536_);
  and (_33105_, _33104_, _32523_);
  and (_33106_, _33105_, _33100_);
  and (_33107_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_33108_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_33109_, _33108_, _32536_);
  or (_33110_, _33109_, _33107_);
  and (_33111_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_33112_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_33113_, _33112_, _32465_);
  or (_33114_, _33113_, _33111_);
  and (_33115_, _33114_, _32544_);
  and (_33116_, _33115_, _33110_);
  or (_33117_, _33116_, _33106_);
  and (_33118_, _33117_, _32530_);
  or (_33119_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_33120_, _32252_, _32835_);
  and (_33121_, _33120_, _33119_);
  or (_33122_, _33121_, _32465_);
  and (_33123_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_33124_, _32252_, _32813_);
  or (_33125_, _33124_, _33123_);
  or (_33126_, _33125_, _32536_);
  and (_33127_, _33126_, _32523_);
  and (_33128_, _33127_, _33122_);
  and (_33129_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_33130_, _32532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_33131_, _33130_, _32536_);
  or (_33132_, _33131_, _33129_);
  nor (_33133_, _32252_, _32685_);
  and (_33134_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_33135_, _33134_, _32465_);
  or (_33136_, _33135_, _33133_);
  and (_33137_, _33136_, _32544_);
  and (_33138_, _33137_, _33132_);
  or (_33139_, _33138_, _33128_);
  and (_33140_, _33139_, _32356_);
  or (_33141_, _33140_, _32529_);
  or (_33142_, _33141_, _33118_);
  or (_33143_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_33144_, _33143_, _35796_);
  and (_36134_[3], _33144_, _33142_);
  and (_33145_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_33146_, _32252_, _32640_);
  or (_33147_, _33146_, _33145_);
  and (_33148_, _33147_, _32465_);
  or (_33149_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_33150_, _32252_, _32663_);
  and (_33151_, _33150_, _33149_);
  and (_33152_, _33151_, _32536_);
  or (_33153_, _33152_, _33148_);
  or (_33154_, _33153_, _32530_);
  and (_33155_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_33156_, _32252_, _32729_);
  or (_33157_, _33156_, _33155_);
  and (_33158_, _33157_, _32465_);
  or (_33159_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_33160_, _32252_, _32750_);
  and (_33161_, _33160_, _33159_);
  and (_33162_, _33161_, _32536_);
  or (_33163_, _33162_, _33158_);
  or (_33164_, _33163_, _32356_);
  and (_33165_, _33164_, _32544_);
  and (_33166_, _33165_, _33154_);
  and (_33167_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_33168_, _32252_, _32816_);
  or (_33169_, _33168_, _33167_);
  and (_33170_, _33169_, _32465_);
  or (_33171_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_33172_, _32252_, _32838_);
  and (_33173_, _33172_, _33171_);
  and (_33174_, _33173_, _32536_);
  or (_33175_, _33174_, _33170_);
  or (_33176_, _33175_, _32530_);
  and (_33177_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_33178_, _32252_, _32902_);
  or (_33179_, _33178_, _33177_);
  and (_33180_, _33179_, _32465_);
  or (_33181_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_33182_, _32252_, _32925_);
  and (_33183_, _33182_, _33181_);
  and (_33184_, _33183_, _32536_);
  or (_33185_, _33184_, _33180_);
  or (_33186_, _33185_, _32356_);
  and (_33187_, _33186_, _32523_);
  and (_33188_, _33187_, _33176_);
  or (_33189_, _33188_, _33166_);
  or (_33190_, _33189_, _32529_);
  or (_33191_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_33192_, _33191_, _35796_);
  and (_36134_[4], _33192_, _33190_);
  and (_33193_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_33194_, _32252_, _32643_);
  or (_33195_, _33194_, _33193_);
  and (_33196_, _33195_, _32465_);
  or (_33197_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_33198_, _32252_, _32666_);
  and (_33199_, _33198_, _33197_);
  and (_33200_, _33199_, _32536_);
  or (_33201_, _33200_, _33196_);
  or (_33202_, _33201_, _32530_);
  and (_33203_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_33204_, _32252_, _32732_);
  or (_33205_, _33204_, _33203_);
  and (_33206_, _33205_, _32465_);
  or (_33207_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_33208_, _32252_, _32753_);
  and (_33209_, _33208_, _33207_);
  and (_33210_, _33209_, _32536_);
  or (_33211_, _33210_, _33206_);
  or (_33212_, _33211_, _32356_);
  and (_33213_, _33212_, _32544_);
  and (_33214_, _33213_, _33202_);
  and (_33215_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_33216_, _32252_, _32819_);
  or (_33217_, _33216_, _33215_);
  and (_33218_, _33217_, _32465_);
  or (_33219_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_33220_, _32252_, _32841_);
  and (_33221_, _33220_, _33219_);
  and (_33222_, _33221_, _32536_);
  or (_33223_, _33222_, _33218_);
  or (_33224_, _33223_, _32530_);
  and (_33225_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_33226_, _32252_, _32905_);
  or (_33227_, _33226_, _33225_);
  and (_33228_, _33227_, _32465_);
  or (_33229_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_33230_, _32252_, _32928_);
  and (_33231_, _33230_, _33229_);
  and (_33232_, _33231_, _32536_);
  or (_33233_, _33232_, _33228_);
  or (_33234_, _33233_, _32356_);
  and (_33235_, _33234_, _32523_);
  and (_33236_, _33235_, _33224_);
  or (_33237_, _33236_, _33214_);
  or (_33238_, _33237_, _32529_);
  or (_33239_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_33240_, _33239_, _35796_);
  and (_36134_[5], _33240_, _33238_);
  and (_33241_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_33242_, _32252_, _32646_);
  or (_33243_, _33242_, _33241_);
  and (_33244_, _33243_, _32465_);
  or (_33245_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand (_33246_, _32252_, _32669_);
  and (_33247_, _33246_, _33245_);
  and (_33248_, _33247_, _32536_);
  or (_33249_, _33248_, _33244_);
  or (_33250_, _33249_, _32530_);
  or (_33251_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nand (_33252_, _32252_, _32714_);
  and (_33253_, _33252_, _32465_);
  and (_33254_, _33253_, _33251_);
  nor (_33255_, _32252_, _32778_);
  and (_33256_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_33257_, _33256_, _33255_);
  and (_33258_, _33257_, _32536_);
  or (_33259_, _33258_, _33254_);
  or (_33260_, _33259_, _32356_);
  and (_33261_, _33260_, _32544_);
  and (_33262_, _33261_, _33250_);
  nand (_33263_, _32252_, _32800_);
  or (_33264_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_33265_, _33264_, _33263_);
  and (_33266_, _33265_, _32465_);
  or (_33267_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_33268_, _32252_, _32844_);
  and (_33269_, _33268_, _33267_);
  and (_33270_, _33269_, _32536_);
  or (_33271_, _33270_, _33266_);
  or (_33272_, _33271_, _32530_);
  and (_33273_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_33274_, _32252_, _32908_);
  or (_33275_, _33274_, _33273_);
  and (_33276_, _33275_, _32465_);
  or (_33277_, _32252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_33278_, _32252_, _32931_);
  and (_33279_, _33278_, _33277_);
  and (_33280_, _33279_, _32536_);
  or (_33281_, _33280_, _33276_);
  or (_33282_, _33281_, _32356_);
  and (_33283_, _33282_, _32523_);
  and (_33284_, _33283_, _33272_);
  or (_33285_, _33284_, _33262_);
  or (_33286_, _33285_, _32529_);
  or (_33287_, _32584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_33288_, _33287_, _35796_);
  and (_36134_[6], _33288_, _33286_);
  or (_33291_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_33293_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_33295_, _33293_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_33297_, _33295_, _33291_);
  nand (_33299_, _33297_, _35796_);
  or (_33301_, \oc8051_gm_cxrom_1.cell0.data [7], _35796_);
  and (_35795_[7], _33301_, _33299_);
  or (_33304_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33306_, \oc8051_gm_cxrom_1.cell0.data [0], _33293_);
  nand (_33308_, _33306_, _33304_);
  nand (_33310_, _33308_, _35796_);
  or (_33312_, \oc8051_gm_cxrom_1.cell0.data [0], _35796_);
  and (_35795_[0], _33312_, _33310_);
  or (_33315_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33317_, \oc8051_gm_cxrom_1.cell0.data [1], _33293_);
  nand (_33319_, _33317_, _33315_);
  nand (_33321_, _33319_, _35796_);
  or (_33323_, \oc8051_gm_cxrom_1.cell0.data [1], _35796_);
  and (_35795_[1], _33323_, _33321_);
  or (_33326_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33328_, \oc8051_gm_cxrom_1.cell0.data [2], _33293_);
  nand (_33330_, _33328_, _33326_);
  nand (_33332_, _33330_, _35796_);
  or (_33334_, \oc8051_gm_cxrom_1.cell0.data [2], _35796_);
  and (_35795_[2], _33334_, _33332_);
  or (_33337_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33339_, \oc8051_gm_cxrom_1.cell0.data [3], _33293_);
  nand (_33340_, _33339_, _33337_);
  nand (_33341_, _33340_, _35796_);
  or (_33342_, \oc8051_gm_cxrom_1.cell0.data [3], _35796_);
  and (_35795_[3], _33342_, _33341_);
  or (_33343_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33344_, \oc8051_gm_cxrom_1.cell0.data [4], _33293_);
  nand (_33345_, _33344_, _33343_);
  nand (_33346_, _33345_, _35796_);
  or (_33347_, \oc8051_gm_cxrom_1.cell0.data [4], _35796_);
  and (_35795_[4], _33347_, _33346_);
  or (_33348_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33349_, \oc8051_gm_cxrom_1.cell0.data [5], _33293_);
  nand (_33350_, _33349_, _33348_);
  nand (_33351_, _33350_, _35796_);
  or (_33352_, \oc8051_gm_cxrom_1.cell0.data [5], _35796_);
  and (_35795_[5], _33352_, _33351_);
  or (_33353_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33354_, \oc8051_gm_cxrom_1.cell0.data [6], _33293_);
  nand (_33355_, _33354_, _33353_);
  nand (_33356_, _33355_, _35796_);
  or (_33357_, \oc8051_gm_cxrom_1.cell0.data [6], _35796_);
  and (_35795_[6], _33357_, _33356_);
  or (_33358_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_33359_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_33360_, _33359_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_33361_, _33360_, _33358_);
  nand (_33362_, _33361_, _35796_);
  or (_33363_, \oc8051_gm_cxrom_1.cell1.data [7], _35796_);
  and (_35797_[7], _33363_, _33362_);
  or (_33364_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33365_, \oc8051_gm_cxrom_1.cell1.data [0], _33359_);
  nand (_33366_, _33365_, _33364_);
  nand (_33367_, _33366_, _35796_);
  or (_33368_, \oc8051_gm_cxrom_1.cell1.data [0], _35796_);
  and (_35797_[0], _33368_, _33367_);
  or (_33369_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33370_, \oc8051_gm_cxrom_1.cell1.data [1], _33359_);
  nand (_33371_, _33370_, _33369_);
  nand (_33372_, _33371_, _35796_);
  or (_33373_, \oc8051_gm_cxrom_1.cell1.data [1], _35796_);
  and (_35797_[1], _33373_, _33372_);
  or (_33374_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33375_, \oc8051_gm_cxrom_1.cell1.data [2], _33359_);
  nand (_33376_, _33375_, _33374_);
  nand (_33377_, _33376_, _35796_);
  or (_33378_, \oc8051_gm_cxrom_1.cell1.data [2], _35796_);
  and (_35797_[2], _33378_, _33377_);
  or (_33379_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33380_, \oc8051_gm_cxrom_1.cell1.data [3], _33359_);
  nand (_33381_, _33380_, _33379_);
  nand (_33382_, _33381_, _35796_);
  or (_33383_, \oc8051_gm_cxrom_1.cell1.data [3], _35796_);
  and (_35797_[3], _33383_, _33382_);
  or (_33384_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33385_, \oc8051_gm_cxrom_1.cell1.data [4], _33359_);
  nand (_33386_, _33385_, _33384_);
  nand (_33387_, _33386_, _35796_);
  or (_33388_, \oc8051_gm_cxrom_1.cell1.data [4], _35796_);
  and (_35797_[4], _33388_, _33387_);
  or (_33389_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33390_, \oc8051_gm_cxrom_1.cell1.data [5], _33359_);
  nand (_33391_, _33390_, _33389_);
  nand (_33392_, _33391_, _35796_);
  or (_33393_, \oc8051_gm_cxrom_1.cell1.data [5], _35796_);
  and (_35797_[5], _33393_, _33392_);
  or (_33394_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33395_, \oc8051_gm_cxrom_1.cell1.data [6], _33359_);
  nand (_33396_, _33395_, _33394_);
  nand (_33397_, _33396_, _35796_);
  or (_33398_, \oc8051_gm_cxrom_1.cell1.data [6], _35796_);
  and (_35797_[6], _33398_, _33397_);
  or (_33399_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_33400_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_33401_, _33400_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_33402_, _33401_, _33399_);
  nand (_33403_, _33402_, _35796_);
  or (_33404_, \oc8051_gm_cxrom_1.cell2.data [7], _35796_);
  and (_35811_[7], _33404_, _33403_);
  or (_33405_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33406_, \oc8051_gm_cxrom_1.cell2.data [0], _33400_);
  nand (_33407_, _33406_, _33405_);
  nand (_33408_, _33407_, _35796_);
  or (_33409_, \oc8051_gm_cxrom_1.cell2.data [0], _35796_);
  and (_35811_[0], _33409_, _33408_);
  or (_33410_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33411_, \oc8051_gm_cxrom_1.cell2.data [1], _33400_);
  nand (_33412_, _33411_, _33410_);
  nand (_33413_, _33412_, _35796_);
  or (_33415_, \oc8051_gm_cxrom_1.cell2.data [1], _35796_);
  and (_35811_[1], _33415_, _33413_);
  or (_33416_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33417_, \oc8051_gm_cxrom_1.cell2.data [2], _33400_);
  nand (_33418_, _33417_, _33416_);
  nand (_33419_, _33418_, _35796_);
  or (_33420_, \oc8051_gm_cxrom_1.cell2.data [2], _35796_);
  and (_35811_[2], _33420_, _33419_);
  or (_33421_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33422_, \oc8051_gm_cxrom_1.cell2.data [3], _33400_);
  nand (_33423_, _33422_, _33421_);
  nand (_33425_, _33423_, _35796_);
  or (_33426_, \oc8051_gm_cxrom_1.cell2.data [3], _35796_);
  and (_35811_[3], _33426_, _33425_);
  or (_33427_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33428_, \oc8051_gm_cxrom_1.cell2.data [4], _33400_);
  nand (_33429_, _33428_, _33427_);
  nand (_33430_, _33429_, _35796_);
  or (_33431_, \oc8051_gm_cxrom_1.cell2.data [4], _35796_);
  and (_35811_[4], _33431_, _33430_);
  or (_33432_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33433_, \oc8051_gm_cxrom_1.cell2.data [5], _33400_);
  nand (_33434_, _33433_, _33432_);
  nand (_33435_, _33434_, _35796_);
  or (_33436_, \oc8051_gm_cxrom_1.cell2.data [5], _35796_);
  and (_35811_[5], _33436_, _33435_);
  or (_33437_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33438_, \oc8051_gm_cxrom_1.cell2.data [6], _33400_);
  nand (_33439_, _33438_, _33437_);
  nand (_33440_, _33439_, _35796_);
  or (_33441_, \oc8051_gm_cxrom_1.cell2.data [6], _35796_);
  and (_35811_[6], _33441_, _33440_);
  or (_33442_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_33443_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_33444_, _33443_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_33445_, _33444_, _33442_);
  nand (_33446_, _33445_, _35796_);
  or (_33447_, \oc8051_gm_cxrom_1.cell3.data [7], _35796_);
  and (_35813_[7], _33447_, _33446_);
  or (_33448_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33449_, \oc8051_gm_cxrom_1.cell3.data [0], _33443_);
  nand (_33450_, _33449_, _33448_);
  nand (_33451_, _33450_, _35796_);
  or (_33452_, \oc8051_gm_cxrom_1.cell3.data [0], _35796_);
  and (_35813_[0], _33452_, _33451_);
  or (_33453_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33454_, \oc8051_gm_cxrom_1.cell3.data [1], _33443_);
  nand (_33455_, _33454_, _33453_);
  nand (_33456_, _33455_, _35796_);
  or (_33457_, \oc8051_gm_cxrom_1.cell3.data [1], _35796_);
  and (_35813_[1], _33457_, _33456_);
  or (_33458_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33459_, \oc8051_gm_cxrom_1.cell3.data [2], _33443_);
  nand (_33460_, _33459_, _33458_);
  nand (_33461_, _33460_, _35796_);
  or (_33462_, \oc8051_gm_cxrom_1.cell3.data [2], _35796_);
  and (_35813_[2], _33462_, _33461_);
  or (_33463_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33464_, \oc8051_gm_cxrom_1.cell3.data [3], _33443_);
  nand (_33465_, _33464_, _33463_);
  nand (_33466_, _33465_, _35796_);
  or (_33467_, \oc8051_gm_cxrom_1.cell3.data [3], _35796_);
  and (_35813_[3], _33467_, _33466_);
  or (_33468_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33469_, \oc8051_gm_cxrom_1.cell3.data [4], _33443_);
  nand (_33470_, _33469_, _33468_);
  nand (_33471_, _33470_, _35796_);
  or (_33472_, \oc8051_gm_cxrom_1.cell3.data [4], _35796_);
  and (_35813_[4], _33472_, _33471_);
  or (_33473_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33474_, \oc8051_gm_cxrom_1.cell3.data [5], _33443_);
  nand (_33475_, _33474_, _33473_);
  nand (_33476_, _33475_, _35796_);
  or (_33477_, \oc8051_gm_cxrom_1.cell3.data [5], _35796_);
  and (_35813_[5], _33477_, _33476_);
  or (_33478_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33479_, \oc8051_gm_cxrom_1.cell3.data [6], _33443_);
  nand (_33480_, _33479_, _33478_);
  nand (_33481_, _33480_, _35796_);
  or (_33482_, \oc8051_gm_cxrom_1.cell3.data [6], _35796_);
  and (_35813_[6], _33482_, _33481_);
  or (_33483_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_33484_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_33485_, _33484_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_33486_, _33485_, _33483_);
  nand (_33487_, _33486_, _35796_);
  or (_33488_, \oc8051_gm_cxrom_1.cell4.data [7], _35796_);
  and (_35815_[7], _33488_, _33487_);
  or (_33489_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33490_, \oc8051_gm_cxrom_1.cell4.data [0], _33484_);
  nand (_33491_, _33490_, _33489_);
  nand (_33492_, _33491_, _35796_);
  or (_33493_, \oc8051_gm_cxrom_1.cell4.data [0], _35796_);
  and (_35815_[0], _33493_, _33492_);
  or (_33494_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33495_, \oc8051_gm_cxrom_1.cell4.data [1], _33484_);
  nand (_33496_, _33495_, _33494_);
  nand (_33497_, _33496_, _35796_);
  or (_33498_, \oc8051_gm_cxrom_1.cell4.data [1], _35796_);
  and (_35815_[1], _33498_, _33497_);
  or (_33499_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33500_, \oc8051_gm_cxrom_1.cell4.data [2], _33484_);
  nand (_33501_, _33500_, _33499_);
  nand (_33502_, _33501_, _35796_);
  or (_33503_, \oc8051_gm_cxrom_1.cell4.data [2], _35796_);
  and (_35815_[2], _33503_, _33502_);
  or (_33504_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33505_, \oc8051_gm_cxrom_1.cell4.data [3], _33484_);
  nand (_33506_, _33505_, _33504_);
  nand (_33507_, _33506_, _35796_);
  or (_33508_, \oc8051_gm_cxrom_1.cell4.data [3], _35796_);
  and (_35815_[3], _33508_, _33507_);
  or (_33509_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33510_, \oc8051_gm_cxrom_1.cell4.data [4], _33484_);
  nand (_33511_, _33510_, _33509_);
  nand (_33512_, _33511_, _35796_);
  or (_33513_, \oc8051_gm_cxrom_1.cell4.data [4], _35796_);
  and (_35815_[4], _33513_, _33512_);
  or (_33514_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33515_, \oc8051_gm_cxrom_1.cell4.data [5], _33484_);
  nand (_33516_, _33515_, _33514_);
  nand (_33517_, _33516_, _35796_);
  or (_33518_, \oc8051_gm_cxrom_1.cell4.data [5], _35796_);
  and (_35815_[5], _33518_, _33517_);
  or (_33519_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33520_, \oc8051_gm_cxrom_1.cell4.data [6], _33484_);
  nand (_33521_, _33520_, _33519_);
  nand (_33522_, _33521_, _35796_);
  or (_33523_, \oc8051_gm_cxrom_1.cell4.data [6], _35796_);
  and (_35815_[6], _33523_, _33522_);
  or (_33524_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_33525_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_33526_, _33525_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_33527_, _33526_, _33524_);
  nand (_33528_, _33527_, _35796_);
  or (_33529_, \oc8051_gm_cxrom_1.cell5.data [7], _35796_);
  and (_35817_[7], _33529_, _33528_);
  or (_33530_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33531_, \oc8051_gm_cxrom_1.cell5.data [0], _33525_);
  nand (_33532_, _33531_, _33530_);
  nand (_33533_, _33532_, _35796_);
  or (_33534_, \oc8051_gm_cxrom_1.cell5.data [0], _35796_);
  and (_35817_[0], _33534_, _33533_);
  or (_33535_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33536_, \oc8051_gm_cxrom_1.cell5.data [1], _33525_);
  nand (_33537_, _33536_, _33535_);
  nand (_33538_, _33537_, _35796_);
  or (_33539_, \oc8051_gm_cxrom_1.cell5.data [1], _35796_);
  and (_35817_[1], _33539_, _33538_);
  or (_33540_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33541_, \oc8051_gm_cxrom_1.cell5.data [2], _33525_);
  nand (_33542_, _33541_, _33540_);
  nand (_33543_, _33542_, _35796_);
  or (_33544_, \oc8051_gm_cxrom_1.cell5.data [2], _35796_);
  and (_35817_[2], _33544_, _33543_);
  or (_33545_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33546_, \oc8051_gm_cxrom_1.cell5.data [3], _33525_);
  nand (_33547_, _33546_, _33545_);
  nand (_33548_, _33547_, _35796_);
  or (_33549_, \oc8051_gm_cxrom_1.cell5.data [3], _35796_);
  and (_35817_[3], _33549_, _33548_);
  or (_33550_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33551_, \oc8051_gm_cxrom_1.cell5.data [4], _33525_);
  nand (_33552_, _33551_, _33550_);
  nand (_33553_, _33552_, _35796_);
  or (_33554_, \oc8051_gm_cxrom_1.cell5.data [4], _35796_);
  and (_35817_[4], _33554_, _33553_);
  or (_33555_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33556_, \oc8051_gm_cxrom_1.cell5.data [5], _33525_);
  nand (_33557_, _33556_, _33555_);
  nand (_33558_, _33557_, _35796_);
  or (_33559_, \oc8051_gm_cxrom_1.cell5.data [5], _35796_);
  and (_35817_[5], _33559_, _33558_);
  or (_33560_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33561_, \oc8051_gm_cxrom_1.cell5.data [6], _33525_);
  nand (_33562_, _33561_, _33560_);
  nand (_33563_, _33562_, _35796_);
  or (_33564_, \oc8051_gm_cxrom_1.cell5.data [6], _35796_);
  and (_35817_[6], _33564_, _33563_);
  or (_33565_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_33566_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_33567_, _33566_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_33568_, _33567_, _33565_);
  nand (_33569_, _33568_, _35796_);
  or (_33570_, \oc8051_gm_cxrom_1.cell6.data [7], _35796_);
  and (_35819_[7], _33570_, _33569_);
  or (_33571_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33572_, \oc8051_gm_cxrom_1.cell6.data [0], _33566_);
  nand (_33573_, _33572_, _33571_);
  nand (_33574_, _33573_, _35796_);
  or (_33575_, \oc8051_gm_cxrom_1.cell6.data [0], _35796_);
  and (_35819_[0], _33575_, _33574_);
  or (_33576_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33577_, \oc8051_gm_cxrom_1.cell6.data [1], _33566_);
  nand (_33578_, _33577_, _33576_);
  nand (_33579_, _33578_, _35796_);
  or (_33580_, \oc8051_gm_cxrom_1.cell6.data [1], _35796_);
  and (_35819_[1], _33580_, _33579_);
  or (_33581_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33582_, \oc8051_gm_cxrom_1.cell6.data [2], _33566_);
  nand (_33583_, _33582_, _33581_);
  nand (_33584_, _33583_, _35796_);
  or (_33585_, \oc8051_gm_cxrom_1.cell6.data [2], _35796_);
  and (_35819_[2], _33585_, _33584_);
  or (_33586_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33587_, \oc8051_gm_cxrom_1.cell6.data [3], _33566_);
  nand (_33588_, _33587_, _33586_);
  nand (_33589_, _33588_, _35796_);
  or (_33590_, \oc8051_gm_cxrom_1.cell6.data [3], _35796_);
  and (_35819_[3], _33590_, _33589_);
  or (_33591_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33592_, \oc8051_gm_cxrom_1.cell6.data [4], _33566_);
  nand (_33593_, _33592_, _33591_);
  nand (_33594_, _33593_, _35796_);
  or (_33595_, \oc8051_gm_cxrom_1.cell6.data [4], _35796_);
  and (_35819_[4], _33595_, _33594_);
  or (_33596_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33597_, \oc8051_gm_cxrom_1.cell6.data [5], _33566_);
  nand (_33598_, _33597_, _33596_);
  nand (_33599_, _33598_, _35796_);
  or (_33600_, \oc8051_gm_cxrom_1.cell6.data [5], _35796_);
  and (_35819_[5], _33600_, _33599_);
  or (_33601_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33602_, \oc8051_gm_cxrom_1.cell6.data [6], _33566_);
  nand (_33603_, _33602_, _33601_);
  nand (_33604_, _33603_, _35796_);
  or (_33605_, \oc8051_gm_cxrom_1.cell6.data [6], _35796_);
  and (_35819_[6], _33605_, _33604_);
  or (_33606_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_33607_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_33608_, _33607_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_33609_, _33608_, _33606_);
  nand (_33610_, _33609_, _35796_);
  or (_33611_, \oc8051_gm_cxrom_1.cell7.data [7], _35796_);
  and (_35821_[7], _33611_, _33610_);
  or (_33612_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33613_, \oc8051_gm_cxrom_1.cell7.data [0], _33607_);
  nand (_33614_, _33613_, _33612_);
  nand (_33615_, _33614_, _35796_);
  or (_33616_, \oc8051_gm_cxrom_1.cell7.data [0], _35796_);
  and (_35821_[0], _33616_, _33615_);
  or (_33617_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33618_, \oc8051_gm_cxrom_1.cell7.data [1], _33607_);
  nand (_33619_, _33618_, _33617_);
  nand (_33620_, _33619_, _35796_);
  or (_33621_, \oc8051_gm_cxrom_1.cell7.data [1], _35796_);
  and (_35821_[1], _33621_, _33620_);
  or (_33622_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33623_, \oc8051_gm_cxrom_1.cell7.data [2], _33607_);
  nand (_33624_, _33623_, _33622_);
  nand (_33625_, _33624_, _35796_);
  or (_33626_, \oc8051_gm_cxrom_1.cell7.data [2], _35796_);
  and (_35821_[2], _33626_, _33625_);
  or (_33627_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33628_, \oc8051_gm_cxrom_1.cell7.data [3], _33607_);
  nand (_33629_, _33628_, _33627_);
  nand (_33630_, _33629_, _35796_);
  or (_33631_, \oc8051_gm_cxrom_1.cell7.data [3], _35796_);
  and (_35821_[3], _33631_, _33630_);
  or (_33632_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33633_, \oc8051_gm_cxrom_1.cell7.data [4], _33607_);
  nand (_33634_, _33633_, _33632_);
  nand (_33635_, _33634_, _35796_);
  or (_33636_, \oc8051_gm_cxrom_1.cell7.data [4], _35796_);
  and (_35821_[4], _33636_, _33635_);
  or (_33637_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33638_, \oc8051_gm_cxrom_1.cell7.data [5], _33607_);
  nand (_33639_, _33638_, _33637_);
  nand (_33640_, _33639_, _35796_);
  or (_33641_, \oc8051_gm_cxrom_1.cell7.data [5], _35796_);
  and (_35821_[5], _33641_, _33640_);
  or (_33642_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33643_, \oc8051_gm_cxrom_1.cell7.data [6], _33607_);
  nand (_33644_, _33643_, _33642_);
  nand (_33645_, _33644_, _35796_);
  or (_33646_, \oc8051_gm_cxrom_1.cell7.data [6], _35796_);
  and (_35821_[6], _33646_, _33645_);
  or (_33647_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_33648_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_33649_, _33648_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_33650_, _33649_, _33647_);
  nand (_33651_, _33650_, _35796_);
  or (_33652_, \oc8051_gm_cxrom_1.cell8.data [7], _35796_);
  and (_35823_[7], _33652_, _33651_);
  or (_33653_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33654_, \oc8051_gm_cxrom_1.cell8.data [0], _33648_);
  nand (_33655_, _33654_, _33653_);
  nand (_33656_, _33655_, _35796_);
  or (_33657_, \oc8051_gm_cxrom_1.cell8.data [0], _35796_);
  and (_35823_[0], _33657_, _33656_);
  or (_33658_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33659_, \oc8051_gm_cxrom_1.cell8.data [1], _33648_);
  nand (_33660_, _33659_, _33658_);
  nand (_33661_, _33660_, _35796_);
  or (_33662_, \oc8051_gm_cxrom_1.cell8.data [1], _35796_);
  and (_35823_[1], _33662_, _33661_);
  or (_33663_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33664_, \oc8051_gm_cxrom_1.cell8.data [2], _33648_);
  nand (_33665_, _33664_, _33663_);
  nand (_33666_, _33665_, _35796_);
  or (_33668_, \oc8051_gm_cxrom_1.cell8.data [2], _35796_);
  and (_35823_[2], _33668_, _33666_);
  or (_33669_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33670_, \oc8051_gm_cxrom_1.cell8.data [3], _33648_);
  nand (_33671_, _33670_, _33669_);
  nand (_33673_, _33671_, _35796_);
  or (_33674_, \oc8051_gm_cxrom_1.cell8.data [3], _35796_);
  and (_35823_[3], _33674_, _33673_);
  or (_33675_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33676_, \oc8051_gm_cxrom_1.cell8.data [4], _33648_);
  nand (_33678_, _33676_, _33675_);
  nand (_33679_, _33678_, _35796_);
  or (_33680_, \oc8051_gm_cxrom_1.cell8.data [4], _35796_);
  and (_35823_[4], _33680_, _33679_);
  or (_33681_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33683_, \oc8051_gm_cxrom_1.cell8.data [5], _33648_);
  nand (_33684_, _33683_, _33681_);
  nand (_33685_, _33684_, _35796_);
  or (_33686_, \oc8051_gm_cxrom_1.cell8.data [5], _35796_);
  and (_35823_[5], _33686_, _33685_);
  or (_33688_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33689_, \oc8051_gm_cxrom_1.cell8.data [6], _33648_);
  nand (_33690_, _33689_, _33688_);
  nand (_33691_, _33690_, _35796_);
  or (_33692_, \oc8051_gm_cxrom_1.cell8.data [6], _35796_);
  and (_35823_[6], _33692_, _33691_);
  or (_33694_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_33695_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_33696_, _33695_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_33697_, _33696_, _33694_);
  nand (_33699_, _33697_, _35796_);
  or (_33700_, \oc8051_gm_cxrom_1.cell9.data [7], _35796_);
  and (_35825_[7], _33700_, _33699_);
  or (_33702_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33703_, \oc8051_gm_cxrom_1.cell9.data [0], _33695_);
  nand (_33704_, _33703_, _33702_);
  nand (_33705_, _33704_, _35796_);
  or (_33706_, \oc8051_gm_cxrom_1.cell9.data [0], _35796_);
  and (_35825_[0], _33706_, _33705_);
  or (_33708_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33709_, \oc8051_gm_cxrom_1.cell9.data [1], _33695_);
  nand (_33710_, _33709_, _33708_);
  nand (_33712_, _33710_, _35796_);
  or (_33713_, \oc8051_gm_cxrom_1.cell9.data [1], _35796_);
  and (_35825_[1], _33713_, _33712_);
  or (_33715_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33716_, \oc8051_gm_cxrom_1.cell9.data [2], _33695_);
  nand (_33717_, _33716_, _33715_);
  nand (_33719_, _33717_, _35796_);
  or (_33720_, \oc8051_gm_cxrom_1.cell9.data [2], _35796_);
  and (_35825_[2], _33720_, _33719_);
  or (_33722_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33723_, \oc8051_gm_cxrom_1.cell9.data [3], _33695_);
  nand (_33724_, _33723_, _33722_);
  nand (_33726_, _33724_, _35796_);
  or (_33727_, \oc8051_gm_cxrom_1.cell9.data [3], _35796_);
  and (_35825_[3], _33727_, _33726_);
  or (_33729_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33730_, \oc8051_gm_cxrom_1.cell9.data [4], _33695_);
  nand (_33732_, _33730_, _33729_);
  nand (_33733_, _33732_, _35796_);
  or (_33734_, \oc8051_gm_cxrom_1.cell9.data [4], _35796_);
  and (_35825_[4], _33734_, _33733_);
  or (_33735_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33736_, \oc8051_gm_cxrom_1.cell9.data [5], _33695_);
  nand (_33737_, _33736_, _33735_);
  nand (_33739_, _33737_, _35796_);
  or (_33740_, \oc8051_gm_cxrom_1.cell9.data [5], _35796_);
  and (_35825_[5], _33740_, _33739_);
  or (_33742_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33743_, \oc8051_gm_cxrom_1.cell9.data [6], _33695_);
  nand (_33744_, _33743_, _33742_);
  nand (_33746_, _33744_, _35796_);
  or (_33747_, \oc8051_gm_cxrom_1.cell9.data [6], _35796_);
  and (_35825_[6], _33747_, _33746_);
  or (_33749_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_33750_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_33751_, _33750_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_33753_, _33751_, _33749_);
  nand (_33754_, _33753_, _35796_);
  or (_33755_, \oc8051_gm_cxrom_1.cell10.data [7], _35796_);
  and (_35799_[7], _33755_, _33754_);
  or (_33757_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33758_, \oc8051_gm_cxrom_1.cell10.data [0], _33750_);
  nand (_33760_, _33758_, _33757_);
  nand (_33761_, _33760_, _35796_);
  or (_33763_, \oc8051_gm_cxrom_1.cell10.data [0], _35796_);
  and (_35799_[0], _33763_, _33761_);
  or (_33764_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33765_, \oc8051_gm_cxrom_1.cell10.data [1], _33750_);
  nand (_33766_, _33765_, _33764_);
  nand (_33768_, _33766_, _35796_);
  or (_33769_, \oc8051_gm_cxrom_1.cell10.data [1], _35796_);
  and (_35799_[1], _33769_, _33768_);
  or (_33771_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33772_, \oc8051_gm_cxrom_1.cell10.data [2], _33750_);
  nand (_33773_, _33772_, _33771_);
  nand (_33775_, _33773_, _35796_);
  or (_33776_, \oc8051_gm_cxrom_1.cell10.data [2], _35796_);
  and (_35799_[2], _33776_, _33775_);
  or (_33778_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33779_, \oc8051_gm_cxrom_1.cell10.data [3], _33750_);
  nand (_33780_, _33779_, _33778_);
  nand (_33782_, _33780_, _35796_);
  or (_33783_, \oc8051_gm_cxrom_1.cell10.data [3], _35796_);
  and (_35799_[3], _33783_, _33782_);
  or (_33785_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33786_, \oc8051_gm_cxrom_1.cell10.data [4], _33750_);
  nand (_33787_, _33786_, _33785_);
  nand (_33789_, _33787_, _35796_);
  or (_33790_, \oc8051_gm_cxrom_1.cell10.data [4], _35796_);
  and (_35799_[4], _33790_, _33789_);
  or (_33792_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33793_, \oc8051_gm_cxrom_1.cell10.data [5], _33750_);
  nand (_33794_, _33793_, _33792_);
  nand (_33795_, _33794_, _35796_);
  or (_33796_, \oc8051_gm_cxrom_1.cell10.data [5], _35796_);
  and (_35799_[5], _33796_, _33795_);
  or (_33798_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33799_, \oc8051_gm_cxrom_1.cell10.data [6], _33750_);
  nand (_33800_, _33799_, _33798_);
  nand (_33801_, _33800_, _35796_);
  or (_33802_, \oc8051_gm_cxrom_1.cell10.data [6], _35796_);
  and (_35799_[6], _33802_, _33801_);
  or (_33803_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_33804_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_33805_, _33804_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_33806_, _33805_, _33803_);
  nand (_33807_, _33806_, _35796_);
  or (_33808_, \oc8051_gm_cxrom_1.cell11.data [7], _35796_);
  and (_35801_[7], _33808_, _33807_);
  or (_33809_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33810_, \oc8051_gm_cxrom_1.cell11.data [0], _33804_);
  nand (_33811_, _33810_, _33809_);
  nand (_33812_, _33811_, _35796_);
  or (_33813_, \oc8051_gm_cxrom_1.cell11.data [0], _35796_);
  and (_35801_[0], _33813_, _33812_);
  or (_33814_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33815_, \oc8051_gm_cxrom_1.cell11.data [1], _33804_);
  nand (_33816_, _33815_, _33814_);
  nand (_33817_, _33816_, _35796_);
  or (_33818_, \oc8051_gm_cxrom_1.cell11.data [1], _35796_);
  and (_35801_[1], _33818_, _33817_);
  or (_33819_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33820_, \oc8051_gm_cxrom_1.cell11.data [2], _33804_);
  nand (_33821_, _33820_, _33819_);
  nand (_33822_, _33821_, _35796_);
  or (_33823_, \oc8051_gm_cxrom_1.cell11.data [2], _35796_);
  and (_35801_[2], _33823_, _33822_);
  or (_33824_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33825_, \oc8051_gm_cxrom_1.cell11.data [3], _33804_);
  nand (_33826_, _33825_, _33824_);
  nand (_33827_, _33826_, _35796_);
  or (_33828_, \oc8051_gm_cxrom_1.cell11.data [3], _35796_);
  and (_35801_[3], _33828_, _33827_);
  or (_33829_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33830_, \oc8051_gm_cxrom_1.cell11.data [4], _33804_);
  nand (_33831_, _33830_, _33829_);
  nand (_33832_, _33831_, _35796_);
  or (_33833_, \oc8051_gm_cxrom_1.cell11.data [4], _35796_);
  and (_35801_[4], _33833_, _33832_);
  or (_33834_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33835_, \oc8051_gm_cxrom_1.cell11.data [5], _33804_);
  nand (_33836_, _33835_, _33834_);
  nand (_33837_, _33836_, _35796_);
  or (_33838_, \oc8051_gm_cxrom_1.cell11.data [5], _35796_);
  and (_35801_[5], _33838_, _33837_);
  or (_33839_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33840_, \oc8051_gm_cxrom_1.cell11.data [6], _33804_);
  nand (_33841_, _33840_, _33839_);
  nand (_33842_, _33841_, _35796_);
  or (_33843_, \oc8051_gm_cxrom_1.cell11.data [6], _35796_);
  and (_35801_[6], _33843_, _33842_);
  or (_33844_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_33845_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_33846_, _33845_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_33847_, _33846_, _33844_);
  nand (_33848_, _33847_, _35796_);
  or (_33849_, \oc8051_gm_cxrom_1.cell12.data [7], _35796_);
  and (_35803_[7], _33849_, _33848_);
  or (_33850_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33851_, \oc8051_gm_cxrom_1.cell12.data [0], _33845_);
  nand (_33852_, _33851_, _33850_);
  nand (_33853_, _33852_, _35796_);
  or (_33854_, \oc8051_gm_cxrom_1.cell12.data [0], _35796_);
  and (_35803_[0], _33854_, _33853_);
  or (_33855_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33856_, \oc8051_gm_cxrom_1.cell12.data [1], _33845_);
  nand (_33857_, _33856_, _33855_);
  nand (_33858_, _33857_, _35796_);
  or (_33859_, \oc8051_gm_cxrom_1.cell12.data [1], _35796_);
  and (_35803_[1], _33859_, _33858_);
  or (_33860_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33861_, \oc8051_gm_cxrom_1.cell12.data [2], _33845_);
  nand (_33862_, _33861_, _33860_);
  nand (_33863_, _33862_, _35796_);
  or (_33864_, \oc8051_gm_cxrom_1.cell12.data [2], _35796_);
  and (_35803_[2], _33864_, _33863_);
  or (_33865_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33866_, \oc8051_gm_cxrom_1.cell12.data [3], _33845_);
  nand (_33867_, _33866_, _33865_);
  nand (_33868_, _33867_, _35796_);
  or (_33869_, \oc8051_gm_cxrom_1.cell12.data [3], _35796_);
  and (_35803_[3], _33869_, _33868_);
  or (_33870_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33871_, \oc8051_gm_cxrom_1.cell12.data [4], _33845_);
  nand (_33872_, _33871_, _33870_);
  nand (_33873_, _33872_, _35796_);
  or (_33874_, \oc8051_gm_cxrom_1.cell12.data [4], _35796_);
  and (_35803_[4], _33874_, _33873_);
  or (_33875_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33876_, \oc8051_gm_cxrom_1.cell12.data [5], _33845_);
  nand (_33877_, _33876_, _33875_);
  nand (_33878_, _33877_, _35796_);
  or (_33879_, \oc8051_gm_cxrom_1.cell12.data [5], _35796_);
  and (_35803_[5], _33879_, _33878_);
  or (_33880_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33881_, \oc8051_gm_cxrom_1.cell12.data [6], _33845_);
  nand (_33882_, _33881_, _33880_);
  nand (_33883_, _33882_, _35796_);
  or (_33884_, \oc8051_gm_cxrom_1.cell12.data [6], _35796_);
  and (_35803_[6], _33884_, _33883_);
  or (_33885_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_33886_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_33887_, _33886_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_33888_, _33887_, _33885_);
  nand (_33889_, _33888_, _35796_);
  or (_33890_, \oc8051_gm_cxrom_1.cell13.data [7], _35796_);
  and (_35805_[7], _33890_, _33889_);
  or (_33891_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33892_, \oc8051_gm_cxrom_1.cell13.data [0], _33886_);
  nand (_33893_, _33892_, _33891_);
  nand (_33894_, _33893_, _35796_);
  or (_33895_, \oc8051_gm_cxrom_1.cell13.data [0], _35796_);
  and (_35805_[0], _33895_, _33894_);
  or (_33896_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33897_, \oc8051_gm_cxrom_1.cell13.data [1], _33886_);
  nand (_33898_, _33897_, _33896_);
  nand (_33899_, _33898_, _35796_);
  or (_33900_, \oc8051_gm_cxrom_1.cell13.data [1], _35796_);
  and (_35805_[1], _33900_, _33899_);
  or (_33901_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33902_, \oc8051_gm_cxrom_1.cell13.data [2], _33886_);
  nand (_33903_, _33902_, _33901_);
  nand (_33904_, _33903_, _35796_);
  or (_33905_, \oc8051_gm_cxrom_1.cell13.data [2], _35796_);
  and (_35805_[2], _33905_, _33904_);
  or (_33906_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33907_, \oc8051_gm_cxrom_1.cell13.data [3], _33886_);
  nand (_33908_, _33907_, _33906_);
  nand (_33909_, _33908_, _35796_);
  or (_33910_, \oc8051_gm_cxrom_1.cell13.data [3], _35796_);
  and (_35805_[3], _33910_, _33909_);
  or (_33911_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33912_, \oc8051_gm_cxrom_1.cell13.data [4], _33886_);
  nand (_33913_, _33912_, _33911_);
  nand (_33914_, _33913_, _35796_);
  or (_33915_, \oc8051_gm_cxrom_1.cell13.data [4], _35796_);
  and (_35805_[4], _33915_, _33914_);
  or (_33916_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33917_, \oc8051_gm_cxrom_1.cell13.data [5], _33886_);
  nand (_33918_, _33917_, _33916_);
  nand (_33919_, _33918_, _35796_);
  or (_33920_, \oc8051_gm_cxrom_1.cell13.data [5], _35796_);
  and (_35805_[5], _33920_, _33919_);
  or (_33921_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33922_, \oc8051_gm_cxrom_1.cell13.data [6], _33886_);
  nand (_33923_, _33922_, _33921_);
  nand (_33924_, _33923_, _35796_);
  or (_33925_, \oc8051_gm_cxrom_1.cell13.data [6], _35796_);
  and (_35805_[6], _33925_, _33924_);
  or (_33926_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_33927_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_33928_, _33927_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_33929_, _33928_, _33926_);
  nand (_33930_, _33929_, _35796_);
  or (_33931_, \oc8051_gm_cxrom_1.cell14.data [7], _35796_);
  and (_35807_[7], _33931_, _33930_);
  or (_33932_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33933_, \oc8051_gm_cxrom_1.cell14.data [0], _33927_);
  nand (_33934_, _33933_, _33932_);
  nand (_33935_, _33934_, _35796_);
  or (_33936_, \oc8051_gm_cxrom_1.cell14.data [0], _35796_);
  and (_35807_[0], _33936_, _33935_);
  or (_33937_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33938_, \oc8051_gm_cxrom_1.cell14.data [1], _33927_);
  nand (_33939_, _33938_, _33937_);
  nand (_33940_, _33939_, _35796_);
  or (_33941_, \oc8051_gm_cxrom_1.cell14.data [1], _35796_);
  and (_35807_[1], _33941_, _33940_);
  or (_33942_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33943_, \oc8051_gm_cxrom_1.cell14.data [2], _33927_);
  nand (_33944_, _33943_, _33942_);
  nand (_33945_, _33944_, _35796_);
  or (_33946_, \oc8051_gm_cxrom_1.cell14.data [2], _35796_);
  and (_35807_[2], _33946_, _33945_);
  or (_33947_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33948_, \oc8051_gm_cxrom_1.cell14.data [3], _33927_);
  nand (_33949_, _33948_, _33947_);
  nand (_33950_, _33949_, _35796_);
  or (_33951_, \oc8051_gm_cxrom_1.cell14.data [3], _35796_);
  and (_35807_[3], _33951_, _33950_);
  or (_33952_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33953_, \oc8051_gm_cxrom_1.cell14.data [4], _33927_);
  nand (_33954_, _33953_, _33952_);
  nand (_33955_, _33954_, _35796_);
  or (_33956_, \oc8051_gm_cxrom_1.cell14.data [4], _35796_);
  and (_35807_[4], _33956_, _33955_);
  or (_33957_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33958_, \oc8051_gm_cxrom_1.cell14.data [5], _33927_);
  nand (_33959_, _33958_, _33957_);
  nand (_33960_, _33959_, _35796_);
  or (_33961_, \oc8051_gm_cxrom_1.cell14.data [5], _35796_);
  and (_35807_[5], _33961_, _33960_);
  or (_33962_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33963_, \oc8051_gm_cxrom_1.cell14.data [6], _33927_);
  nand (_33964_, _33963_, _33962_);
  nand (_33965_, _33964_, _35796_);
  or (_33966_, \oc8051_gm_cxrom_1.cell14.data [6], _35796_);
  and (_35807_[6], _33966_, _33965_);
  or (_33967_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_33968_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_33969_, _33968_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_33970_, _33969_, _33967_);
  nand (_33971_, _33970_, _35796_);
  or (_33972_, \oc8051_gm_cxrom_1.cell15.data [7], _35796_);
  and (_35809_[7], _33972_, _33971_);
  or (_33973_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33974_, \oc8051_gm_cxrom_1.cell15.data [0], _33968_);
  nand (_33975_, _33974_, _33973_);
  nand (_33976_, _33975_, _35796_);
  or (_33977_, \oc8051_gm_cxrom_1.cell15.data [0], _35796_);
  and (_35809_[0], _33977_, _33976_);
  or (_33978_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33979_, \oc8051_gm_cxrom_1.cell15.data [1], _33968_);
  nand (_33980_, _33979_, _33978_);
  nand (_33981_, _33980_, _35796_);
  or (_33982_, \oc8051_gm_cxrom_1.cell15.data [1], _35796_);
  and (_35809_[1], _33982_, _33981_);
  or (_33983_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33984_, \oc8051_gm_cxrom_1.cell15.data [2], _33968_);
  nand (_33985_, _33984_, _33983_);
  nand (_33986_, _33985_, _35796_);
  or (_33987_, \oc8051_gm_cxrom_1.cell15.data [2], _35796_);
  and (_35809_[2], _33987_, _33986_);
  or (_33988_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33989_, \oc8051_gm_cxrom_1.cell15.data [3], _33968_);
  nand (_33990_, _33989_, _33988_);
  nand (_33991_, _33990_, _35796_);
  or (_33992_, \oc8051_gm_cxrom_1.cell15.data [3], _35796_);
  and (_35809_[3], _33992_, _33991_);
  or (_33993_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33994_, \oc8051_gm_cxrom_1.cell15.data [4], _33968_);
  nand (_33995_, _33994_, _33993_);
  nand (_33996_, _33995_, _35796_);
  or (_33997_, \oc8051_gm_cxrom_1.cell15.data [4], _35796_);
  and (_35809_[4], _33997_, _33996_);
  or (_33998_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33999_, \oc8051_gm_cxrom_1.cell15.data [5], _33968_);
  nand (_34000_, _33999_, _33998_);
  nand (_34001_, _34000_, _35796_);
  or (_34002_, \oc8051_gm_cxrom_1.cell15.data [5], _35796_);
  and (_35809_[5], _34002_, _34001_);
  or (_34003_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_34004_, \oc8051_gm_cxrom_1.cell15.data [6], _33968_);
  nand (_34005_, _34004_, _34003_);
  nand (_34006_, _34005_, _35796_);
  or (_34007_, \oc8051_gm_cxrom_1.cell15.data [6], _35796_);
  and (_35809_[6], _34007_, _34006_);
  nor (_35986_[2], _30743_, rst);
  and (_34008_, _30494_, _35796_);
  nand (_34009_, _34008_, _30784_);
  nor (_34010_, _30735_, _30705_);
  or (_35987_[2], _34010_, _34009_);
  not (_34011_, _30527_);
  nor (_34012_, _30699_, _34011_);
  nor (_34013_, _30550_, _30574_);
  and (_34014_, _34013_, _30597_);
  and (_34015_, _34014_, _34012_);
  not (_34016_, _30597_);
  not (_34017_, _30574_);
  nor (_34018_, _30550_, _34017_);
  and (_34019_, _34018_, _34016_);
  not (_34020_, _30676_);
  and (_34021_, _30699_, _34020_);
  nor (_34022_, _30649_, _34011_);
  and (_34023_, _34022_, _34021_);
  or (_34024_, _34023_, _34012_);
  and (_34025_, _34024_, _34019_);
  or (_34026_, _34025_, _34015_);
  and (_34027_, _34021_, _30649_);
  nor (_34028_, _30597_, _34011_);
  and (_34029_, _34028_, _34018_);
  and (_34030_, _34029_, _34027_);
  not (_34031_, _30649_);
  and (_34032_, _30699_, _30676_);
  and (_34033_, _34032_, _34031_);
  and (_34034_, _34033_, _30624_);
  and (_34035_, _30550_, _30574_);
  and (_34036_, _34035_, _30597_);
  and (_34037_, _34036_, _34034_);
  or (_34038_, _34037_, _34030_);
  or (_34039_, _34038_, _34026_);
  and (_34040_, _30649_, _30624_);
  and (_34041_, _34040_, _34021_);
  and (_34042_, _34041_, _34011_);
  and (_34043_, _34042_, _34018_);
  and (_34044_, _34013_, _34016_);
  and (_34045_, _34044_, _34033_);
  or (_34046_, _34045_, _34043_);
  or (_34047_, _34046_, _34039_);
  not (_34048_, _30624_);
  nor (_34049_, _30597_, _30527_);
  and (_34050_, _30550_, _34017_);
  and (_34051_, _34050_, _34049_);
  nor (_34052_, _34051_, _34048_);
  and (_34053_, _34032_, _30649_);
  not (_34054_, _34053_);
  nor (_34055_, _34054_, _34052_);
  not (_34056_, _34055_);
  and (_34057_, _34040_, _34032_);
  and (_34058_, _34035_, _34028_);
  and (_34059_, _34058_, _34057_);
  and (_34060_, _30597_, _34011_);
  and (_34061_, _34050_, _34060_);
  and (_34062_, _34061_, _34057_);
  nor (_34063_, _34062_, _34059_);
  and (_34064_, _34063_, _34056_);
  and (_34065_, _34060_, _34018_);
  and (_34066_, _34057_, _34065_);
  and (_34067_, _34018_, _30597_);
  and (_34068_, _34033_, _34048_);
  and (_34069_, _34068_, _34067_);
  or (_34070_, _34069_, _34066_);
  and (_34071_, _30597_, _30527_);
  or (_34072_, _34049_, _34071_);
  and (_34073_, _34072_, _34035_);
  and (_34074_, _34073_, _34057_);
  and (_34075_, _34035_, _34016_);
  and (_34076_, _34075_, _34034_);
  or (_34077_, _34076_, _34074_);
  or (_34078_, _34077_, _34070_);
  and (_34079_, _34050_, _34028_);
  and (_34080_, _34079_, _34068_);
  and (_34081_, _34071_, _34013_);
  and (_34082_, _34027_, _34048_);
  and (_34083_, _34082_, _34081_);
  or (_34084_, _34083_, _34080_);
  and (_34085_, _34050_, _30527_);
  and (_34086_, _34085_, _34057_);
  and (_34087_, _34057_, _34044_);
  or (_34088_, _34087_, _34086_);
  or (_34089_, _34088_, _34084_);
  nor (_34090_, _34089_, _34078_);
  nand (_34091_, _34090_, _34064_);
  or (_34092_, _34091_, _34047_);
  and (_34093_, _34092_, _30495_);
  not (_34094_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_34095_, _30493_, _15260_);
  and (_34096_, _34095_, _30731_);
  nor (_34097_, _34096_, _34094_);
  or (_34098_, _34097_, rst);
  or (_35988_[1], _34098_, _34093_);
  nand (_34099_, _30550_, _30489_);
  or (_34100_, _30489_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_34101_, _34100_, _35796_);
  and (_35989_[7], _34101_, _34099_);
  and (_34102_, \oc8051_top_1.oc8051_sfr1.wait_data , _35796_);
  and (_34103_, _34102_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_34104_, _30736_, _30809_);
  and (_34105_, _30798_, _30705_);
  and (_34106_, _30735_, _30720_);
  or (_34107_, _34106_, _34105_);
  and (_34108_, _30706_, _30767_);
  or (_34109_, _34108_, _34107_);
  or (_34110_, _34109_, _34104_);
  not (_34111_, _30783_);
  and (_34112_, _30724_, _30785_);
  and (_34113_, _30706_, _30712_);
  and (_34114_, _34113_, _30532_);
  or (_34115_, _34114_, _34112_);
  or (_34116_, _34115_, _34111_);
  or (_34117_, _34116_, _34110_);
  and (_34118_, _34117_, _34008_);
  or (_35990_, _34118_, _34103_);
  and (_34119_, _30735_, _30713_);
  or (_34120_, _34119_, _30707_);
  nor (_34121_, _30703_, _30709_);
  and (_34122_, _30765_, _34121_);
  and (_34123_, _34122_, _30555_);
  or (_34124_, _34123_, _30860_);
  and (_34125_, _30722_, _30655_);
  and (_34126_, _34125_, _30767_);
  or (_34127_, _34126_, _34124_);
  or (_34128_, _34127_, _34120_);
  and (_34129_, _34128_, _30494_);
  and (_34130_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34131_, \oc8051_top_1.oc8051_decoder1.state [0], _15260_);
  and (_34132_, _34131_, _34094_);
  not (_34133_, _30727_);
  and (_34134_, _34133_, _34132_);
  or (_34135_, _34134_, _34130_);
  or (_34136_, _34135_, _34129_);
  and (_35991_[1], _34136_, _35796_);
  and (_34137_, _34102_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_34138_, _30724_, _30788_);
  nor (_34139_, _30798_, _30788_);
  nor (_34140_, _34139_, _30823_);
  or (_34141_, _34140_, _34138_);
  and (_34142_, _34125_, _30780_);
  or (_34143_, _34142_, _34141_);
  not (_34144_, _30856_);
  nor (_34145_, _34139_, _30703_);
  nor (_34146_, _30703_, _30532_);
  and (_34147_, _34146_, _30779_);
  or (_34148_, _34147_, _34145_);
  or (_34149_, _34148_, _34144_);
  and (_34150_, _30724_, _30820_);
  and (_34151_, _30807_, _30756_);
  or (_34152_, _34151_, _34120_);
  or (_34153_, _34152_, _34150_);
  or (_34154_, _34153_, _34149_);
  or (_34155_, _34154_, _34143_);
  and (_34156_, _34155_, _34008_);
  or (_35992_[1], _34156_, _34137_);
  and (_34157_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34158_, _30751_, _30494_);
  or (_34159_, _34158_, _34157_);
  or (_34160_, _34159_, _34134_);
  and (_35993_[2], _34160_, _35796_);
  not (_34161_, _34010_);
  and (_34162_, _34161_, _30785_);
  nor (_34163_, _34162_, _34113_);
  not (_34164_, _34163_);
  and (_34165_, _34164_, _34132_);
  or (_34166_, _34165_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34167_, _30749_, _30704_);
  and (_34168_, _30779_, _30747_);
  nor (_34169_, _34168_, _34167_);
  nor (_34170_, _34169_, _30532_);
  not (_34171_, _30490_);
  and (_34172_, _34114_, _34171_);
  or (_34173_, _34172_, _34170_);
  and (_34174_, _34173_, _30731_);
  or (_34175_, _34174_, _34166_);
  or (_34176_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _15260_);
  and (_34177_, _34176_, _35796_);
  and (_35994_[2], _34177_, _34175_);
  and (_34178_, _34102_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_34179_, _34146_, _30766_);
  or (_34180_, _34179_, _34147_);
  or (_34181_, _30707_, _30799_);
  or (_34182_, _34181_, _34180_);
  or (_34183_, _34142_, _34105_);
  and (_34184_, _30791_, _30767_);
  and (_34185_, _30791_, _30780_);
  or (_34186_, _34185_, _34184_);
  or (_34187_, _34186_, _34183_);
  or (_34188_, _30827_, _30808_);
  or (_34189_, _34123_, _30768_);
  or (_34190_, _34189_, _34188_);
  or (_34191_, _34190_, _34187_);
  or (_34192_, _34191_, _34182_);
  and (_34193_, _34192_, _34008_);
  or (_35995_[1], _34193_, _34178_);
  and (_34194_, _34102_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  nand (_34195_, _30724_, _30802_);
  nand (_34196_, _34195_, _30813_);
  and (_34197_, _30853_, _30766_);
  and (_34198_, _30792_, _30765_);
  or (_34199_, _34198_, _30868_);
  or (_34200_, _34199_, _34197_);
  or (_34201_, _34200_, _34148_);
  or (_34202_, _34201_, _34196_);
  nor (_34203_, _30855_, _30817_);
  nand (_34204_, _34203_, _30805_);
  and (_34205_, _34125_, _30770_);
  or (_34206_, _34205_, _34126_);
  and (_34207_, _30715_, _34121_);
  or (_34208_, _34207_, _34122_);
  and (_34209_, _30706_, _30753_);
  or (_34210_, _34209_, _34208_);
  or (_34211_, _34210_, _34206_);
  or (_34212_, _34211_, _34204_);
  or (_34213_, _34212_, _34143_);
  or (_34214_, _34213_, _34202_);
  and (_34215_, _34214_, _34008_);
  or (_35996_[3], _34215_, _34194_);
  and (_34216_, _34146_, _30712_);
  and (_34217_, _30791_, _30754_);
  and (_34218_, _34125_, _30754_);
  or (_34219_, _34218_, _34217_);
  or (_34220_, _34219_, _34216_);
  and (_34221_, _30754_, _30756_);
  or (_34222_, _34221_, _30861_);
  or (_34223_, _34222_, _34220_);
  and (_34224_, _34125_, _30713_);
  or (_34225_, _34224_, _34223_);
  and (_34226_, _34225_, _30494_);
  nand (_34227_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_34228_, _34227_, _30740_);
  or (_34229_, _34228_, _34226_);
  and (_35997_[1], _34229_, _35796_);
  or (_34230_, _30826_, _30768_);
  or (_34231_, _34140_, _30819_);
  or (_34232_, _34231_, _34230_);
  or (_34233_, _30812_, _30800_);
  and (_34234_, _30780_, _30747_);
  and (_34235_, _30750_, _30709_);
  and (_34236_, _34235_, _30714_);
  or (_34237_, _34236_, _34234_);
  or (_34238_, _34237_, _34233_);
  nand (_34239_, _30810_, _30752_);
  or (_34240_, _34239_, _34238_);
  or (_34241_, _34240_, _34232_);
  and (_34242_, _30853_, _30714_);
  or (_34243_, _34242_, _30855_);
  or (_34244_, _34243_, _30793_);
  and (_34245_, _34146_, _30714_);
  or (_34246_, _34245_, _30757_);
  or (_34247_, _34246_, _34124_);
  or (_34248_, _34247_, _34244_);
  and (_34249_, _34167_, _30709_);
  or (_34250_, _34249_, _30857_);
  and (_34251_, _30720_, _30756_);
  or (_34252_, _34251_, _30763_);
  or (_34253_, _34252_, _34250_);
  or (_34254_, _34253_, _34148_);
  or (_34255_, _34254_, _34248_);
  or (_34256_, _34255_, _34241_);
  and (_34257_, _34256_, _30494_);
  and (_34258_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34259_, _30733_, _30841_);
  or (_34260_, _34234_, _34249_);
  and (_34261_, _34260_, _30733_);
  or (_34262_, _34261_, _34134_);
  or (_34263_, _34262_, _34259_);
  or (_34264_, _34263_, _34258_);
  or (_34265_, _34264_, _34257_);
  and (_35998_, _34265_, _35796_);
  nor (_35986_[0], _30884_, rst);
  nor (_35986_[1], _30848_, rst);
  nand (_35987_[0], _34164_, _34008_);
  nand (_34266_, _34008_, _34113_);
  or (_34267_, _34009_, _30777_);
  and (_35987_[1], _34267_, _34266_);
  or (_34268_, _34069_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_34269_, _34268_, _34076_);
  or (_34270_, _34269_, _34043_);
  and (_34271_, _34270_, _34096_);
  nor (_34272_, _34095_, _30731_);
  or (_34273_, _34272_, rst);
  or (_35988_[0], _34273_, _34271_);
  nand (_34274_, _30624_, _30489_);
  or (_34275_, _30489_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_34276_, _34275_, _35796_);
  and (_35989_[0], _34276_, _34274_);
  nand (_34277_, _30649_, _30489_);
  or (_34278_, _30489_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_34279_, _34278_, _35796_);
  and (_35989_[1], _34279_, _34277_);
  nand (_34280_, _30676_, _30489_);
  or (_34281_, _30489_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_34282_, _34281_, _35796_);
  and (_35989_[2], _34282_, _34280_);
  nand (_34283_, _30699_, _30489_);
  or (_34284_, _30489_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_34285_, _34284_, _35796_);
  and (_35989_[3], _34285_, _34283_);
  nand (_34286_, _34011_, _30489_);
  or (_34287_, _30489_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_34288_, _34287_, _35796_);
  and (_35989_[4], _34288_, _34286_);
  nand (_34289_, _30597_, _30489_);
  or (_34290_, _30489_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_34291_, _34290_, _35796_);
  and (_35989_[5], _34291_, _34289_);
  nand (_34292_, _30574_, _30489_);
  or (_34293_, _30489_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_34294_, _34293_, _35796_);
  and (_35989_[6], _34294_, _34292_);
  or (_34295_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _15260_);
  and (_34296_, _34295_, _34166_);
  and (_34297_, _34125_, _30802_);
  or (_34298_, _34297_, _34119_);
  or (_34299_, _34298_, _34220_);
  and (_34300_, _34146_, _30761_);
  or (_34301_, _34300_, _34221_);
  or (_34302_, _30798_, _30779_);
  and (_34303_, _34302_, _30724_);
  or (_34304_, _34303_, _34301_);
  or (_34305_, _34304_, _34299_);
  or (_34306_, _34112_, _30786_);
  or (_34307_, _30873_, _30868_);
  or (_34308_, _34307_, _34306_);
  and (_34309_, _30784_, _34121_);
  and (_34310_, _30761_, _34121_);
  or (_34311_, _34310_, _34207_);
  or (_34312_, _34311_, _34309_);
  and (_34313_, _30791_, _30713_);
  or (_34314_, _30707_, _34313_);
  or (_34315_, _34314_, _34312_);
  or (_34316_, _34315_, _34308_);
  and (_34317_, _30724_, _30716_);
  and (_34318_, _30784_, _30709_);
  and (_34319_, _34318_, _30724_);
  and (_34320_, _34125_, _30762_);
  or (_34321_, _34320_, _34319_);
  or (_34322_, _34321_, _34317_);
  or (_34323_, _34209_, _34205_);
  and (_34324_, _30791_, _30762_);
  or (_34325_, _34324_, _34224_);
  or (_34326_, _34325_, _34323_);
  or (_34327_, _34326_, _34322_);
  or (_34328_, _34327_, _34316_);
  or (_34329_, _34328_, _34305_);
  and (_34330_, _34329_, _30494_);
  or (_34331_, _34330_, _34296_);
  and (_35991_[0], _34331_, _35796_);
  and (_34332_, _34102_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_34333_, _30769_, _30747_);
  nor (_34334_, _34333_, _34208_);
  nand (_34335_, _34334_, _30772_);
  and (_34336_, _34146_, _30603_);
  and (_34337_, _34336_, _30555_);
  nor (_34338_, _34337_, _30854_);
  not (_34339_, _34338_);
  or (_34340_, _34339_, _34298_);
  or (_34341_, _34340_, _34335_);
  or (_34342_, _34200_, _34115_);
  or (_34343_, _34342_, _34341_);
  not (_34344_, _30770_);
  nand (_34345_, _30824_, _34344_);
  or (_34346_, _34345_, _30820_);
  and (_34347_, _34346_, _30724_);
  or (_34348_, _34347_, _34343_);
  and (_34349_, _34348_, _34008_);
  or (_35992_[0], _34349_, _34332_);
  or (_34350_, _34253_, _34241_);
  and (_34351_, _34350_, _30494_);
  and (_34352_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34353_, _34352_, _34263_);
  or (_34354_, _34353_, _34351_);
  and (_35993_[0], _34354_, _35796_);
  and (_34355_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34356_, _34355_, _34262_);
  and (_34357_, _34356_, _35796_);
  and (_34358_, _30816_, _30532_);
  or (_34359_, _34358_, _30860_);
  or (_34360_, _34359_, _34244_);
  or (_34361_, _34360_, _34170_);
  and (_34362_, _34361_, _34008_);
  or (_35993_[1], _34362_, _34357_);
  or (_34363_, _30726_, _34113_);
  and (_34364_, _34218_, _30709_);
  or (_34365_, _34364_, _34320_);
  or (_34366_, _34365_, _34363_);
  or (_34367_, _34216_, _30865_);
  or (_34368_, _34367_, _34170_);
  or (_34369_, _34368_, _34366_);
  and (_34370_, _34125_, _30807_);
  or (_34371_, _34370_, _34112_);
  or (_34372_, _34319_, _30725_);
  or (_34373_, _34372_, _34303_);
  or (_34374_, _34373_, _34371_);
  and (_34375_, _30724_, _30767_);
  or (_34376_, _34224_, _34209_);
  or (_34377_, _34376_, _34375_);
  or (_34378_, _34377_, _34301_);
  and (_34379_, _30762_, _30747_);
  and (_34380_, _34218_, _30532_);
  or (_34381_, _34380_, _34379_);
  and (_34382_, _30706_, _30716_);
  and (_34383_, _34235_, _30784_);
  or (_34384_, _34383_, _34382_);
  or (_34385_, _34384_, _34381_);
  and (_34386_, _30724_, _30769_);
  or (_34387_, _34245_, _34242_);
  or (_34388_, _34387_, _34386_);
  or (_34389_, _34317_, _34313_);
  or (_34390_, _34389_, _34388_);
  or (_34391_, _34390_, _34385_);
  or (_34392_, _34391_, _34378_);
  or (_34393_, _34392_, _34374_);
  or (_34394_, _34393_, _34369_);
  and (_34395_, _34394_, _30494_);
  and (_34396_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34397_, _34165_, _30741_);
  or (_34398_, _34397_, _34396_);
  or (_34399_, _34398_, _34395_);
  and (_35994_[0], _34399_, _35796_);
  and (_34400_, _34245_, _30555_);
  or (_34401_, _34400_, _34313_);
  or (_34402_, _30726_, _30763_);
  or (_34403_, _34402_, _34401_);
  or (_34404_, _30718_, _30825_);
  or (_34405_, _34404_, _34403_);
  or (_34406_, _34236_, _34119_);
  and (_34407_, _30853_, _30784_);
  and (_34408_, _30706_, _30769_);
  or (_34409_, _34408_, _34407_);
  or (_34410_, _34409_, _34406_);
  or (_34411_, _34410_, _34367_);
  or (_34412_, _34411_, _34405_);
  or (_34413_, _34378_, _34374_);
  or (_34414_, _34413_, _34412_);
  and (_34415_, _34414_, _30494_);
  or (_34416_, _34415_, _34397_);
  and (_34417_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34418_, _34417_, _34416_);
  and (_35994_[1], _34418_, _35796_);
  and (_34419_, _34102_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_34420_, _34336_, _30554_);
  and (_34421_, _30706_, _30807_);
  or (_34422_, _34421_, _34420_);
  and (_34423_, _30706_, _30778_);
  or (_34424_, _34423_, _34422_);
  or (_34425_, _34424_, _34182_);
  and (_34426_, _30706_, _30779_);
  and (_34427_, _34426_, _30709_);
  and (_34428_, _34105_, _30629_);
  or (_34429_, _34428_, _34427_);
  not (_34430_, _32137_);
  or (_34431_, _34224_, _34430_);
  or (_34432_, _34431_, _34429_);
  or (_34433_, _34432_, _34425_);
  or (_34434_, _34216_, _34123_);
  and (_34435_, _30724_, _30798_);
  or (_34436_, _34435_, _34142_);
  or (_34437_, _34436_, _34230_);
  or (_34438_, _34437_, _34434_);
  and (_34439_, _34217_, _30709_);
  or (_34440_, _34439_, _34364_);
  or (_34441_, _34440_, _34186_);
  nor (_34442_, _34313_, _30748_);
  nand (_34443_, _34442_, _32135_);
  or (_34444_, _34443_, _34441_);
  or (_34445_, _34444_, _34438_);
  or (_34446_, _34445_, _34433_);
  and (_34447_, _34446_, _34008_);
  or (_35995_[0], _34447_, _34419_);
  or (_34448_, _34198_, _34197_);
  or (_34449_, _34380_, _34382_);
  or (_34450_, _34449_, _34448_);
  or (_34451_, _34450_, _34196_);
  or (_34452_, _34451_, _34366_);
  or (_34453_, _34423_, _34435_);
  or (_34454_, _34427_, _34301_);
  or (_34455_, _34454_, _34453_);
  or (_34456_, _34122_, _30707_);
  or (_34457_, _34126_, _30803_);
  or (_34458_, _34457_, _34456_);
  not (_34459_, _30764_);
  or (_34460_, _30865_, _34459_);
  or (_34461_, _34460_, _34458_);
  or (_34462_, _34461_, _34455_);
  or (_34463_, _34462_, _34452_);
  and (_34464_, _34463_, _34008_);
  and (_34465_, _30490_, _35796_);
  and (_34466_, _34465_, _30726_);
  and (_34467_, _34102_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_34468_, _34467_, _34466_);
  or (_35996_[0], _34468_, _34464_);
  or (_34469_, _34320_, _30763_);
  or (_34470_, _34469_, _30760_);
  and (_34471_, _30706_, _30754_);
  or (_34472_, _34224_, _34151_);
  or (_34473_, _34472_, _34471_);
  or (_34474_, _34126_, _32134_);
  or (_34475_, _34474_, _30863_);
  or (_34476_, _34475_, _34473_);
  or (_34477_, _34476_, _34470_);
  or (_34478_, _34434_, _34371_);
  and (_34479_, _30807_, _30705_);
  or (_34480_, _34479_, _34319_);
  and (_34481_, _30853_, _30761_);
  or (_34482_, _34300_, _34481_);
  or (_34483_, _34482_, _34480_);
  or (_34484_, _34483_, _34478_);
  or (_34485_, _34484_, _34149_);
  or (_34486_, _34485_, _34143_);
  or (_34487_, _34486_, _34477_);
  and (_34488_, _34487_, _30494_);
  and (_34489_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34490_, _34489_, _30738_);
  or (_34491_, _34490_, _34488_);
  and (_35996_[1], _34491_, _35796_);
  or (_34492_, _34480_, _34469_);
  or (_34493_, _34492_, _34482_);
  or (_34494_, _30860_, _30855_);
  nor (_34495_, _34494_, _34426_);
  nand (_34496_, _34495_, _32137_);
  or (_34497_, _34436_, _34189_);
  or (_34498_, _34497_, _34496_);
  or (_34499_, _34148_, _34141_);
  or (_34500_, _34499_, _34498_);
  or (_34501_, _34500_, _34493_);
  and (_34502_, _34501_, _30494_);
  and (_34503_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34504_, _34503_, _30739_);
  or (_34505_, _34504_, _34502_);
  and (_35996_[2], _34505_, _35796_);
  and (_34506_, _34102_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_34507_, _34108_, _30827_);
  not (_34508_, _30704_);
  and (_34509_, _30807_, _34508_);
  or (_34510_, _34509_, _34421_);
  or (_34511_, _34510_, _34507_);
  not (_34512_, _32135_);
  or (_34513_, _34453_, _34512_);
  or (_34514_, _34513_, _34511_);
  or (_34515_, _34429_, _34223_);
  or (_34516_, _34515_, _34431_);
  or (_34517_, _34516_, _34514_);
  and (_34518_, _34517_, _34008_);
  or (_35997_[0], _34518_, _34506_);
  nor (_35983_[7], _30550_, rst);
  nor (_35984_[7], _32126_, rst);
  nor (_34519_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_34520_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_34521_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_34522_, _34521_, _34520_);
  and (_34523_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_34524_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_34525_, _34524_, _34523_);
  and (_34526_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_34527_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_34528_, _34527_, _34526_);
  and (_34529_, _34528_, _34525_);
  and (_34530_, _34529_, _34522_);
  and (_34531_, _34530_, _30632_);
  nor (_34532_, _34531_, _34519_);
  nor (_34533_, _34532_, _32110_);
  nor (_34534_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  nor (_34535_, _34534_, _34533_);
  and (_35985_[7], _34535_, _35796_);
  nor (_35983_[0], _30624_, rst);
  nor (_35983_[1], _30649_, rst);
  nor (_35983_[2], _30676_, rst);
  nor (_35983_[3], _30699_, rst);
  and (_35983_[4], _30527_, _35796_);
  nor (_35983_[5], _30597_, rst);
  nor (_35983_[6], _30574_, rst);
  nor (_35984_[0], _32245_, rst);
  nor (_35984_[1], _32458_, rst);
  nor (_35984_[2], _32349_, rst);
  nor (_35984_[3], _32197_, rst);
  nor (_35984_[4], _32400_, rst);
  nor (_35984_[5], _32297_, rst);
  nor (_35984_[6], _32514_, rst);
  nor (_34536_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_34537_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_34538_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_34539_, _34538_, _34537_);
  and (_34540_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_34541_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_34542_, _34541_, _34540_);
  and (_34543_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_34544_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_34545_, _34544_, _34543_);
  and (_34546_, _34545_, _34542_);
  and (_34547_, _34546_, _34539_);
  and (_34548_, _34547_, _30632_);
  nor (_34549_, _34548_, _34536_);
  nor (_34550_, _34549_, _32110_);
  nor (_34551_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  nor (_34552_, _34551_, _34550_);
  and (_35985_[0], _34552_, _35796_);
  nor (_34553_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_34554_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_34555_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_34556_, _34555_, _34554_);
  and (_34557_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_34558_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_34559_, _34558_, _34557_);
  and (_34560_, _34559_, _34556_);
  and (_34561_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_34562_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_34563_, _34562_, _34561_);
  and (_34564_, _34563_, _34560_);
  and (_34565_, _34564_, _30632_);
  nor (_34566_, _34565_, _34553_);
  nor (_34567_, _34566_, _32110_);
  nor (_34568_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  nor (_34569_, _34568_, _34567_);
  and (_35985_[1], _34569_, _35796_);
  nor (_34570_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_34571_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_34572_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_34573_, _34572_, _34571_);
  and (_34574_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_34575_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_34576_, _34575_, _34574_);
  and (_34577_, _34576_, _34573_);
  and (_34578_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_34579_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_34580_, _34579_, _34578_);
  and (_34581_, _34580_, _34577_);
  and (_34582_, _34581_, _30632_);
  nor (_34583_, _34582_, _34570_);
  nor (_34584_, _34583_, _32110_);
  nor (_34585_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  nor (_34586_, _34585_, _34584_);
  and (_35985_[2], _34586_, _35796_);
  nor (_34587_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_34588_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_34589_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_34590_, _34589_, _34588_);
  and (_34591_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_34592_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_34593_, _34592_, _34591_);
  and (_34594_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_34595_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_34596_, _34595_, _34594_);
  and (_34597_, _34596_, _34593_);
  and (_34598_, _34597_, _34590_);
  and (_34599_, _34598_, _30632_);
  nor (_34600_, _34599_, _34587_);
  nor (_34601_, _34600_, _32110_);
  nor (_34602_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  nor (_34603_, _34602_, _34601_);
  and (_35985_[3], _34603_, _35796_);
  nor (_34604_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_34605_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_34606_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_34607_, _34606_, _34605_);
  and (_34608_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_34609_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_34610_, _34609_, _34608_);
  and (_34611_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_34612_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_34613_, _34612_, _34611_);
  and (_34614_, _34613_, _34610_);
  and (_34615_, _34614_, _34607_);
  and (_34616_, _34615_, _30632_);
  nor (_34617_, _34616_, _34604_);
  nor (_34618_, _34617_, _32110_);
  nor (_34619_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  nor (_34620_, _34619_, _34618_);
  and (_35985_[4], _34620_, _35796_);
  nor (_34621_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_34622_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_34623_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34624_, _34623_, _34622_);
  and (_34625_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34626_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_34627_, _34626_, _34625_);
  and (_34628_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_34629_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_34630_, _34629_, _34628_);
  and (_34631_, _34630_, _34627_);
  and (_34632_, _34631_, _34624_);
  and (_34633_, _34632_, _30632_);
  nor (_34634_, _34633_, _34621_);
  nor (_34635_, _34634_, _32110_);
  nor (_34636_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  nor (_34637_, _34636_, _34635_);
  and (_35985_[5], _34637_, _35796_);
  nor (_34638_, _30632_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_34639_, _30516_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_34640_, _30504_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_34641_, _34640_, _34639_);
  and (_34642_, _30508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34643_, _30511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_34644_, _34643_, _34642_);
  and (_34645_, _30500_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_34646_, _30514_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_34647_, _34646_, _34645_);
  and (_34648_, _34647_, _34644_);
  and (_34649_, _34648_, _34641_);
  and (_34650_, _34649_, _30632_);
  nor (_34651_, _34650_, _34638_);
  nor (_34652_, _34651_, _32110_);
  nor (_34653_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  nor (_34654_, _34653_, _34652_);
  and (_35985_[6], _34654_, _35796_);
  and (_34655_, _30495_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_34656_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_34657_, _34655_, _31070_);
  and (_34658_, _34657_, _35796_);
  and (_36000_[15], _34658_, _34656_);
  not (_34659_, _34655_);
  or (_34660_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _34655_, _35796_);
  and (_34661_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _35796_);
  or (_34662_, _34661_, _00000_);
  and (_36001_[15], _34662_, _34660_);
  nor (_36002_, _32133_, rst);
  and (_36003_, \oc8051_top_1.oc8051_memory_interface1.dstb_o , _35796_);
  nor (_36004_[4], _32407_, rst);
  and (_36005_[7], _32105_, _35796_);
  nor (_34663_, _32133_, _28274_);
  and (_34664_, _32133_, _28274_);
  nor (_34665_, _34664_, _34663_);
  nor (_34666_, _32202_, _24213_);
  and (_34667_, _32202_, _24213_);
  nor (_34668_, _34667_, _34666_);
  and (_34669_, _34668_, _34665_);
  nor (_34670_, _32413_, _32078_);
  and (_34671_, _32413_, _32078_);
  nor (_34672_, _34671_, _34670_);
  nor (_34673_, _32521_, _30890_);
  and (_34674_, _32521_, _30890_);
  nor (_34675_, _34674_, _34673_);
  nor (_34676_, _32305_, _24532_);
  and (_34677_, _32305_, _24532_);
  nor (_34678_, _34677_, _34676_);
  and (_34679_, _34678_, _34675_);
  and (_34680_, _34679_, _34672_);
  and (_34681_, _34680_, _34669_);
  nor (_34682_, _32463_, _30163_);
  and (_34683_, _32463_, _30163_);
  or (_34684_, _34683_, _34682_);
  nor (_34685_, _34684_, _31713_);
  nor (_34686_, _32250_, _24653_);
  and (_34687_, _32250_, _24653_);
  nor (_34688_, _34687_, _34686_);
  nor (_34689_, _32354_, _24894_);
  and (_34690_, _32354_, _24894_);
  nor (_34691_, _34690_, _34689_);
  nor (_34692_, _34691_, _34688_);
  and (_34693_, _34692_, _34685_);
  and (_34694_, _34693_, _34681_);
  nor (_34695_, _23877_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_34696_, _34695_, _34694_);
  not (_34697_, _34696_);
  nor (_34698_, _30783_, _34131_);
  and (_34699_, _30476_, _27711_);
  and (_34700_, _34699_, _34698_);
  and (_34701_, _34700_, _34681_);
  nor (_34702_, _34106_, _34382_);
  nor (_34703_, _28461_, _26498_);
  and (_34704_, _34703_, _29707_);
  and (_34705_, _34704_, _30203_);
  and (_34706_, _34705_, _30347_);
  and (_34707_, _34706_, _30429_);
  not (_34708_, _30840_);
  and (_34709_, _32146_, _34708_);
  nor (_34710_, _34709_, _34131_);
  or (_34711_, _34710_, _30737_);
  nor (_34712_, _34711_, _30273_);
  and (_34713_, _34712_, _34707_);
  and (_34714_, _34713_, _26694_);
  nor (_34715_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_34716_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_34717_, _34716_, _34715_);
  nor (_34718_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_34719_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_34720_, _34719_, _34718_);
  and (_34721_, _34720_, _34717_);
  and (_34722_, _34721_, _30882_);
  not (_34723_, _30737_);
  nor (_34724_, _34698_, _30601_);
  nor (_34725_, _34724_, _34723_);
  and (_34726_, _34725_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_34727_, _34726_, _34722_);
  nor (_34728_, _34727_, _34714_);
  nand (_34729_, _34710_, _25686_);
  and (_34730_, _34729_, _34728_);
  not (_34731_, _34179_);
  nor (_34732_, _34370_, _30799_);
  and (_34733_, _34732_, _34731_);
  or (_34734_, _30716_, _30778_);
  nor (_34735_, _34734_, _30762_);
  nor (_34736_, _34735_, _30777_);
  nor (_34737_, _34736_, _34339_);
  and (_34738_, _34737_, _34733_);
  not (_34739_, _34738_);
  and (_34740_, _34739_, _34730_);
  and (_34741_, _30736_, _30532_);
  not (_34742_, _34741_);
  and (_34743_, _34742_, _30842_);
  nor (_34744_, _34743_, _34730_);
  nor (_34745_, _34744_, _34740_);
  and (_34746_, _34745_, _34702_);
  nor (_34747_, _34746_, _30843_);
  nor (_34748_, _34169_, _30490_);
  nor (_34749_, _34748_, _30879_);
  not (_34750_, _34749_);
  nor (_34751_, _34750_, _34747_);
  not (_34752_, _30882_);
  and (_34753_, _31503_, _31554_);
  nor (_34754_, _34753_, _34752_);
  nor (_34755_, _31386_, _31380_);
  and (_34756_, _34755_, _31446_);
  not (_34757_, _34756_);
  and (_34758_, _34757_, _34725_);
  nor (_34759_, _34758_, _34754_);
  not (_34760_, _34759_);
  nor (_34761_, _34760_, _34751_);
  not (_34762_, _34761_);
  nor (_34763_, _34762_, _34701_);
  and (_34764_, _34763_, _34697_);
  nor (_34765_, _30880_, rst);
  and (_36008_, _34765_, _34764_);
  and (_36009_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _35796_);
  nor (_34766_, \oc8051_top_1.oc8051_memory_interface1.dstb_o , rst);
  and (_34767_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_34768_, _36003_, xram_data_in_reg[7]);
  or (_36010_[7], _34768_, _34767_);
  nor (_34769_, _30507_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_34770_, _34769_, _32110_);
  nor (_34771_, _34770_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_34772_, _34771_);
  and (_34773_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_34774_, _34773_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_34775_, _34774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_34776_, _34775_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_34777_, _34776_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_34778_, _34777_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_34779_, _34778_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_34780_, _34779_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_34781_, _34780_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_34782_, _34781_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_34783_, _34782_, _34772_);
  and (_34784_, _34783_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_34785_, _34784_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_34786_, _34785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_34787_, _34694_, _28274_);
  and (_34788_, _34787_, _27668_);
  not (_34789_, _34788_);
  or (_34790_, _34747_, _30879_);
  nor (_34791_, _34790_, _34748_);
  and (_34792_, _30737_, _30601_);
  and (_34793_, _34757_, _34792_);
  or (_34794_, _34793_, _34791_);
  and (_34795_, _30715_, _30735_);
  nand (_34796_, _34795_, _30733_);
  nor (_34797_, _34753_, _34796_);
  and (_34798_, _34710_, _30476_);
  and (_34799_, _34798_, _27711_);
  and (_34800_, _34799_, _34681_);
  or (_34801_, _34800_, _34797_);
  nor (_34802_, _34801_, _34794_);
  and (_34803_, _34802_, _34789_);
  and (_34804_, _34785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_34805_, _34804_, _34803_);
  and (_34806_, _34805_, _34786_);
  and (_34807_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_34808_, _34807_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_34809_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_34810_, _34809_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_34811_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_34812_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34813_, _34812_, _34811_);
  and (_34814_, _34813_, _34810_);
  and (_34815_, _34814_, _34808_);
  and (_34816_, _34815_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_34817_, _34816_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34818_, _34817_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_34819_, _34818_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_34820_, _34819_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_34821_, _34819_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_34822_, _34821_, _34820_);
  nor (_34823_, _34339_, _30736_);
  and (_34824_, _34823_, _34702_);
  and (_34825_, _34733_, _30783_);
  and (_34826_, _34825_, _34824_);
  nor (_34827_, _34826_, _30843_);
  not (_34828_, _34827_);
  and (_34829_, _30735_, _34171_);
  and (_34830_, _34829_, _30754_);
  not (_34831_, _34830_);
  and (_34832_, _34732_, _34338_);
  and (_34833_, _34832_, _34709_);
  nor (_34834_, _34833_, _30843_);
  not (_34835_, _34834_);
  and (_34836_, _34168_, _34171_);
  nor (_34837_, _34836_, _30836_);
  and (_34838_, _34837_, _34835_);
  and (_34839_, _34838_, _34831_);
  and (_34840_, _34382_, _30733_);
  nor (_34841_, _34840_, _34748_);
  not (_34842_, _34841_);
  and (_34843_, _34842_, _34839_);
  and (_34844_, _34843_, _34828_);
  and (_34845_, _34844_, _34822_);
  nor (_34846_, _30837_, _27635_);
  not (_34847_, _34840_);
  nor (_34848_, _34847_, _31119_);
  and (_34849_, _34836_, _32127_);
  not (_34850_, _30880_);
  and (_34851_, _30775_, _34171_);
  nor (_34852_, _34851_, _34836_);
  and (_34853_, _34852_, _34850_);
  and (_34854_, _34853_, _34835_);
  nor (_34855_, _34827_, _34842_);
  and (_34856_, _34855_, _34854_);
  and (_34857_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_34858_, _34857_, _34849_);
  or (_34859_, _34858_, _34848_);
  or (_34860_, _34859_, _34846_);
  or (_34861_, _34860_, _34845_);
  and (_34862_, _34854_, _32126_);
  nor (_34863_, _34854_, _34535_);
  nor (_34864_, _34863_, _34862_);
  not (_34865_, _34864_);
  and (_34866_, _34864_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_34867_, _34864_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_34868_, _34854_, _32514_);
  nor (_34869_, _34854_, _34654_);
  nor (_34870_, _34869_, _34868_);
  and (_34871_, _34870_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_34872_, _34870_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_34873_, _34872_, _34871_);
  and (_34874_, _34854_, _32297_);
  nor (_34875_, _34854_, _34637_);
  nor (_34876_, _34875_, _34874_);
  and (_34877_, _34876_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_34878_, _34876_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_34879_, _34854_, _32400_);
  nor (_34880_, _34854_, _34620_);
  nor (_34881_, _34880_, _34879_);
  nand (_34882_, _34881_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34883_, _34854_, _32197_);
  nor (_34884_, _34854_, _34603_);
  nor (_34885_, _34884_, _34883_);
  and (_34886_, _34885_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_34887_, _34885_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_34888_, _34854_, _32349_);
  nor (_34889_, _34854_, _34586_);
  nor (_34890_, _34889_, _34888_);
  and (_34891_, _34890_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_34892_, _34854_, _32458_);
  nor (_34893_, _34854_, _34569_);
  nor (_34894_, _34893_, _34892_);
  and (_34895_, _34894_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_34896_, _34854_, _32245_);
  nor (_34897_, _34854_, _34552_);
  nor (_34898_, _34897_, _34896_);
  and (_34899_, _34898_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_34900_, _34894_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_34901_, _34900_, _34895_);
  and (_34902_, _34901_, _34899_);
  nor (_34903_, _34902_, _34895_);
  not (_34904_, _34903_);
  nor (_34905_, _34890_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_34906_, _34905_, _34891_);
  and (_34907_, _34906_, _34904_);
  nor (_34908_, _34907_, _34891_);
  nor (_34909_, _34908_, _34887_);
  or (_34910_, _34909_, _34886_);
  or (_34911_, _34881_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34912_, _34911_, _34882_);
  nand (_34913_, _34912_, _34910_);
  and (_34914_, _34913_, _34882_);
  nor (_34915_, _34914_, _34878_);
  or (_34916_, _34915_, _34877_);
  and (_34917_, _34916_, _34873_);
  nor (_34918_, _34917_, _34871_);
  nor (_34919_, _34918_, _34867_);
  or (_34920_, _34919_, _34866_);
  nor (_34921_, _34920_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_34922_, _34921_, _31048_);
  and (_34923_, _34922_, _31053_);
  and (_34924_, _34923_, _31038_);
  nor (_34925_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34926_, _34925_, _34924_);
  and (_34927_, _34926_, _31065_);
  nor (_34928_, _34927_, _34865_);
  and (_34929_, \oc8051_top_1.oc8051_memory_interface1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_34930_, _34929_, _34807_);
  and (_34931_, _34930_, _34920_);
  and (_34932_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34933_, _34932_, _34931_);
  and (_34934_, _34933_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_34935_, _34934_, _34864_);
  nor (_34936_, _34935_, _34928_);
  or (_34937_, _34936_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_34938_, _34936_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_34939_, _34938_, _34937_);
  nor (_34940_, _34827_, _34830_);
  nor (_34941_, _34940_, _34843_);
  and (_34942_, _34941_, _34939_);
  or (_34943_, _34942_, _34861_);
  and (_34944_, _34943_, _34803_);
  or (_34945_, _34944_, _34806_);
  and (_36011_[15], _34945_, _35796_);
  and (_34946_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _35796_);
  and (_34947_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_34948_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_34949_, _30494_, _34948_);
  not (_34950_, _34949_);
  not (_34951_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_34952_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_34953_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_34954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_34955_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_34956_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_34957_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_34958_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_34959_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_34960_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_34961_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_34962_, _34961_, _34960_);
  and (_34963_, _34962_, _34959_);
  and (_34964_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34965_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_34966_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_34967_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_34968_, _34967_, _34965_);
  and (_34969_, _34968_, _34966_);
  nor (_34970_, _34969_, _34965_);
  nor (_34971_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_34972_, _34971_, _34964_);
  not (_34973_, _34972_);
  nor (_34974_, _34973_, _34970_);
  nor (_34975_, _34974_, _34964_);
  and (_34976_, _34975_, _34963_);
  and (_34977_, _34976_, _34958_);
  and (_34978_, _34977_, _34957_);
  and (_34979_, _34978_, _34956_);
  and (_34980_, _34979_, _34955_);
  and (_34981_, _34980_, _34954_);
  and (_34982_, _34981_, _34953_);
  and (_34983_, _34982_, _34952_);
  and (_34984_, _34983_, _34951_);
  and (_34985_, _34984_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_34986_, _34984_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_34987_, _34986_, _34985_);
  nor (_34988_, _34983_, _34951_);
  or (_34989_, _34988_, _34984_);
  nor (_34990_, _34982_, _34952_);
  nor (_34991_, _34990_, _34983_);
  not (_34992_, _34991_);
  nor (_34993_, _34981_, _34953_);
  or (_34994_, _34993_, _34982_);
  nor (_34995_, _34980_, _34954_);
  nor (_34996_, _34995_, _34981_);
  not (_34997_, _34996_);
  nor (_34998_, _34979_, _34955_);
  nor (_34999_, _34998_, _34980_);
  not (_35000_, _34999_);
  nor (_35001_, _34978_, _34956_);
  or (_35002_, _35001_, _34979_);
  nor (_35003_, _34977_, _34957_);
  nor (_35004_, _35003_, _34978_);
  not (_35005_, _35004_);
  nor (_35006_, _34976_, _34958_);
  nor (_35007_, _35006_, _34977_);
  not (_35008_, _35007_);
  and (_35009_, _34975_, _34962_);
  nor (_35010_, _35009_, _34959_);
  nor (_35011_, _35010_, _34976_);
  not (_35012_, _35011_);
  and (_35013_, _34975_, _34961_);
  nor (_35014_, _35013_, _34960_);
  nor (_35015_, _35014_, _35009_);
  not (_35016_, _35015_);
  not (_35017_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_35018_, _34975_, _35017_);
  nor (_35019_, _34975_, _35017_);
  nor (_35020_, _35019_, _35018_);
  not (_35021_, _35020_);
  and (_35022_, _34082_, _34029_);
  nor (_35023_, _34083_, _34074_);
  and (_35024_, _34041_, _34029_);
  and (_35025_, _34050_, _34071_);
  and (_35026_, _35025_, _34068_);
  nor (_35027_, _35026_, _35024_);
  nand (_35028_, _35027_, _35023_);
  nor (_35029_, _35028_, _35022_);
  not (_35030_, _34082_);
  nor (_35031_, _34079_, _34065_);
  and (_35032_, _34028_, _34013_);
  not (_35033_, _35032_);
  and (_35034_, _34060_, _34013_);
  not (_35035_, _35034_);
  and (_35036_, _34018_, _34071_);
  nor (_35037_, _35036_, _34061_);
  and (_35038_, _35037_, _35035_);
  and (_35039_, _35038_, _35033_);
  and (_35040_, _35039_, _35031_);
  nor (_35041_, _35040_, _35030_);
  not (_35042_, _35041_);
  not (_35043_, _35025_);
  nor (_35044_, _34034_, _34027_);
  nor (_35045_, _35044_, _35043_);
  not (_35046_, _35045_);
  and (_35047_, _34075_, _34042_);
  not (_35048_, _34041_);
  nor (_35049_, _34079_, _34058_);
  nor (_35050_, _35049_, _35048_);
  nor (_35051_, _35050_, _35047_);
  and (_35052_, _35051_, _35046_);
  and (_35053_, _35052_, _35042_);
  and (_35054_, _35053_, _35029_);
  not (_35055_, _34034_);
  nor (_35056_, _34029_, _34014_);
  and (_35057_, _34072_, _34018_);
  nor (_35058_, _35057_, _34079_);
  and (_35059_, _35058_, _35056_);
  nor (_35060_, _35059_, _35055_);
  not (_35061_, _35060_);
  and (_35062_, _34049_, _34018_);
  not (_35063_, _35062_);
  and (_35064_, _35031_, _35063_);
  nor (_35065_, _35064_, _30699_);
  not (_35066_, _35065_);
  and (_35067_, _35066_, _34064_);
  and (_35068_, _35067_, _35061_);
  nor (_35069_, _34037_, _34025_);
  nor (_35070_, _34086_, _34066_);
  and (_35071_, _35070_, _35069_);
  and (_35072_, _34057_, _34018_);
  and (_35073_, _35072_, _30527_);
  not (_35074_, _35073_);
  nor (_35075_, _30649_, _30527_);
  and (_35076_, _35075_, _34018_);
  and (_35077_, _35076_, _34021_);
  not (_35078_, _35077_);
  and (_35079_, _34050_, _34016_);
  and (_35080_, _35079_, _34023_);
  nor (_35081_, _35080_, _34015_);
  and (_35082_, _35081_, _35078_);
  and (_35083_, _35082_, _35074_);
  and (_35084_, _35083_, _35071_);
  and (_35085_, _34049_, _34013_);
  and (_35086_, _35085_, _34082_);
  and (_35087_, _34065_, _34034_);
  nor (_35088_, _35087_, _35086_);
  nor (_35089_, _34033_, _34027_);
  not (_35090_, _35089_);
  and (_35091_, _34061_, _30624_);
  and (_35092_, _35091_, _35090_);
  not (_35093_, _34057_);
  nor (_35094_, _35062_, _34014_);
  nor (_35095_, _35094_, _35093_);
  nor (_35096_, _35095_, _35092_);
  and (_35097_, _35096_, _35088_);
  and (_35098_, _35090_, _34051_);
  and (_35099_, _35036_, _34041_);
  nor (_35100_, _35099_, _35098_);
  and (_35101_, _34068_, _34061_);
  and (_35102_, _34082_, _34035_);
  nor (_35103_, _35102_, _35101_);
  and (_35104_, _35103_, _35100_);
  and (_35105_, _35104_, _35097_);
  and (_35106_, _35105_, _35084_);
  and (_35107_, _35106_, _35068_);
  and (_35108_, _35107_, _35054_);
  not (_35109_, _35108_);
  nor (_35110_, _34968_, _34966_);
  nor (_35111_, _35110_, _34969_);
  nand (_35112_, _35111_, _35109_);
  and (_35113_, _35036_, _34057_);
  nor (_35114_, _35031_, _35030_);
  or (_35115_, _35114_, _35113_);
  and (_35116_, _34050_, _34011_);
  and (_35117_, _35116_, _34068_);
  nor (_35118_, _35117_, _34059_);
  nand (_35119_, _35118_, _35069_);
  nor (_35120_, _35119_, _35115_);
  nand (_35121_, _35120_, _35029_);
  or (_35122_, _35121_, _35108_);
  nor (_35123_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_35124_, _35123_, _34966_);
  and (_35125_, _35124_, _35122_);
  or (_35126_, _35111_, _35109_);
  and (_35127_, _35126_, _35112_);
  nand (_35128_, _35127_, _35125_);
  and (_35129_, _35128_, _35112_);
  not (_35130_, _35129_);
  and (_35131_, _34973_, _34970_);
  nor (_35132_, _35131_, _34974_);
  and (_35133_, _35132_, _35130_);
  and (_35134_, _35133_, _35021_);
  not (_35135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_35136_, _35018_, _35135_);
  or (_35137_, _35136_, _35013_);
  and (_35138_, _35137_, _35134_);
  and (_35139_, _35138_, _35016_);
  and (_35140_, _35139_, _35012_);
  and (_35141_, _35140_, _35008_);
  and (_35142_, _35141_, _35005_);
  and (_35143_, _35142_, _35002_);
  and (_35144_, _35143_, _35000_);
  and (_35145_, _35144_, _34997_);
  and (_35146_, _35145_, _34994_);
  and (_35147_, _35146_, _34992_);
  and (_35148_, _35147_, _34989_);
  and (_35149_, _35148_, _34987_);
  nor (_35150_, _35148_, _34987_);
  or (_35151_, _35150_, _35149_);
  or (_35152_, _35151_, _34950_);
  or (_35153_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_35154_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_35155_, _35154_, _35153_);
  and (_35156_, _35155_, _35152_);
  or (_36012_[15], _35156_, _34947_);
  nor (_35157_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_36013_, _35157_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_36014_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _35796_);
  and (_35158_, \oc8051_top_1.oc8051_rom1.ea_int , _30491_);
  nand (_35159_, _35158_, _30494_);
  and (_36015_, _35159_, _36014_);
  and (_36016_[7], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _35796_);
  nor (_35160_, _34771_, _32110_);
  or (_35161_, _35108_, _30502_);
  and (_35162_, _35122_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_35163_, _35108_, _30502_);
  and (_35164_, _35163_, _35161_);
  nand (_35165_, _35164_, _35162_);
  and (_35166_, _35165_, _35161_);
  nor (_35167_, _35166_, _32110_);
  and (_35168_, _35167_, _30498_);
  nor (_35169_, _35167_, _30498_);
  nor (_35170_, _35169_, _35168_);
  nor (_35171_, _35170_, _35160_);
  and (_35172_, _30503_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_35173_, _35172_, _35160_);
  and (_35174_, _35173_, _35121_);
  or (_35175_, _35174_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_35176_, _35175_, _35171_);
  and (_36017_[2], _35176_, _35796_);
  nor (_35177_, _30618_, _30568_);
  not (_35178_, _30546_);
  and (_35179_, _30591_, _35178_);
  and (_35180_, _35179_, _35177_);
  not (_35181_, _30520_);
  and (_35182_, _30495_, _35796_);
  and (_35183_, _35182_, _30669_);
  and (_35184_, _35183_, _35181_);
  nor (_35185_, _30693_, _30644_);
  and (_35186_, _35185_, _35184_);
  and (_36020_, _35186_, _35180_);
  nor (_35187_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_35188_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_35189_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_36022_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _35796_);
  and (_35190_, _36022_, _35189_);
  or (_36021_[7], _35190_, _35188_);
  not (_35191_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_35192_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_35193_, _35192_, _35191_);
  and (_35194_, _35192_, _35191_);
  nor (_35195_, _35194_, _35193_);
  not (_35196_, _35195_);
  and (_35197_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_35198_, _35197_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_35199_, _35197_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_35200_, _35199_, _35198_);
  or (_35201_, _35200_, _35192_);
  and (_35202_, _35201_, _35196_);
  nor (_35203_, _35193_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_35204_, _35193_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_35205_, _35204_, _35203_);
  or (_35206_, _35198_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_36024_[3], _35206_, _35796_);
  and (_35207_, _36024_[3], _35205_);
  and (_36023_, _35207_, _35202_);
  not (_35208_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_35209_, _34771_, _35208_);
  and (_35210_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_35211_, _35209_);
  and (_35212_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_35213_, _35212_, _35210_);
  and (_36025_[31], _35213_, _35796_);
  and (_35214_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_35215_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_35216_, _35215_, _35214_);
  and (_36026_[31], _35216_, _35796_);
  not (_35217_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  nor (_35218_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  nor (_35219_, _35218_, _35217_);
  and (_35220_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_35221_, _35220_, _35218_);
  or (_35222_, _35221_, _35219_);
  and (_36027_[7], _35222_, _35796_);
  not (_35223_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_35224_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _35223_);
  and (_35225_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_35226_, _35225_, _35224_);
  and (_36028_, _35226_, _34766_);
  and (_36029_, _35218_, _35796_);
  not (_35227_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  nor (_35228_, _35218_, _35227_);
  not (_35229_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_35230_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_35231_, _35230_, _35218_);
  or (_35232_, _35231_, _35228_);
  and (_36030_[15], _35232_, _35796_);
  or (_35233_, _35223_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_36031_, _35233_, _34766_);
  nor (_35234_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_35235_, _35234_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_35236_, _35235_, _35796_);
  and (_35237_, _36022_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_36032_, _35237_, _35236_);
  and (_35238_, _35208_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_35239_, _35238_, _35235_);
  and (_36033_, _35239_, _35796_);
  nand (_35240_, _35235_, _31119_);
  or (_35241_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_35242_, _35241_, _35796_);
  and (_36034_[15], _35242_, _35240_);
  nand (_35243_, _30745_, _35796_);
  nor (_36035_, _35243_, _30886_);
  or (_35244_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_35245_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_35246_, _34655_, _35245_);
  and (_35247_, _35246_, _35796_);
  and (_36000_[0], _35247_, _35244_);
  or (_35248_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_35249_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_35250_, _34655_, _35249_);
  and (_35251_, _35250_, _35796_);
  and (_36000_[1], _35251_, _35248_);
  or (_35252_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_35253_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], _35796_);
  or (_35254_, _35253_, _00000_);
  and (_36000_[2], _35254_, _35252_);
  or (_35255_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_35256_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_35257_, _34655_, _35256_);
  and (_35258_, _35257_, _35796_);
  and (_36000_[3], _35258_, _35255_);
  or (_35259_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_35260_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_35261_, _34655_, _35260_);
  and (_35262_, _35261_, _35796_);
  and (_36000_[4], _35262_, _35259_);
  or (_35263_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_35264_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_35265_, _34655_, _35264_);
  and (_35266_, _35265_, _35796_);
  and (_36000_[5], _35266_, _35263_);
  or (_35267_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_35268_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_35269_, _34655_, _35268_);
  and (_35270_, _35269_, _35796_);
  and (_36000_[6], _35270_, _35267_);
  or (_35271_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_35272_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_35273_, _34655_, _35272_);
  and (_35274_, _35273_, _35796_);
  and (_36000_[7], _35274_, _35271_);
  or (_35275_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_35276_, _34655_, _31042_);
  and (_35277_, _35276_, _35796_);
  and (_36000_[8], _35277_, _35275_);
  or (_35278_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_35279_, _34655_, _31048_);
  and (_35280_, _35279_, _35796_);
  and (_36000_[9], _35280_, _35278_);
  or (_35281_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_35282_, _34655_, _31053_);
  and (_35283_, _35282_, _35796_);
  and (_36000_[10], _35283_, _35281_);
  or (_35284_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_35285_, _34655_, _31038_);
  and (_35286_, _35285_, _35796_);
  and (_36000_[11], _35286_, _35284_);
  or (_35287_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_35288_, _34655_, _31059_);
  and (_35289_, _35288_, _35796_);
  and (_36000_[12], _35289_, _35287_);
  or (_35290_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_35291_, _34655_, _31034_);
  and (_35292_, _35291_, _35796_);
  and (_36000_[13], _35292_, _35290_);
  or (_35293_, _34655_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_35294_, _34655_, _31065_);
  and (_35295_, _35294_, _35796_);
  and (_36000_[14], _35295_, _35293_);
  or (_35296_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_35297_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _35796_);
  or (_35298_, _35297_, _00000_);
  and (_36001_[0], _35298_, _35296_);
  or (_35299_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_35300_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _35796_);
  or (_35301_, _35300_, _00000_);
  and (_36001_[1], _35301_, _35299_);
  or (_35302_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_35303_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _35796_);
  or (_35304_, _35303_, _00000_);
  and (_36001_[2], _35304_, _35302_);
  or (_35305_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_35306_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _35796_);
  or (_35307_, _35306_, _00000_);
  and (_36001_[3], _35307_, _35305_);
  or (_35308_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_35309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _35796_);
  or (_35310_, _35309_, _00000_);
  and (_36001_[4], _35310_, _35308_);
  or (_35311_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_35312_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _35796_);
  or (_35313_, _35312_, _00000_);
  and (_36001_[5], _35313_, _35311_);
  or (_35314_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_35315_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _35796_);
  or (_35316_, _35315_, _00000_);
  and (_36001_[6], _35316_, _35314_);
  or (_35317_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_35318_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _35796_);
  or (_35319_, _35318_, _00000_);
  and (_36001_[7], _35319_, _35317_);
  or (_35320_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_35321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _35796_);
  or (_35322_, _35321_, _00000_);
  and (_36001_[8], _35322_, _35320_);
  or (_35323_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_35324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _35796_);
  or (_35325_, _35324_, _00000_);
  and (_36001_[9], _35325_, _35323_);
  or (_35326_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_35327_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _35796_);
  or (_35328_, _35327_, _00000_);
  and (_36001_[10], _35328_, _35326_);
  or (_35329_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_35330_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _35796_);
  or (_35331_, _35330_, _00000_);
  and (_36001_[11], _35331_, _35329_);
  or (_35332_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_35333_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _35796_);
  or (_35334_, _35333_, _00000_);
  and (_36001_[12], _35334_, _35332_);
  or (_35335_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_35336_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _35796_);
  or (_35337_, _35336_, _00000_);
  and (_36001_[13], _35337_, _35335_);
  or (_35338_, _34659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_35339_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _35796_);
  or (_35340_, _35339_, _00000_);
  and (_36001_[14], _35340_, _35338_);
  and (_35341_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_35342_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_35343_, _35342_, _35341_);
  and (_36025_[0], _35343_, _35796_);
  and (_35344_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_35345_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_35346_, _35345_, _35344_);
  and (_36025_[1], _35346_, _35796_);
  and (_35347_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_35348_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_35349_, _35348_, _35347_);
  and (_36025_[2], _35349_, _35796_);
  and (_35350_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_35351_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_35352_, _35351_, _35350_);
  and (_36025_[3], _35352_, _35796_);
  and (_35353_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_35354_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_35355_, _35354_, _35209_);
  or (_35356_, _35355_, _35353_);
  and (_36025_[4], _35356_, _35796_);
  and (_35357_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_35358_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_35359_, _35358_, _35209_);
  or (_35360_, _35359_, _35357_);
  and (_36025_[5], _35360_, _35796_);
  and (_35361_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_35362_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_35363_, _35362_, _35361_);
  and (_36025_[6], _35363_, _35796_);
  and (_35364_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_35365_, _35209_, _35189_);
  or (_35366_, _35365_, _35364_);
  and (_36025_[7], _35366_, _35796_);
  and (_35367_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_35368_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_35369_, _35368_, _35367_);
  and (_36025_[8], _35369_, _35796_);
  and (_35370_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_35371_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_35372_, _35371_, _35370_);
  and (_36025_[9], _35372_, _35796_);
  and (_35373_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_35374_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_35375_, _35374_, _35373_);
  and (_36025_[10], _35375_, _35796_);
  and (_35376_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_35377_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_35378_, _35377_, _35376_);
  and (_36025_[11], _35378_, _35796_);
  and (_35379_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_35380_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_35381_, _35380_, _35379_);
  and (_36025_[12], _35381_, _35796_);
  and (_35382_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_35383_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_35384_, _35383_, _35382_);
  and (_36025_[13], _35384_, _35796_);
  and (_35385_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_35386_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_35387_, _35386_, _35385_);
  and (_36025_[14], _35387_, _35796_);
  and (_35388_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_35389_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_35390_, _35389_, _35388_);
  and (_36025_[15], _35390_, _35796_);
  and (_35391_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_35392_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_35393_, _35392_, _35391_);
  and (_36025_[16], _35393_, _35796_);
  and (_35394_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_35395_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_35396_, _35395_, _35394_);
  and (_36025_[17], _35396_, _35796_);
  and (_35397_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_35398_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_35399_, _35398_, _35397_);
  and (_36025_[18], _35399_, _35796_);
  and (_35400_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_35401_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_35402_, _35401_, _35400_);
  and (_36025_[19], _35402_, _35796_);
  and (_35403_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_35404_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_35405_, _35404_, _35403_);
  and (_36025_[20], _35405_, _35796_);
  and (_35406_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_35407_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_35408_, _35407_, _35406_);
  and (_36025_[21], _35408_, _35796_);
  and (_35409_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_35410_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_35411_, _35410_, _35409_);
  and (_36025_[22], _35411_, _35796_);
  and (_35412_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_35413_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_35414_, _35413_, _35412_);
  and (_36025_[23], _35414_, _35796_);
  and (_35415_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_35416_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_35417_, _35416_, _35415_);
  and (_36025_[24], _35417_, _35796_);
  and (_35418_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_35419_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_35420_, _35419_, _35418_);
  and (_36025_[25], _35420_, _35796_);
  and (_35421_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_35422_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_35423_, _35422_, _35421_);
  and (_36025_[26], _35423_, _35796_);
  and (_35424_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_35425_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_35426_, _35425_, _35424_);
  and (_36025_[27], _35426_, _35796_);
  and (_35427_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_35428_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_35429_, _35428_, _35427_);
  and (_36025_[28], _35429_, _35796_);
  and (_35430_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_35431_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_35432_, _35431_, _35430_);
  and (_36025_[29], _35432_, _35796_);
  and (_35433_, _35209_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_35434_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_35435_, _35434_, _35433_);
  and (_36025_[30], _35435_, _35796_);
  nor (_36004_[0], _30628_, rst);
  nor (_36004_[1], _30655_, rst);
  nor (_36004_[2], _30680_, rst);
  nor (_36004_[3], _32048_, rst);
  and (_36005_[0], _32225_, _35796_);
  and (_36005_[1], _32443_, _35796_);
  and (_36005_[2], _32329_, _35796_);
  and (_36005_[3], _32173_, _35796_);
  and (_36005_[4], _32382_, _35796_);
  nor (_36005_[5], _32279_, rst);
  nor (_36005_[6], _32497_, rst);
  and (_35436_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0]);
  and (_35437_, _36003_, xram_data_in_reg[0]);
  or (_36010_[0], _35437_, _35436_);
  and (_35438_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1]);
  and (_35439_, _36003_, xram_data_in_reg[1]);
  or (_36010_[1], _35439_, _35438_);
  and (_35440_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2]);
  and (_35441_, _36003_, xram_data_in_reg[2]);
  or (_36010_[2], _35441_, _35440_);
  and (_35442_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3]);
  and (_35443_, _36003_, xram_data_in_reg[3]);
  or (_36010_[3], _35443_, _35442_);
  and (_35444_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4]);
  and (_35445_, _36003_, xram_data_in_reg[4]);
  or (_36010_[4], _35445_, _35444_);
  and (_35446_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5]);
  and (_35447_, _36003_, xram_data_in_reg[5]);
  or (_36010_[5], _35447_, _35446_);
  and (_35448_, _34766_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6]);
  and (_35449_, _36003_, xram_data_in_reg[6]);
  or (_36010_[6], _35449_, _35448_);
  or (_35450_, _34764_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_35451_, _35450_, _35796_);
  or (_35452_, _34856_, _34840_);
  and (_35453_, _35452_, _28750_);
  or (_35454_, _34898_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_35455_, _34899_);
  and (_35456_, _34842_, _34854_);
  nor (_35457_, _34827_, _34851_);
  nor (_35458_, _35457_, _35456_);
  and (_35459_, _35458_, _35455_);
  and (_35460_, _35459_, _35454_);
  and (_35461_, _34828_, _35456_);
  and (_35462_, _35461_, _32246_);
  and (_35463_, _34836_, _34552_);
  and (_35464_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_35465_, _35464_, _35463_);
  or (_35466_, _35465_, _35462_);
  nor (_35467_, _35466_, _35460_);
  nand (_35468_, _35467_, _34764_);
  or (_35469_, _35468_, _35453_);
  and (_36011_[0], _35469_, _35451_);
  or (_35470_, _34764_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_35471_, _35470_, _35796_);
  and (_35472_, _35452_, _29390_);
  or (_35473_, _34901_, _34899_);
  not (_35474_, _34902_);
  and (_35475_, _35458_, _35474_);
  and (_35476_, _35475_, _35473_);
  and (_35477_, _34836_, _34569_);
  and (_35478_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_35479_, _35461_, _32459_);
  or (_35480_, _35479_, _35478_);
  or (_35481_, _35480_, _35477_);
  nor (_35482_, _35481_, _35476_);
  nand (_35483_, _35482_, _34764_);
  or (_35484_, _35483_, _35472_);
  and (_36011_[1], _35484_, _35471_);
  not (_35485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_35486_, _34771_, _35485_);
  and (_35487_, _34771_, _35485_);
  nor (_35488_, _35487_, _35486_);
  or (_35489_, _35488_, _34764_);
  and (_35490_, _35489_, _35796_);
  and (_35491_, _35452_, _30035_);
  or (_35492_, _34906_, _34904_);
  not (_35493_, _34907_);
  and (_35494_, _35458_, _35493_);
  and (_35495_, _35494_, _35492_);
  and (_35496_, _34836_, _34586_);
  and (_35497_, _35461_, _32350_);
  and (_35498_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_35499_, _35498_, _35497_);
  or (_35500_, _35499_, _35496_);
  nor (_35501_, _35500_, _35495_);
  nand (_35502_, _35501_, _34764_);
  or (_35503_, _35502_, _35491_);
  and (_36011_[2], _35503_, _35490_);
  and (_35504_, _35486_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_35505_, _35486_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_35506_, _35505_, _35504_);
  or (_35507_, _35506_, _34764_);
  and (_35508_, _35507_, _35796_);
  and (_35509_, _35452_, _30248_);
  or (_35510_, _34887_, _34886_);
  nand (_35511_, _35510_, _34908_);
  or (_35512_, _35510_, _34908_);
  and (_35513_, _35512_, _35458_);
  and (_35514_, _35513_, _35511_);
  and (_35515_, _34836_, _34603_);
  and (_35516_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_35517_, _35461_, _32198_);
  or (_35518_, _35517_, _35516_);
  or (_35519_, _35518_, _35515_);
  nor (_35520_, _35519_, _35514_);
  nand (_35521_, _35520_, _34764_);
  or (_35522_, _35521_, _35509_);
  and (_36011_[3], _35522_, _35508_);
  and (_35523_, _34774_, _34772_);
  nor (_35524_, _35504_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_35525_, _35524_, _35523_);
  or (_35526_, _35525_, _34764_);
  and (_35527_, _35526_, _35796_);
  and (_35528_, _35452_, _30320_);
  or (_35529_, _34912_, _34910_);
  and (_35530_, _35458_, _34913_);
  and (_35531_, _35530_, _35529_);
  and (_35532_, _34836_, _34620_);
  and (_35533_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_35534_, _35461_, _32401_);
  or (_35535_, _35534_, _35533_);
  or (_35536_, _35535_, _35532_);
  nor (_35537_, _35536_, _35531_);
  nand (_35538_, _35537_, _34764_);
  or (_35539_, _35538_, _35528_);
  and (_36011_[4], _35539_, _35527_);
  not (_35540_, _34775_);
  nor (_35541_, _35540_, _34771_);
  nor (_35542_, _35523_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_35543_, _35542_, _35541_);
  or (_35544_, _35543_, _34764_);
  and (_35545_, _35544_, _35796_);
  and (_35546_, _35452_, _30397_);
  or (_35547_, _34878_, _34877_);
  or (_35548_, _35547_, _34914_);
  nand (_35549_, _35547_, _34914_);
  and (_35550_, _35549_, _35458_);
  and (_35551_, _35550_, _35548_);
  and (_35552_, _35461_, _32298_);
  and (_35553_, _34836_, _34637_);
  and (_35554_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_35555_, _35554_, _35553_);
  or (_35556_, _35555_, _35552_);
  nor (_35557_, _35556_, _35551_);
  nand (_35558_, _35557_, _34764_);
  or (_35559_, _35558_, _35546_);
  and (_36011_[5], _35559_, _35545_);
  nor (_35560_, _35541_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35561_, _35541_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_35562_, _35561_, _35560_);
  or (_35563_, _35562_, _34764_);
  and (_35564_, _35563_, _35796_);
  and (_35565_, _35452_, _30469_);
  or (_35566_, _34916_, _34873_);
  not (_35567_, _34917_);
  and (_35568_, _35458_, _35567_);
  nand (_35569_, _35568_, _35566_);
  and (_35570_, _34836_, _34654_);
  and (_35571_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35572_, _35461_, _32515_);
  or (_35573_, _35572_, _35571_);
  nor (_35574_, _35573_, _35570_);
  and (_35575_, _35574_, _35569_);
  nand (_35576_, _35575_, _34764_);
  or (_35577_, _35576_, _35565_);
  and (_36011_[6], _35577_, _35564_);
  nor (_35578_, _35561_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_35579_, _35561_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_35580_, _35579_, _35578_);
  or (_35581_, _35580_, _34764_);
  and (_35582_, _35581_, _35796_);
  and (_35583_, _35452_, _27646_);
  or (_35584_, _34866_, _34867_);
  or (_35585_, _35584_, _34918_);
  nand (_35586_, _35584_, _34918_);
  and (_35587_, _35586_, _35458_);
  and (_35588_, _35587_, _35585_);
  and (_35589_, _34836_, _34535_);
  and (_35590_, _30880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_35591_, _35461_, _32127_);
  or (_35592_, _35591_, _35590_);
  nor (_35593_, _35592_, _35589_);
  nand (_35594_, _35593_, _34764_);
  or (_35595_, _35594_, _35588_);
  or (_35596_, _35595_, _35583_);
  and (_36011_[7], _35596_, _35582_);
  not (_35597_, _34803_);
  nor (_35598_, _34847_, _31157_);
  and (_35599_, _34920_, _31042_);
  nor (_35600_, _34920_, _31042_);
  nor (_35601_, _35600_, _35599_);
  or (_35602_, _35601_, _34865_);
  nand (_35603_, _35601_, _34865_);
  and (_35604_, _35603_, _35458_);
  and (_35605_, _35604_, _35602_);
  and (_35606_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_35607_, _34836_, _32246_);
  or (_35608_, _35607_, _35606_);
  and (_35609_, _35461_, _34016_);
  or (_35610_, _35609_, _35608_);
  or (_35611_, _35610_, _35605_);
  or (_35612_, _35611_, _35598_);
  nor (_35613_, _30837_, _28739_);
  or (_35614_, _35613_, _35612_);
  or (_35615_, _35614_, _35597_);
  or (_35616_, _35579_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_35617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35618_, _35617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_35619_, _35618_, _35541_);
  and (_35620_, _35619_, _35616_);
  or (_35621_, _35620_, _34803_);
  and (_35622_, _35621_, _35796_);
  and (_36011_[8], _35622_, _35615_);
  nor (_35623_, _30837_, _29380_);
  nor (_35624_, _34847_, _31189_);
  and (_35625_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_35626_, _34836_, _32459_);
  and (_35627_, _35461_, _34017_);
  or (_35628_, _35627_, _35626_);
  or (_35629_, _35628_, _35625_);
  or (_35630_, _35629_, _35624_);
  and (_35631_, _34920_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_35632_, _35631_, _34865_);
  and (_35633_, _34921_, _34864_);
  nor (_35634_, _35633_, _35632_);
  and (_35635_, _35634_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_35636_, _35634_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_35637_, _35636_, _35635_);
  and (_35638_, _35637_, _35458_);
  or (_35639_, _35638_, _35630_);
  or (_35640_, _35639_, _35597_);
  or (_35641_, _35640_, _35623_);
  nand (_35642_, _35619_, _34956_);
  or (_35643_, _35619_, _34956_);
  and (_35644_, _35643_, _35642_);
  or (_35645_, _35644_, _34803_);
  and (_35646_, _35645_, _35796_);
  and (_36011_[9], _35646_, _35641_);
  and (_35647_, _35618_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_35648_, _35647_, _35541_);
  and (_35649_, _35648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_35650_, _35648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_35651_, _35650_, _35649_);
  or (_35652_, _35651_, _34764_);
  and (_35653_, _35652_, _35796_);
  nor (_35654_, _30837_, _30024_);
  nor (_35655_, _34847_, _31219_);
  and (_35656_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_35657_, _34836_, _32350_);
  not (_35658_, _30550_);
  and (_35659_, _35461_, _35658_);
  or (_35660_, _35659_, _35657_);
  or (_35661_, _35660_, _35656_);
  or (_35662_, _35661_, _35655_);
  and (_35663_, _34922_, _34864_);
  and (_35664_, _35632_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_35665_, _35664_, _35663_);
  nand (_35666_, _35665_, _31053_);
  or (_35667_, _35665_, _31053_);
  and (_35668_, _35667_, _35666_);
  and (_35669_, _35668_, _34941_);
  or (_35670_, _35669_, _35662_);
  or (_35671_, _35670_, _35654_);
  or (_35672_, _35671_, _35597_);
  and (_36011_[10], _35672_, _35653_);
  nor (_35673_, _35649_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_35674_, _34779_, _34772_);
  and (_35675_, _35674_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_35676_, _35675_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_35677_, _35676_, _35673_);
  or (_35678_, _35677_, _34764_);
  and (_35679_, _35678_, _35796_);
  nor (_35680_, _30837_, _30247_);
  nor (_35681_, _34847_, _31250_);
  and (_35682_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_35683_, _34836_, _32198_);
  and (_35684_, _34814_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_35685_, _35684_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_35686_, _35685_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_35687_, _35686_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_35688_, _35686_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_35689_, _35688_, _35687_);
  and (_35690_, _35689_, _35461_);
  or (_35691_, _35690_, _35683_);
  or (_35692_, _35691_, _35682_);
  or (_35693_, _35692_, _35681_);
  and (_35694_, _34808_, _34920_);
  and (_35695_, _35694_, _34865_);
  and (_35696_, _34923_, _34864_);
  nor (_35697_, _35696_, _35695_);
  nor (_35698_, _35697_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_35699_, _35697_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_35700_, _35699_, _35698_);
  and (_35701_, _35700_, _34941_);
  or (_35702_, _35701_, _35693_);
  or (_35703_, _35702_, _35680_);
  or (_35704_, _35703_, _35597_);
  and (_36011_[11], _35704_, _35679_);
  and (_35705_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_35706_, _35705_, _35649_);
  nor (_35707_, _35676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_35708_, _35707_, _35706_);
  or (_35709_, _35708_, _34764_);
  and (_35710_, _35709_, _35796_);
  nor (_35711_, _34850_, _30319_);
  and (_35712_, _34931_, _34865_);
  and (_35713_, _34924_, _34864_);
  nor (_35714_, _35713_, _35712_);
  nand (_35715_, _35714_, _31059_);
  or (_35716_, _35714_, _31059_);
  and (_35717_, _35716_, _35458_);
  and (_35718_, _35717_, _35715_);
  nor (_35719_, _34847_, _31281_);
  and (_35720_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_35721_, _34836_, _32401_);
  or (_35722_, _35721_, _35720_);
  nor (_35723_, _34816_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_35724_, _35723_, _34817_);
  and (_35725_, _35724_, _35461_);
  or (_35726_, _35725_, _35722_);
  nor (_35727_, _35726_, _35719_);
  nand (_35728_, _35727_, _34764_);
  or (_35729_, _35728_, _35718_);
  or (_35730_, _35729_, _35711_);
  and (_36011_[12], _35730_, _35710_);
  and (_35731_, _35706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_35732_, _35706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_35733_, _35732_, _35731_);
  or (_35734_, _35733_, _34764_);
  and (_35735_, _35734_, _35796_);
  nor (_35736_, _34850_, _30396_);
  nand (_35737_, _35712_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_35738_, _35713_, _31059_);
  and (_35739_, _35738_, _35737_);
  nand (_35740_, _35739_, _31034_);
  or (_35741_, _35739_, _31034_);
  and (_35742_, _35741_, _35458_);
  and (_35743_, _35742_, _35740_);
  nor (_35744_, _34847_, _31315_);
  and (_35745_, _34836_, _32298_);
  and (_35746_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_35747_, _34817_, _31034_);
  and (_35748_, _34817_, _31034_);
  or (_35749_, _35748_, _35747_);
  and (_35750_, _35749_, _35461_);
  or (_35751_, _35750_, _35746_);
  or (_35752_, _35751_, _35745_);
  nor (_35753_, _35752_, _35744_);
  nand (_35754_, _35753_, _34764_);
  or (_35755_, _35754_, _35743_);
  or (_35756_, _35755_, _35736_);
  and (_36011_[13], _35756_, _35735_);
  nor (_35757_, _35731_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_35758_, _35757_, _34785_);
  or (_35759_, _35758_, _34764_);
  and (_35760_, _35759_, _35796_);
  nor (_35761_, _34933_, _34864_);
  nor (_35762_, _34926_, _34865_);
  nor (_35763_, _35762_, _35761_);
  nand (_35764_, _35763_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_35765_, _35763_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_35766_, _35765_, _34941_);
  and (_35767_, _35766_, _35764_);
  nor (_35768_, _34818_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_35769_, _35768_, _34819_);
  and (_35770_, _35769_, _34844_);
  nor (_35771_, _30837_, _30468_);
  nor (_35772_, _34847_, _31344_);
  and (_35773_, _34836_, _32515_);
  and (_35774_, _34856_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_35775_, _35774_, _35773_);
  or (_35776_, _35775_, _35772_);
  or (_35777_, _35776_, _35771_);
  or (_35778_, _35777_, _35770_);
  or (_35779_, _35778_, _35767_);
  or (_35780_, _35779_, _35597_);
  and (_36011_[14], _35780_, _35760_);
  and (_35781_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_35782_, _35124_, _35122_);
  nor (_35783_, _35782_, _35125_);
  or (_35784_, _35783_, _34950_);
  or (_35785_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35786_, _35785_, _35154_);
  and (_35787_, _35786_, _35784_);
  or (_36012_[0], _35787_, _35781_);
  or (_35788_, _35127_, _35125_);
  and (_35789_, _35788_, _35128_);
  or (_35790_, _35789_, _34950_);
  or (_35791_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_35792_, _35791_, _35154_);
  and (_35793_, _35792_, _35790_);
  and (_35794_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_36012_[1], _35794_, _35793_);
  and (_00009_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00010_, _35132_, _35130_);
  nor (_00011_, _00010_, _35133_);
  or (_00012_, _00011_, _34950_);
  or (_00013_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00014_, _00013_, _35154_);
  and (_00015_, _00014_, _00012_);
  or (_36012_[2], _00015_, _00009_);
  and (_00016_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00017_, _35133_, _35021_);
  nor (_00018_, _00017_, _35134_);
  or (_00019_, _00018_, _34950_);
  or (_00020_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00021_, _00020_, _35154_);
  and (_00022_, _00021_, _00019_);
  or (_36012_[3], _00022_, _00016_);
  nor (_00023_, _35137_, _35134_);
  nor (_00024_, _00023_, _35138_);
  or (_00025_, _00024_, _34950_);
  or (_00026_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00027_, _00026_, _35154_);
  and (_00028_, _00027_, _00025_);
  and (_00029_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_36012_[4], _00029_, _00028_);
  nor (_00030_, _35138_, _35016_);
  nor (_00031_, _00030_, _35139_);
  or (_00032_, _00031_, _34950_);
  or (_00033_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00034_, _00033_, _35154_);
  and (_00035_, _00034_, _00032_);
  and (_00036_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_36012_[5], _00036_, _00035_);
  and (_00037_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00038_, _35139_, _35012_);
  nor (_00039_, _00038_, _35140_);
  or (_00040_, _00039_, _34950_);
  or (_00041_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00042_, _00041_, _35154_);
  and (_00043_, _00042_, _00040_);
  or (_36012_[6], _00043_, _00037_);
  nor (_00044_, _35140_, _35008_);
  nor (_00045_, _00044_, _35141_);
  or (_00046_, _00045_, _34950_);
  or (_00047_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00048_, _00047_, _35154_);
  and (_00049_, _00048_, _00046_);
  and (_00050_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_36012_[7], _00050_, _00049_);
  nor (_00051_, _35141_, _35005_);
  nor (_00052_, _00051_, _35142_);
  or (_00053_, _00052_, _34950_);
  or (_00054_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00055_, _00054_, _35154_);
  and (_00056_, _00055_, _00053_);
  and (_00057_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_36012_[8], _00057_, _00056_);
  nor (_00058_, _35142_, _35002_);
  nor (_00059_, _00058_, _35143_);
  or (_00060_, _00059_, _34950_);
  or (_00061_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00062_, _00061_, _35154_);
  and (_00063_, _00062_, _00060_);
  and (_00064_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_36012_[9], _00064_, _00063_);
  or (_00065_, _35143_, _35000_);
  nor (_00066_, _35144_, _34950_);
  and (_00067_, _00066_, _00065_);
  nor (_00068_, _34949_, _31053_);
  or (_00069_, _00068_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00070_, _00069_, _00067_);
  or (_00071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _30491_);
  and (_00072_, _00071_, _35796_);
  and (_36012_[10], _00072_, _00070_);
  nor (_00073_, _35144_, _34997_);
  nor (_00074_, _00073_, _35145_);
  or (_00075_, _00074_, _34950_);
  or (_00076_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00077_, _00076_, _35154_);
  and (_00078_, _00077_, _00075_);
  and (_00079_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_36012_[11], _00079_, _00078_);
  nor (_00080_, _35145_, _34994_);
  nor (_00081_, _00080_, _35146_);
  or (_00082_, _00081_, _34950_);
  or (_00083_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00084_, _00083_, _35154_);
  and (_00085_, _00084_, _00082_);
  and (_00086_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_36012_[12], _00086_, _00085_);
  and (_00087_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_00088_, _35146_, _34992_);
  nor (_00089_, _00088_, _35147_);
  or (_00090_, _00089_, _34950_);
  or (_00091_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00092_, _00091_, _35154_);
  and (_00093_, _00092_, _00090_);
  or (_36012_[13], _00093_, _00087_);
  nor (_00094_, _35147_, _34989_);
  nor (_00095_, _00094_, _35148_);
  or (_00096_, _00095_, _34950_);
  or (_00097_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00098_, _00097_, _35154_);
  and (_00099_, _00098_, _00096_);
  and (_00100_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_36012_[14], _00100_, _00099_);
  and (_36016_[0], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _35796_);
  and (_36016_[1], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _35796_);
  and (_36016_[2], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _35796_);
  and (_36016_[3], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _35796_);
  and (_36016_[4], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _35796_);
  and (_36016_[5], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _35796_);
  and (_36016_[6], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _35796_);
  and (_00101_, _35122_, _30494_);
  nand (_00102_, _00101_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00103_, _00101_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00104_, _00103_, _35154_);
  and (_36017_[0], _00104_, _00102_);
  or (_00105_, _35164_, _35162_);
  and (_00106_, _00105_, _35165_);
  or (_00107_, _00106_, _32110_);
  or (_00108_, _30494_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00109_, _00108_, _35154_);
  and (_36017_[1], _00109_, _00107_);
  and (_00110_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00111_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_00112_, _00111_, _36022_);
  or (_36021_[0], _00112_, _00110_);
  and (_00113_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00114_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00115_, _00114_, _36022_);
  or (_36021_[1], _00115_, _00113_);
  and (_00116_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00117_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00118_, _00117_, _36022_);
  or (_36021_[2], _00118_, _00116_);
  and (_00119_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00120_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00121_, _00120_, _36022_);
  or (_36021_[3], _00121_, _00119_);
  and (_00122_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00123_, _35354_, _36022_);
  or (_36021_[4], _00123_, _00122_);
  and (_00124_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00125_, _35358_, _36022_);
  or (_36021_[5], _00125_, _00124_);
  and (_00126_, _35187_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00127_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00128_, _00127_, _36022_);
  or (_36021_[6], _00128_, _00126_);
  and (_36024_[0], _35195_, _35796_);
  nor (_36024_[1], _35205_, rst);
  and (_36024_[2], _35201_, _35796_);
  and (_00129_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00130_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00131_, _00130_, _00129_);
  and (_36026_[0], _00131_, _35796_);
  and (_00132_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00133_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00134_, _00133_, _00132_);
  and (_36026_[1], _00134_, _35796_);
  and (_00135_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00136_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00137_, _00136_, _00135_);
  and (_36026_[2], _00137_, _35796_);
  and (_00138_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00139_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00140_, _00139_, _00138_);
  and (_36026_[3], _00140_, _35796_);
  and (_00141_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00142_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00143_, _00142_, _00141_);
  and (_36026_[4], _00143_, _35796_);
  and (_00144_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00145_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00146_, _00145_, _00144_);
  and (_36026_[5], _00146_, _35796_);
  and (_00147_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00148_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00149_, _00148_, _00147_);
  and (_36026_[6], _00149_, _35796_);
  and (_00150_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00151_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00152_, _00151_, _00150_);
  and (_36026_[7], _00152_, _35796_);
  and (_00153_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00154_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00155_, _00154_, _00153_);
  and (_36026_[8], _00155_, _35796_);
  and (_00156_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00157_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00158_, _00157_, _00156_);
  and (_36026_[9], _00158_, _35796_);
  and (_00159_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00160_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00161_, _00160_, _00159_);
  and (_36026_[10], _00161_, _35796_);
  and (_00162_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00163_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00164_, _00163_, _00162_);
  and (_36026_[11], _00164_, _35796_);
  and (_00165_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00166_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00167_, _00166_, _00165_);
  and (_36026_[12], _00167_, _35796_);
  and (_00168_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00169_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00170_, _00169_, _00168_);
  and (_36026_[13], _00170_, _35796_);
  and (_00171_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00172_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00173_, _00172_, _00171_);
  and (_36026_[14], _00173_, _35796_);
  and (_00174_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00175_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00176_, _00175_, _00174_);
  and (_36026_[15], _00176_, _35796_);
  and (_00177_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00178_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00179_, _00178_, _00177_);
  and (_36026_[16], _00179_, _35796_);
  and (_00180_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00181_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00182_, _00181_, _00180_);
  and (_36026_[17], _00182_, _35796_);
  and (_00183_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00184_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00185_, _00184_, _00183_);
  and (_36026_[18], _00185_, _35796_);
  and (_00186_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00187_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00188_, _00187_, _00186_);
  and (_36026_[19], _00188_, _35796_);
  and (_00189_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00190_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00191_, _00190_, _00189_);
  and (_36026_[20], _00191_, _35796_);
  and (_00192_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00193_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00194_, _00193_, _00192_);
  and (_36026_[21], _00194_, _35796_);
  and (_00195_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00196_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00197_, _00196_, _00195_);
  and (_36026_[22], _00197_, _35796_);
  and (_00198_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00199_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00200_, _00199_, _00198_);
  and (_36026_[23], _00200_, _35796_);
  and (_00201_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00202_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00203_, _00202_, _00201_);
  and (_36026_[24], _00203_, _35796_);
  and (_00204_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00205_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00206_, _00205_, _00204_);
  and (_36026_[25], _00206_, _35796_);
  and (_00207_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00208_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00209_, _00208_, _00207_);
  and (_36026_[26], _00209_, _35796_);
  and (_00210_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00211_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00212_, _00211_, _00210_);
  and (_36026_[27], _00212_, _35796_);
  and (_00213_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00214_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00215_, _00214_, _00213_);
  and (_36026_[28], _00215_, _35796_);
  and (_00216_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00217_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00218_, _00217_, _00216_);
  and (_36026_[29], _00218_, _35796_);
  and (_00219_, _35209_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00220_, _35211_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00221_, _00220_, _00219_);
  and (_36026_[30], _00221_, _35796_);
  not (_00222_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  nor (_00223_, _35218_, _00222_);
  and (_00224_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_00225_, _00224_, _35218_);
  or (_00226_, _00225_, _00223_);
  and (_36027_[0], _00226_, _35796_);
  not (_00227_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  nor (_00228_, _35218_, _00227_);
  and (_00229_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00230_, _00229_, _35218_);
  or (_00231_, _00230_, _00228_);
  and (_36027_[1], _00231_, _35796_);
  not (_00232_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  nor (_00233_, _35218_, _00232_);
  and (_00234_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00235_, _00234_, _35218_);
  or (_00236_, _00235_, _00233_);
  and (_36027_[2], _00236_, _35796_);
  not (_00237_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  nor (_00238_, _35218_, _00237_);
  and (_00239_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00240_, _00239_, _35218_);
  or (_00241_, _00240_, _00238_);
  and (_36027_[3], _00241_, _35796_);
  not (_00242_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  nor (_00243_, _35218_, _00242_);
  and (_00244_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_00245_, _00244_, _35218_);
  or (_00246_, _00245_, _00243_);
  and (_36027_[4], _00246_, _35796_);
  not (_00247_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  nor (_00248_, _35218_, _00247_);
  and (_00249_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_00250_, _00249_, _35218_);
  or (_00251_, _00250_, _00248_);
  and (_36027_[5], _00251_, _35796_);
  not (_00252_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  nor (_00253_, _35218_, _00252_);
  and (_00254_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00255_, _00254_, _35218_);
  or (_00256_, _00255_, _00253_);
  and (_36027_[6], _00256_, _35796_);
  not (_00257_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  nor (_00258_, _35218_, _00257_);
  or (_00259_, _32225_, _35229_);
  or (_00260_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00261_, _00260_, _35218_);
  and (_00262_, _00261_, _00259_);
  or (_00263_, _00262_, _00258_);
  and (_36030_[0], _00263_, _35796_);
  not (_00264_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  nor (_00265_, _35218_, _00264_);
  or (_00266_, _32443_, _35229_);
  or (_00267_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00268_, _00267_, _35218_);
  and (_00269_, _00268_, _00266_);
  or (_00270_, _00269_, _00265_);
  and (_36030_[1], _00270_, _35796_);
  not (_00271_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  nor (_00272_, _35218_, _00271_);
  or (_00273_, _32329_, _35229_);
  or (_00274_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00275_, _00274_, _35218_);
  and (_00276_, _00275_, _00273_);
  or (_00277_, _00276_, _00272_);
  and (_36030_[2], _00277_, _35796_);
  not (_00278_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  nor (_00279_, _35218_, _00278_);
  or (_00280_, _32173_, _35229_);
  or (_00281_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00282_, _00281_, _35218_);
  and (_00283_, _00282_, _00280_);
  or (_00284_, _00283_, _00279_);
  and (_36030_[3], _00284_, _35796_);
  not (_00285_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  nor (_00286_, _35218_, _00285_);
  or (_00287_, _32382_, _35229_);
  or (_00288_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00289_, _00288_, _35218_);
  and (_00290_, _00289_, _00287_);
  or (_00291_, _00290_, _00286_);
  and (_36030_[4], _00291_, _35796_);
  not (_00292_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  nor (_00293_, _35218_, _00292_);
  nand (_00294_, _32279_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00295_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00296_, _00295_, _35218_);
  and (_00297_, _00296_, _00294_);
  or (_00298_, _00297_, _00293_);
  and (_36030_[5], _00298_, _35796_);
  not (_00299_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  nor (_00300_, _35218_, _00299_);
  nand (_00301_, _32497_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00302_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00303_, _00302_, _35218_);
  and (_00304_, _00303_, _00301_);
  or (_00305_, _00304_, _00300_);
  and (_36030_[6], _00305_, _35796_);
  not (_00306_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  nor (_00307_, _35218_, _00306_);
  or (_00308_, _32105_, _35229_);
  or (_00309_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00310_, _00309_, _35218_);
  and (_00311_, _00310_, _00308_);
  or (_00312_, _00311_, _00307_);
  and (_36030_[7], _00312_, _35796_);
  not (_00313_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  nor (_00314_, _35218_, _00313_);
  and (_00315_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_00316_, _00315_, _35218_);
  or (_00317_, _00316_, _00314_);
  and (_36030_[8], _00317_, _35796_);
  not (_00318_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  nor (_00319_, _35218_, _00318_);
  and (_00320_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_00321_, _00320_, _35218_);
  or (_00322_, _00321_, _00319_);
  and (_36030_[9], _00322_, _35796_);
  not (_00323_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  nor (_00324_, _35218_, _00323_);
  and (_00325_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_00326_, _00325_, _35218_);
  or (_00327_, _00326_, _00324_);
  and (_36030_[10], _00327_, _35796_);
  not (_00328_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  nor (_00329_, _35218_, _00328_);
  and (_00330_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_00331_, _00330_, _35218_);
  or (_00332_, _00331_, _00329_);
  and (_36030_[11], _00332_, _35796_);
  not (_00333_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  nor (_00334_, _35218_, _00333_);
  and (_00335_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_00336_, _00335_, _35218_);
  or (_00337_, _00336_, _00334_);
  and (_36030_[12], _00337_, _35796_);
  not (_00338_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  nor (_00339_, _35218_, _00338_);
  and (_00340_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_00341_, _00340_, _35218_);
  or (_00342_, _00341_, _00339_);
  and (_36030_[13], _00342_, _35796_);
  not (_00343_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  nor (_00344_, _35218_, _00343_);
  and (_00345_, _35229_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_00346_, _00345_, _35218_);
  or (_00347_, _00346_, _00344_);
  and (_36030_[14], _00347_, _35796_);
  nand (_00348_, _35235_, _28739_);
  or (_00349_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00350_, _00349_, _35796_);
  and (_36034_[0], _00350_, _00348_);
  nand (_00351_, _35235_, _29380_);
  or (_00352_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00353_, _00352_, _35796_);
  and (_36034_[1], _00353_, _00351_);
  nand (_00354_, _35235_, _30024_);
  or (_00355_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00356_, _00355_, _35796_);
  and (_36034_[2], _00356_, _00354_);
  nand (_00357_, _35235_, _30247_);
  or (_00358_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00359_, _00358_, _35796_);
  and (_36034_[3], _00359_, _00357_);
  nand (_00360_, _35235_, _30319_);
  or (_00361_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00362_, _00361_, _35796_);
  and (_36034_[4], _00362_, _00360_);
  nand (_00363_, _35235_, _30396_);
  or (_00364_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00365_, _00364_, _35796_);
  and (_36034_[5], _00365_, _00363_);
  nand (_00366_, _35235_, _30468_);
  or (_00367_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00368_, _00367_, _35796_);
  and (_36034_[6], _00368_, _00366_);
  nand (_00369_, _35235_, _27635_);
  or (_00370_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00371_, _00370_, _35796_);
  and (_36034_[7], _00371_, _00369_);
  nand (_00372_, _35235_, _31157_);
  or (_00373_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00374_, _00373_, _35796_);
  and (_36034_[8], _00374_, _00372_);
  nand (_00375_, _35235_, _31189_);
  or (_00376_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00377_, _00376_, _35796_);
  and (_36034_[9], _00377_, _00375_);
  nand (_00378_, _35235_, _31219_);
  or (_00379_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00380_, _00379_, _35796_);
  and (_36034_[10], _00380_, _00378_);
  nand (_00381_, _35235_, _31250_);
  or (_00382_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00383_, _00382_, _35796_);
  and (_36034_[11], _00383_, _00381_);
  nand (_00384_, _35235_, _31281_);
  or (_00385_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00386_, _00385_, _35796_);
  and (_36034_[12], _00386_, _00384_);
  nand (_00387_, _35235_, _31315_);
  or (_00388_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00389_, _00388_, _35796_);
  and (_36034_[13], _00389_, _00387_);
  nand (_00390_, _35235_, _31344_);
  or (_00391_, _35235_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00392_, _00391_, _35796_);
  and (_36034_[14], _00392_, _00390_);
  nor (_35999_, _32148_, rst);
  nor (_00393_, _32203_, _32133_);
  and (_00394_, _00393_, _32521_);
  and (_00395_, _00393_, _32413_);
  nor (_00396_, _32521_, _32305_);
  and (_00397_, _00396_, _00395_);
  nor (_00398_, _32521_, _32133_);
  and (_00399_, _32414_, _32305_);
  and (_00400_, _00399_, _32202_);
  and (_00401_, _00400_, _00398_);
  and (_00402_, _00393_, _32414_);
  and (_00403_, _00396_, _00402_);
  or (_00404_, _00403_, _00401_);
  or (_00405_, _00404_, _00397_);
  nor (_00406_, _00405_, _00394_);
  not (_00407_, _31385_);
  and (_00408_, _30761_, _30756_);
  or (_00409_, _00408_, _34207_);
  nor (_00410_, _00409_, _30771_);
  nor (_00411_, _30826_, _30789_);
  and (_00412_, _00411_, _00410_);
  not (_00413_, _34203_);
  nor (_00414_, _00413_, _34145_);
  and (_00415_, _00414_, _00412_);
  and (_00416_, _30792_, _30734_);
  or (_00417_, _34324_, _34147_);
  or (_00418_, _00417_, _00416_);
  nor (_00419_, _00418_, _34470_);
  and (_00420_, _00419_, _00415_);
  and (_00421_, _00420_, _30815_);
  nor (_00422_, _00421_, _30490_);
  not (_00423_, _00422_);
  and (_00424_, _00423_, _00394_);
  nor (_00425_, _00424_, _00407_);
  nand (_00426_, _00425_, _34681_);
  nor (_00427_, _00426_, _00406_);
  not (_00428_, _32354_);
  nor (_00429_, _31534_, _31522_);
  and (_00430_, _31534_, _31522_);
  nor (_00431_, _00430_, _00429_);
  nor (_00432_, _31562_, _31546_);
  and (_00433_, _31562_, _31546_);
  nor (_00434_, _00433_, _00432_);
  nor (_00435_, _00434_, _00431_);
  and (_00436_, _00434_, _00431_);
  or (_00437_, _00436_, _00435_);
  nor (_00438_, _31586_, _31574_);
  and (_00439_, _31586_, _31574_);
  nor (_00440_, _00439_, _00438_);
  not (_00441_, _31510_);
  nor (_00442_, _31598_, _00441_);
  and (_00443_, _31598_, _00441_);
  nor (_00444_, _00443_, _00442_);
  nor (_00445_, _00444_, _00440_);
  and (_00446_, _00444_, _00440_);
  or (_00447_, _00446_, _00445_);
  or (_00448_, _00447_, _00437_);
  nand (_00449_, _00447_, _00437_);
  and (_00450_, _00449_, _00448_);
  or (_00451_, _00450_, _00428_);
  and (_00452_, _32250_, _32463_);
  or (_00453_, _32354_, _31455_);
  and (_00454_, _00453_, _00452_);
  and (_00455_, _00454_, _00451_);
  or (_00456_, _32354_, _31464_);
  not (_00457_, _32250_);
  and (_00458_, _00457_, _32463_);
  or (_00459_, _00428_, _31399_);
  and (_00460_, _00459_, _00458_);
  and (_00461_, _00460_, _00456_);
  nor (_00462_, _32250_, _32463_);
  and (_00463_, _00462_, _00428_);
  and (_00464_, _00463_, _31390_);
  and (_00465_, _00462_, _32354_);
  and (_00466_, _00465_, _31445_);
  or (_00467_, _00466_, _00464_);
  or (_00468_, _00467_, _00461_);
  or (_00469_, _00428_, _31434_);
  nor (_00470_, _00457_, _32463_);
  or (_00471_, _32354_, _31480_);
  and (_00472_, _00471_, _00470_);
  and (_00473_, _00472_, _00469_);
  or (_00474_, _00473_, _00468_);
  or (_00475_, _00474_, _00455_);
  and (_00476_, _00475_, _00401_);
  and (_00477_, _34659_, p0in_reg[7]);
  and (_00478_, _34655_, p0_in[7]);
  or (_00479_, _00478_, _00477_);
  or (_00480_, _00479_, _00422_);
  nand (_00481_, _00422_, _31609_);
  and (_00482_, _00481_, _00480_);
  and (_00483_, _00482_, _00463_);
  and (_00484_, _34659_, p0in_reg[3]);
  and (_00485_, _34655_, p0_in[3]);
  or (_00486_, _00485_, _00484_);
  or (_00487_, _00486_, _00422_);
  or (_00488_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_00489_, _00488_, _00487_);
  and (_00490_, _00489_, _00465_);
  or (_00491_, _00490_, _00483_);
  and (_00492_, _34659_, p0in_reg[4]);
  and (_00493_, _34655_, p0_in[4]);
  or (_00494_, _00493_, _00492_);
  or (_00495_, _00494_, _00422_);
  or (_00496_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_00497_, _00496_, _00495_);
  or (_00498_, _00497_, _32354_);
  and (_00499_, _34659_, p0in_reg[0]);
  and (_00500_, _34655_, p0_in[0]);
  or (_00501_, _00500_, _00499_);
  or (_00502_, _00501_, _00422_);
  nand (_00503_, _00422_, _31671_);
  and (_00504_, _00503_, _00502_);
  or (_00505_, _00504_, _00428_);
  and (_00506_, _00505_, _00452_);
  and (_00507_, _00506_, _00498_);
  and (_00508_, _34659_, p0in_reg[6]);
  and (_00509_, _34655_, p0_in[6]);
  or (_00510_, _00509_, _00508_);
  or (_00511_, _00510_, _00422_);
  nand (_00512_, _00422_, _31743_);
  and (_00513_, _00512_, _00511_);
  and (_00514_, _00513_, _00428_);
  and (_00515_, _34659_, p0in_reg[2]);
  and (_00516_, _34655_, p0_in[2]);
  or (_00517_, _00516_, _00515_);
  or (_00518_, _00517_, _00422_);
  nand (_00519_, _00422_, _31698_);
  and (_00520_, _00519_, _00518_);
  and (_00521_, _00520_, _32354_);
  or (_00522_, _00521_, _00514_);
  and (_00523_, _00522_, _00470_);
  and (_00524_, _34659_, p0in_reg[5]);
  and (_00525_, _34655_, p0_in[5]);
  or (_00526_, _00525_, _00524_);
  or (_00527_, _00526_, _00422_);
  or (_00528_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_00529_, _00528_, _00527_);
  and (_00530_, _00529_, _00428_);
  and (_00531_, _34659_, p0in_reg[1]);
  and (_00532_, _34655_, p0_in[1]);
  or (_00533_, _00532_, _00531_);
  or (_00534_, _00533_, _00422_);
  nand (_00535_, _00422_, _31682_);
  and (_00536_, _00535_, _00534_);
  and (_00537_, _00536_, _32354_);
  or (_00538_, _00537_, _00530_);
  and (_00539_, _00538_, _00458_);
  or (_00540_, _00539_, _00523_);
  or (_00541_, _00540_, _00507_);
  or (_00542_, _00541_, _00491_);
  and (_00543_, _32413_, _32305_);
  and (_00544_, _00543_, _00542_);
  and (_00545_, _34659_, p1in_reg[3]);
  and (_00546_, _34655_, p1_in[3]);
  or (_00547_, _00546_, _00545_);
  or (_00548_, _00547_, _00422_);
  or (_00549_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00550_, _00549_, _00548_);
  and (_00551_, _00550_, _00465_);
  and (_00552_, _34659_, p1in_reg[7]);
  and (_00553_, _34655_, p1_in[7]);
  or (_00554_, _00553_, _00552_);
  or (_00555_, _00554_, _00422_);
  nand (_00556_, _00422_, _31622_);
  and (_00557_, _00556_, _00555_);
  and (_00558_, _00557_, _00463_);
  or (_00559_, _00558_, _00551_);
  and (_00560_, _34659_, p1in_reg[4]);
  and (_00561_, _34655_, p1_in[4]);
  or (_00562_, _00561_, _00560_);
  or (_00563_, _00562_, _00422_);
  or (_00564_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_00565_, _00564_, _00563_);
  or (_00566_, _00565_, _32354_);
  and (_00567_, _34659_, p1in_reg[0]);
  and (_00568_, _34655_, p1_in[0]);
  or (_00569_, _00568_, _00567_);
  or (_00570_, _00569_, _00422_);
  nand (_00571_, _00422_, _31761_);
  and (_00572_, _00571_, _00570_);
  or (_00573_, _00572_, _00428_);
  and (_00574_, _00573_, _00452_);
  and (_00575_, _00574_, _00566_);
  and (_00576_, _34659_, p1in_reg[6]);
  and (_00577_, _34655_, p1_in[6]);
  or (_00578_, _00577_, _00576_);
  or (_00579_, _00578_, _00422_);
  nand (_00580_, _00422_, _31836_);
  and (_00581_, _00580_, _00579_);
  and (_00582_, _00581_, _00428_);
  and (_00583_, _34659_, p1in_reg[2]);
  and (_00584_, _34655_, p1_in[2]);
  or (_00585_, _00584_, _00583_);
  or (_00586_, _00585_, _00422_);
  nand (_00587_, _00422_, _31787_);
  and (_00588_, _00587_, _00586_);
  and (_00589_, _00588_, _32354_);
  or (_00590_, _00589_, _00582_);
  and (_00591_, _00590_, _00470_);
  or (_00592_, _00591_, _00575_);
  and (_00593_, _34659_, p1in_reg[5]);
  and (_00594_, _34655_, p1_in[5]);
  or (_00595_, _00594_, _00593_);
  or (_00596_, _00595_, _00422_);
  or (_00597_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_00598_, _00597_, _00596_);
  and (_00599_, _00598_, _00428_);
  and (_00600_, _34659_, p1in_reg[1]);
  and (_00601_, _34655_, p1_in[1]);
  or (_00602_, _00601_, _00600_);
  or (_00603_, _00602_, _00422_);
  nand (_00604_, _00422_, _31774_);
  and (_00605_, _00604_, _00603_);
  and (_00606_, _00605_, _32354_);
  or (_00607_, _00606_, _00599_);
  and (_00608_, _00607_, _00458_);
  or (_00609_, _00608_, _00592_);
  or (_00610_, _00609_, _00559_);
  and (_00611_, _00610_, _00399_);
  or (_00612_, _00611_, _00544_);
  and (_00613_, _00612_, _00394_);
  and (_00614_, _32521_, _32306_);
  and (_00615_, _34659_, p3in_reg[7]);
  and (_00616_, _34655_, p3_in[7]);
  or (_00617_, _00616_, _00615_);
  or (_00618_, _00617_, _00422_);
  nand (_00619_, _00422_, _31648_);
  and (_00620_, _00619_, _00618_);
  and (_00621_, _00620_, _00463_);
  and (_00622_, _34659_, p3in_reg[4]);
  and (_00623_, _34655_, p3_in[4]);
  or (_00624_, _00623_, _00622_);
  or (_00625_, _00624_, _00422_);
  or (_00626_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_00627_, _00626_, _00625_);
  or (_00628_, _00627_, _32354_);
  and (_00629_, _34659_, p3in_reg[0]);
  and (_00630_, _34655_, p3_in[0]);
  or (_00631_, _00630_, _00629_);
  or (_00632_, _00631_, _00422_);
  nand (_00633_, _00422_, _31934_);
  and (_00634_, _00633_, _00632_);
  or (_00635_, _00634_, _00428_);
  and (_00636_, _00635_, _00452_);
  and (_00637_, _00636_, _00628_);
  and (_00638_, _34659_, p3in_reg[3]);
  and (_00639_, _34655_, p3_in[3]);
  or (_00640_, _00639_, _00638_);
  or (_00641_, _00640_, _00422_);
  or (_00642_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_00643_, _00642_, _00641_);
  and (_00644_, _00643_, _00465_);
  or (_00645_, _00644_, _00637_);
  or (_00646_, _00645_, _00621_);
  and (_00647_, _34659_, p3in_reg[6]);
  and (_00648_, _34655_, p3_in[6]);
  or (_00649_, _00648_, _00647_);
  or (_00650_, _00649_, _00422_);
  nand (_00651_, _00422_, _32014_);
  and (_00652_, _00651_, _00650_);
  and (_00653_, _00652_, _00428_);
  and (_00654_, _34659_, p3in_reg[2]);
  and (_00655_, _34655_, p3_in[2]);
  or (_00656_, _00655_, _00654_);
  or (_00657_, _00656_, _00422_);
  nand (_00658_, _00422_, _31960_);
  and (_00659_, _00658_, _00657_);
  and (_00660_, _00659_, _32354_);
  or (_00661_, _00660_, _00653_);
  and (_00662_, _00661_, _00470_);
  and (_00663_, _34659_, p3in_reg[5]);
  and (_00664_, _34655_, p3_in[5]);
  or (_00665_, _00664_, _00663_);
  or (_00666_, _00665_, _00422_);
  or (_00667_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00668_, _00667_, _00666_);
  and (_00669_, _00668_, _00428_);
  and (_00670_, _34659_, p3in_reg[1]);
  and (_00671_, _34655_, p3_in[1]);
  or (_00672_, _00671_, _00670_);
  or (_00673_, _00672_, _00422_);
  nand (_00674_, _00422_, _31949_);
  and (_00675_, _00674_, _00673_);
  and (_00676_, _00675_, _32354_);
  or (_00677_, _00676_, _00669_);
  and (_00678_, _00677_, _00458_);
  or (_00679_, _00678_, _00662_);
  or (_00680_, _00679_, _00646_);
  and (_00681_, _00680_, _00402_);
  and (_00682_, _34659_, p2in_reg[7]);
  and (_00683_, _34655_, p2_in[7]);
  or (_00684_, _00683_, _00682_);
  or (_00685_, _00684_, _00422_);
  nand (_00686_, _00422_, _31640_);
  and (_00687_, _00686_, _00685_);
  and (_00688_, _00687_, _00463_);
  and (_00689_, _34659_, p2in_reg[4]);
  and (_00690_, _34655_, p2_in[4]);
  or (_00691_, _00690_, _00689_);
  or (_00692_, _00691_, _00422_);
  or (_00693_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_00694_, _00693_, _00692_);
  or (_00695_, _00694_, _32354_);
  and (_00696_, _34659_, p2in_reg[0]);
  and (_00697_, _34655_, p2_in[0]);
  or (_00698_, _00697_, _00696_);
  or (_00699_, _00698_, _00422_);
  nand (_00700_, _00422_, _31848_);
  and (_00701_, _00700_, _00699_);
  or (_00702_, _00701_, _00428_);
  and (_00703_, _00702_, _00452_);
  and (_00704_, _00703_, _00695_);
  and (_00705_, _34659_, p2in_reg[3]);
  and (_00706_, _34655_, p2_in[3]);
  or (_00707_, _00706_, _00705_);
  or (_00708_, _00707_, _00422_);
  or (_00709_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00710_, _00709_, _00708_);
  and (_00711_, _00710_, _00465_);
  or (_00712_, _00711_, _00704_);
  or (_00713_, _00712_, _00688_);
  and (_00714_, _34659_, p2in_reg[6]);
  and (_00715_, _34655_, p2_in[6]);
  or (_00716_, _00715_, _00714_);
  or (_00717_, _00716_, _00422_);
  nand (_00718_, _00422_, _31923_);
  and (_00719_, _00718_, _00717_);
  and (_00720_, _00719_, _00428_);
  and (_00721_, _34659_, p2in_reg[2]);
  and (_00722_, _34655_, p2_in[2]);
  or (_00723_, _00722_, _00721_);
  or (_00724_, _00723_, _00422_);
  nand (_00725_, _00422_, _31874_);
  and (_00726_, _00725_, _00724_);
  and (_00727_, _00726_, _32354_);
  or (_00728_, _00727_, _00720_);
  and (_00729_, _00728_, _00470_);
  and (_00730_, _34659_, p2in_reg[5]);
  and (_00731_, _34655_, p2_in[5]);
  or (_00732_, _00731_, _00730_);
  or (_00733_, _00732_, _00422_);
  or (_00734_, _00423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_00735_, _00734_, _00733_);
  and (_00736_, _00735_, _00428_);
  and (_00737_, _34659_, p2in_reg[1]);
  and (_00738_, _34655_, p2_in[1]);
  or (_00739_, _00738_, _00737_);
  or (_00740_, _00739_, _00422_);
  nand (_00741_, _00422_, _31861_);
  and (_00742_, _00741_, _00740_);
  and (_00743_, _00742_, _32354_);
  or (_00744_, _00743_, _00736_);
  and (_00745_, _00744_, _00458_);
  or (_00746_, _00745_, _00729_);
  or (_00747_, _00746_, _00713_);
  and (_00748_, _00747_, _00395_);
  or (_00749_, _00748_, _00681_);
  and (_00750_, _00749_, _00614_);
  and (_00751_, _00463_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_00752_, _32354_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_00753_, _32354_, _28772_);
  and (_00754_, _00753_, _00452_);
  and (_00755_, _00754_, _00752_);
  and (_00756_, _00465_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00757_, _00756_, _00755_);
  or (_00758_, _00757_, _00751_);
  nor (_00759_, _32354_, _30471_);
  and (_00760_, _32354_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00761_, _00760_, _00759_);
  and (_00762_, _00761_, _00470_);
  nor (_00763_, _32354_, _30399_);
  and (_00764_, _32354_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_00765_, _00764_, _00763_);
  and (_00766_, _00765_, _00458_);
  or (_00767_, _00766_, _00762_);
  or (_00768_, _00767_, _00758_);
  and (_00769_, _00768_, _00403_);
  and (_00770_, _00428_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_00771_, _32354_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00772_, _00771_, _00770_);
  and (_00773_, _00772_, _00452_);
  and (_00774_, _00458_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00775_, _00774_, _00428_);
  and (_00776_, _00470_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00777_, _00462_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00778_, _00777_, _00776_);
  or (_00779_, _00778_, _00775_);
  and (_00780_, _00458_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00781_, _00780_, _32354_);
  and (_00782_, _00470_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00783_, _00462_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_00784_, _00783_, _00782_);
  or (_00785_, _00784_, _00781_);
  and (_00786_, _00785_, _00779_);
  or (_00787_, _00786_, _00773_);
  and (_00788_, _00787_, _00397_);
  nor (_00789_, _00406_, _27668_);
  and (_00790_, _00789_, _34694_);
  or (_00791_, _00790_, _00788_);
  or (_00792_, _00791_, _00769_);
  or (_00793_, _00792_, _00750_);
  or (_00794_, _00793_, _00613_);
  or (_00795_, _00794_, _00476_);
  and (_00796_, _00790_, _28243_);
  and (_00797_, _00397_, _31486_);
  nor (_00798_, _00797_, _00796_);
  and (_00799_, _00798_, _00795_);
  and (_00800_, _00452_, _31522_);
  and (_00801_, _00458_, _31534_);
  not (_00802_, _00462_);
  nor (_00803_, _00802_, _31562_);
  and (_00804_, _00470_, _31546_);
  or (_00805_, _00804_, _00803_);
  or (_00806_, _00805_, _00801_);
  or (_00807_, _00806_, _00800_);
  and (_00808_, _00807_, _32354_);
  and (_00809_, _00463_, _31510_);
  and (_00810_, _00452_, _31574_);
  and (_00811_, _00470_, _31598_);
  and (_00812_, _00458_, _31586_);
  or (_00813_, _00812_, _00811_);
  or (_00814_, _00813_, _00810_);
  and (_00815_, _00814_, _00428_);
  or (_00816_, _00815_, _00809_);
  or (_00817_, _00816_, _00808_);
  and (_00818_, _00817_, _00797_);
  nor (_00819_, _00818_, _00799_);
  nor (_00820_, _00819_, _00427_);
  or (_00821_, _32354_, _32474_);
  nand (_00822_, _32354_, _30947_);
  and (_00823_, _00822_, _00470_);
  and (_00824_, _00823_, _00821_);
  or (_00825_, _32354_, _32361_);
  nand (_00826_, _32354_, _30962_);
  and (_00827_, _00826_, _00452_);
  and (_00828_, _00827_, _00825_);
  or (_00829_, _00828_, _00824_);
  and (_00830_, _00465_, _32151_);
  and (_00831_, _00463_, _30908_);
  nor (_00832_, _00428_, _30954_);
  nor (_00833_, _32354_, _30925_);
  or (_00834_, _00833_, _00832_);
  and (_00835_, _00834_, _00458_);
  or (_00836_, _00835_, _00831_);
  or (_00837_, _00836_, _00830_);
  or (_00838_, _00837_, _00829_);
  and (_00839_, _00838_, _00427_);
  or (_00840_, _00839_, _00820_);
  and (_36135_, _00840_, _35796_);
  not (_00841_, _32133_);
  and (_00842_, _32521_, _00841_);
  and (_00843_, _00543_, _00842_);
  and (_00844_, _32202_, _32354_);
  and (_00845_, _00844_, _00462_);
  and (_00846_, _00845_, _00843_);
  and (_00847_, _00846_, _31029_);
  and (_00848_, _00844_, _00452_);
  and (_00849_, _00848_, _00398_);
  and (_00850_, _00849_, _00399_);
  and (_00851_, _00850_, _31380_);
  nor (_00852_, _00851_, _00847_);
  nor (_00853_, _00852_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_00854_, _00853_);
  not (_00855_, _31438_);
  nor (_00856_, _00463_, _00855_);
  and (_00857_, _00856_, _34681_);
  or (_00858_, _31486_, _31482_);
  nor (_00859_, _32414_, _32305_);
  and (_00860_, _00859_, _00849_);
  and (_00861_, _00860_, _00858_);
  nor (_00862_, _00861_, _00857_);
  and (_00863_, _00862_, _34697_);
  and (_00864_, _00863_, _00854_);
  and (_00865_, _00844_, _00470_);
  and (_00866_, _00865_, _00843_);
  and (_00867_, _00866_, _31029_);
  or (_00868_, _00867_, rst);
  nor (_36136_, _00868_, _00864_);
  nand (_00869_, _00867_, _27635_);
  or (_00870_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_00871_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_00872_, _00850_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_00873_, _00872_, _00871_);
  and (_00874_, _00848_, _00842_);
  and (_00875_, _00874_, _00399_);
  and (_00876_, _00875_, _00557_);
  and (_00877_, _00874_, _00859_);
  and (_00878_, _00877_, _00687_);
  or (_00879_, _00878_, _00876_);
  or (_00880_, _00879_, _00873_);
  and (_00881_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00882_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_00883_, _00882_, _00881_);
  and (_00884_, _00844_, _00458_);
  and (_00885_, _00884_, _00843_);
  and (_00886_, _00885_, _32130_);
  and (_00887_, _00848_, _00843_);
  and (_00888_, _00887_, _00482_);
  or (_00889_, _00888_, _00886_);
  or (_00890_, _00889_, _00883_);
  nor (_00891_, _32413_, _32305_);
  and (_00892_, _00891_, _00849_);
  and (_00893_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_00894_, _00891_, _00874_);
  and (_00895_, _00894_, _00620_);
  or (_00896_, _00895_, _00893_);
  or (_00897_, _00896_, _00890_);
  nor (_00898_, _00897_, _00880_);
  nand (_00899_, _00898_, _00864_);
  and (_00900_, _00899_, _00870_);
  or (_00901_, _00900_, _00867_);
  and (_00902_, _00901_, _35796_);
  and (_36137_[7], _00902_, _00869_);
  and (_00903_, _00850_, _00450_);
  and (_00904_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00905_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_00906_, _00877_, _00701_);
  or (_00907_, _00906_, _00905_);
  or (_00908_, _00907_, _00904_);
  and (_00909_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_00910_, _00885_, _32228_);
  or (_00911_, _00910_, _00909_);
  and (_00912_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00913_, _00887_, _00504_);
  or (_00914_, _00913_, _00912_);
  or (_00916_, _00914_, _00911_);
  and (_00917_, _00875_, _00572_);
  and (_00918_, _00894_, _00634_);
  or (_00919_, _00918_, _00917_);
  or (_00920_, _00919_, _00916_);
  nor (_00921_, _00920_, _00908_);
  nand (_00922_, _00921_, _00864_);
  or (_00923_, _00922_, _00903_);
  or (_00924_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_00925_, _00924_, _00923_);
  or (_00926_, _00925_, _00867_);
  nand (_00927_, _00867_, _28739_);
  and (_00928_, _00927_, _35796_);
  and (_36137_[0], _00928_, _00926_);
  nand (_00929_, _00867_, _29380_);
  or (_00930_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_00931_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00932_, _00850_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_00933_, _00932_, _00931_);
  and (_00934_, _00875_, _00605_);
  and (_00935_, _00877_, _00742_);
  or (_00936_, _00935_, _00934_);
  or (_00937_, _00936_, _00933_);
  and (_00938_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00939_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00940_, _00939_, _00938_);
  and (_00941_, _00885_, _32417_);
  and (_00942_, _00887_, _00536_);
  or (_00943_, _00942_, _00941_);
  or (_00944_, _00943_, _00940_);
  and (_00946_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00947_, _00894_, _00675_);
  or (_00948_, _00947_, _00946_);
  or (_00949_, _00948_, _00944_);
  nor (_00950_, _00949_, _00937_);
  nand (_00951_, _00950_, _00864_);
  and (_00952_, _00951_, _00930_);
  or (_00953_, _00952_, _00867_);
  and (_00954_, _00953_, _35796_);
  and (_36137_[1], _00954_, _00929_);
  nand (_00955_, _00867_, _30024_);
  or (_00956_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_00957_, _00850_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_00958_, _00875_, _00588_);
  or (_00959_, _00958_, _00957_);
  and (_00960_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00961_, _00894_, _00659_);
  or (_00962_, _00961_, _00960_);
  or (_00963_, _00962_, _00959_);
  and (_00964_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00966_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00967_, _00966_, _00964_);
  and (_00968_, _00885_, _32332_);
  and (_00969_, _00887_, _00520_);
  or (_00970_, _00969_, _00968_);
  or (_00971_, _00970_, _00967_);
  and (_00972_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00973_, _00877_, _00726_);
  or (_00974_, _00973_, _00972_);
  or (_00975_, _00974_, _00971_);
  nor (_00976_, _00975_, _00963_);
  nand (_00977_, _00976_, _00864_);
  and (_00978_, _00977_, _00956_);
  or (_00979_, _00978_, _00867_);
  and (_00980_, _00979_, _35796_);
  and (_36137_[2], _00980_, _00955_);
  nand (_00981_, _00867_, _30247_);
  or (_00982_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_00983_, _00850_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_00984_, _00875_, _00550_);
  or (_00985_, _00984_, _00983_);
  and (_00986_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00987_, _00877_, _00710_);
  or (_00988_, _00987_, _00986_);
  or (_00989_, _00988_, _00985_);
  and (_00990_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00991_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00992_, _00991_, _00990_);
  and (_00993_, _00885_, _32176_);
  and (_00994_, _00887_, _00489_);
  or (_00995_, _00994_, _00993_);
  or (_00996_, _00995_, _00992_);
  and (_00997_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00998_, _00894_, _00643_);
  or (_00999_, _00998_, _00997_);
  or (_01000_, _00999_, _00996_);
  nor (_01001_, _01000_, _00989_);
  nand (_01002_, _01001_, _00864_);
  and (_01003_, _01002_, _00982_);
  or (_01004_, _01003_, _00867_);
  and (_01005_, _01004_, _35796_);
  and (_36137_[3], _01005_, _00981_);
  nand (_01006_, _00867_, _30319_);
  or (_01007_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_01008_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01009_, _00850_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_01010_, _01009_, _01008_);
  and (_01011_, _00875_, _00565_);
  and (_01012_, _00894_, _00627_);
  or (_01013_, _01012_, _01011_);
  or (_01014_, _01013_, _01010_);
  and (_01015_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01016_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01017_, _01016_, _01015_);
  and (_01018_, _00885_, _32385_);
  and (_01019_, _00887_, _00497_);
  or (_01020_, _01019_, _01018_);
  or (_01021_, _01020_, _01017_);
  and (_01022_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01023_, _00877_, _00694_);
  or (_01024_, _01023_, _01022_);
  or (_01025_, _01024_, _01021_);
  nor (_01026_, _01025_, _01014_);
  nand (_01027_, _01026_, _00864_);
  and (_01028_, _01027_, _01007_);
  or (_01029_, _01028_, _00867_);
  and (_01030_, _01029_, _35796_);
  and (_36137_[4], _01030_, _01006_);
  nand (_01031_, _00867_, _30396_);
  or (_01032_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_01033_, _00850_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01034_, _00875_, _00598_);
  or (_01035_, _01034_, _01033_);
  and (_01036_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01037_, _00894_, _00668_);
  or (_01038_, _01037_, _01036_);
  or (_01039_, _01038_, _01035_);
  and (_01040_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_01041_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_01042_, _01041_, _01040_);
  and (_01043_, _00885_, _32282_);
  and (_01044_, _00887_, _00529_);
  or (_01045_, _01044_, _01043_);
  or (_01046_, _01045_, _01042_);
  and (_01047_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01048_, _00877_, _00735_);
  or (_01049_, _01048_, _01047_);
  or (_01050_, _01049_, _01046_);
  nor (_01051_, _01050_, _01039_);
  nand (_01052_, _01051_, _00864_);
  and (_01053_, _01052_, _01032_);
  or (_01054_, _01053_, _00867_);
  and (_01055_, _01054_, _35796_);
  and (_36137_[5], _01055_, _01031_);
  nand (_01056_, _00867_, _30468_);
  or (_01057_, _00864_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_01058_, _00850_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01059_, _00894_, _00652_);
  or (_01060_, _01059_, _01058_);
  and (_01061_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01062_, _00875_, _00581_);
  or (_01063_, _01062_, _01061_);
  or (_01064_, _01063_, _01060_);
  and (_01065_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_01066_, _00887_, _00513_);
  or (_01067_, _01066_, _01065_);
  and (_01068_, _00866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01069_, _00885_, _32499_);
  or (_01070_, _01069_, _01068_);
  or (_01071_, _01070_, _01067_);
  and (_01072_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01073_, _00877_, _00719_);
  or (_01074_, _01073_, _01072_);
  or (_01075_, _01074_, _01071_);
  nor (_01076_, _01075_, _01064_);
  nand (_01077_, _01076_, _00864_);
  and (_01078_, _01077_, _01057_);
  or (_01079_, _01078_, _00867_);
  and (_01080_, _01079_, _35796_);
  and (_36137_[6], _01080_, _01056_);
  and (_36036_, _32529_, _35796_);
  nor (_36037_[7], _32064_, rst);
  nor (_36039_[2], _32354_, rst);
  and (_36037_[0], _32212_, _35796_);
  nor (_36037_[1], _32430_, rst);
  and (_36037_[2], _32317_, _35796_);
  and (_36037_[3], _32160_, _35796_);
  and (_36037_[4], _32370_, _35796_);
  nor (_36037_[5], _32266_, rst);
  nor (_36037_[6], _32484_, rst);
  nor (_36039_[0], _32250_, rst);
  nor (_36039_[1], _32463_, rst);
  not (_01081_, _33486_);
  nor (_01082_, _35506_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01083_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01084_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01083_);
  nor (_01085_, _01084_, _01082_);
  not (_01086_, _01085_);
  nor (_01087_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01088_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01083_);
  nor (_01089_, _01088_, _01087_);
  nor (_01090_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01091_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01083_);
  nor (_01092_, _01091_, _01090_);
  nor (_01093_, _01092_, _01089_);
  not (_01094_, _01093_);
  nor (_01095_, _35488_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01083_);
  nor (_01097_, _01096_, _01095_);
  and (_01098_, _01097_, _01094_);
  nor (_01099_, _01097_, _01094_);
  nor (_01100_, _01099_, _01098_);
  and (_01101_, _01100_, _01086_);
  not (_01102_, _01089_);
  nor (_01103_, _01092_, _01102_);
  and (_01104_, _01103_, _01101_);
  and (_01105_, _01104_, _01081_);
  not (_01106_, _33361_);
  and (_01107_, _01092_, _01102_);
  or (_01108_, _01085_, _01099_);
  or (_01109_, _01086_, _01098_);
  and (_01110_, _01109_, _01108_);
  and (_01111_, _01110_, _01107_);
  and (_01112_, _01111_, _01106_);
  or (_01113_, _01112_, _01105_);
  not (_01114_, _33888_);
  and (_01115_, _01100_, _01085_);
  and (_01116_, _01115_, _01107_);
  and (_01117_, _01116_, _01114_);
  not (_01118_, _33847_);
  and (_01119_, _01115_, _01103_);
  and (_01120_, _01119_, _01118_);
  or (_01121_, _01120_, _01117_);
  or (_01122_, _01121_, _01113_);
  not (_01123_, _33568_);
  and (_01124_, _01092_, _01089_);
  and (_01125_, _01124_, _01101_);
  and (_01126_, _01125_, _01123_);
  not (_01127_, _33402_);
  and (_01128_, _01110_, _01124_);
  and (_01129_, _01128_, _01127_);
  or (_01130_, _01129_, _01126_);
  not (_01131_, _33297_);
  and (_01132_, _01110_, _01103_);
  and (_01133_, _01132_, _01131_);
  not (_01134_, _33929_);
  and (_01135_, _01115_, _01124_);
  and (_01136_, _01135_, _01134_);
  or (_01137_, _01136_, _01133_);
  or (_01138_, _01137_, _01130_);
  not (_01139_, _33650_);
  and (_01140_, _01086_, _01097_);
  and (_01141_, _01140_, _01103_);
  and (_01142_, _01141_, _01139_);
  not (_01143_, _33697_);
  and (_01144_, _01140_, _01107_);
  and (_01145_, _01144_, _01143_);
  not (_01146_, _33753_);
  and (_01147_, _01140_, _01124_);
  and (_01148_, _01147_, _01146_);
  or (_01149_, _01148_, _01145_);
  or (_01150_, _01149_, _01142_);
  not (_01151_, _33527_);
  and (_01152_, _01107_, _01101_);
  and (_01153_, _01152_, _01151_);
  not (_01154_, _33970_);
  and (_01155_, _01097_, _01093_);
  and (_01156_, _01155_, _01085_);
  and (_01157_, _01156_, _01154_);
  not (_01158_, _33609_);
  and (_01159_, _01155_, _01086_);
  and (_01160_, _01159_, _01158_);
  or (_01161_, _01160_, _01157_);
  not (_01162_, _33445_);
  and (_01163_, _01086_, _01099_);
  and (_01164_, _01163_, _01162_);
  not (_01165_, _33806_);
  and (_01166_, _01085_, _01099_);
  and (_01167_, _01166_, _01165_);
  or (_01168_, _01167_, _01164_);
  or (_01169_, _01168_, _01161_);
  or (_01170_, _01169_, _01153_);
  or (_01171_, _01170_, _01150_);
  or (_01172_, _01171_, _01138_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01172_, _01122_);
  and (_01173_, _01104_, _01127_);
  and (_01174_, _01125_, _01081_);
  or (_01175_, _01174_, _01173_);
  and (_01176_, _01111_, _01154_);
  and (_01177_, _01128_, _01131_);
  or (_01178_, _01177_, _01176_);
  or (_01179_, _01178_, _01175_);
  and (_01180_, _01119_, _01146_);
  and (_01181_, _01116_, _01165_);
  or (_01182_, _01181_, _01180_);
  and (_01183_, _01152_, _01162_);
  and (_01184_, _01135_, _01118_);
  or (_01185_, _01184_, _01183_);
  or (_01186_, _01185_, _01182_);
  and (_01187_, _01144_, _01158_);
  and (_01188_, _01141_, _01123_);
  and (_01189_, _01147_, _01139_);
  or (_01190_, _01189_, _01188_);
  or (_01191_, _01190_, _01187_);
  and (_01192_, _01132_, _01134_);
  and (_01193_, _01166_, _01143_);
  and (_01194_, _01156_, _01114_);
  or (_01195_, _01194_, _01193_);
  and (_01196_, _01163_, _01106_);
  and (_01197_, _01159_, _01151_);
  or (_01198_, _01197_, _01196_);
  or (_01199_, _01198_, _01195_);
  or (_01200_, _01199_, _01192_);
  or (_01201_, _01200_, _01191_);
  or (_01202_, _01201_, _01186_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01202_, _01179_);
  and (_01203_, _01116_, _01118_);
  and (_01204_, _01119_, _01165_);
  or (_01205_, _01204_, _01203_);
  and (_01206_, _01152_, _01081_);
  and (_01207_, _01104_, _01162_);
  or (_01208_, _01207_, _01206_);
  or (_01209_, _01208_, _01205_);
  and (_01210_, _01111_, _01131_);
  and (_01211_, _01128_, _01106_);
  or (_01212_, _01211_, _01210_);
  and (_01213_, _01132_, _01154_);
  and (_01214_, _01125_, _01151_);
  or (_01215_, _01214_, _01213_);
  or (_01216_, _01215_, _01212_);
  and (_01217_, _01141_, _01158_);
  and (_01218_, _01144_, _01139_);
  or (_01219_, _01218_, _01217_);
  and (_01220_, _01147_, _01143_);
  or (_01221_, _01220_, _01219_);
  and (_01222_, _01135_, _01114_);
  and (_01223_, _01166_, _01146_);
  and (_01224_, _01156_, _01134_);
  or (_01225_, _01224_, _01223_);
  and (_01226_, _01163_, _01127_);
  and (_01227_, _01159_, _01123_);
  or (_01228_, _01227_, _01226_);
  or (_01229_, _01228_, _01225_);
  or (_01230_, _01229_, _01222_);
  or (_01231_, _01230_, _01221_);
  or (_01232_, _01231_, _01216_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01232_, _01209_);
  and (_01233_, _01116_, _01146_);
  and (_01234_, _01111_, _01134_);
  or (_01235_, _01234_, _01233_);
  and (_01236_, _01152_, _01127_);
  and (_01237_, _01135_, _01165_);
  or (_01238_, _01237_, _01236_);
  or (_01239_, _01238_, _01235_);
  and (_01240_, _01125_, _01162_);
  and (_01241_, _01132_, _01114_);
  or (_01242_, _01241_, _01240_);
  and (_01243_, _01128_, _01154_);
  and (_01244_, _01119_, _01143_);
  or (_01245_, _01244_, _01243_);
  or (_01246_, _01245_, _01242_);
  and (_01247_, _01144_, _01123_);
  and (_01248_, _01141_, _01151_);
  or (_01249_, _01248_, _01247_);
  and (_01250_, _01147_, _01158_);
  or (_01251_, _01250_, _01249_);
  and (_01252_, _01104_, _01106_);
  and (_01253_, _01163_, _01131_);
  and (_01254_, _01156_, _01118_);
  or (_01255_, _01254_, _01253_);
  and (_01256_, _01159_, _01081_);
  and (_01257_, _01166_, _01139_);
  or (_01258_, _01257_, _01256_);
  or (_01259_, _01258_, _01255_);
  or (_01260_, _01259_, _01252_);
  or (_01261_, _01260_, _01251_);
  or (_01262_, _01261_, _01246_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01262_, _01239_);
  not (_01263_, _33308_);
  and (_01264_, _01132_, _01263_);
  not (_01265_, _33407_);
  and (_01266_, _01128_, _01265_);
  or (_01267_, _01266_, _01264_);
  not (_01268_, _33573_);
  and (_01269_, _01125_, _01268_);
  not (_01270_, _33491_);
  and (_01271_, _01104_, _01270_);
  or (_01272_, _01271_, _01269_);
  or (_01273_, _01272_, _01267_);
  not (_01274_, _33893_);
  and (_01275_, _01116_, _01274_);
  not (_01276_, _33852_);
  and (_01277_, _01119_, _01276_);
  or (_01278_, _01277_, _01275_);
  not (_01279_, _33366_);
  and (_01280_, _01111_, _01279_);
  not (_01281_, _33532_);
  and (_01282_, _01152_, _01281_);
  or (_01283_, _01282_, _01280_);
  or (_01284_, _01283_, _01278_);
  not (_01285_, _33760_);
  and (_01286_, _01147_, _01285_);
  not (_01287_, _33704_);
  and (_01288_, _01144_, _01287_);
  or (_01289_, _01288_, _01286_);
  not (_01290_, _33655_);
  and (_01291_, _01141_, _01290_);
  or (_01292_, _01291_, _01289_);
  not (_01293_, _33934_);
  and (_01294_, _01135_, _01293_);
  not (_01295_, _33975_);
  and (_01296_, _01156_, _01295_);
  not (_01297_, _33811_);
  and (_01298_, _01166_, _01297_);
  or (_01299_, _01298_, _01296_);
  not (_01300_, _33614_);
  and (_01301_, _01159_, _01300_);
  not (_01302_, _33450_);
  and (_01303_, _01163_, _01302_);
  or (_01304_, _01303_, _01301_);
  or (_01305_, _01304_, _01299_);
  or (_01306_, _01305_, _01294_);
  or (_01307_, _01306_, _01292_);
  or (_01308_, _01307_, _01284_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01308_, _01273_);
  not (_01309_, _33496_);
  and (_01310_, _01104_, _01309_);
  not (_01311_, _33412_);
  and (_01312_, _01128_, _01311_);
  or (_01313_, _01312_, _01310_);
  not (_01314_, _33578_);
  and (_01315_, _01125_, _01314_);
  not (_01316_, _33319_);
  and (_01317_, _01132_, _01316_);
  or (_01318_, _01317_, _01315_);
  or (_01319_, _01318_, _01313_);
  not (_01320_, _33939_);
  and (_01321_, _01135_, _01320_);
  not (_01322_, _33857_);
  and (_01323_, _01119_, _01322_);
  or (_01324_, _01323_, _01321_);
  not (_01325_, _33898_);
  and (_01326_, _01116_, _01325_);
  not (_01327_, _33371_);
  and (_01328_, _01111_, _01327_);
  or (_01329_, _01328_, _01326_);
  or (_01330_, _01329_, _01324_);
  not (_01331_, _33710_);
  and (_01332_, _01144_, _01331_);
  not (_01333_, _33766_);
  and (_01334_, _01147_, _01333_);
  or (_01335_, _01334_, _01332_);
  not (_01336_, _33660_);
  and (_01337_, _01141_, _01336_);
  or (_01338_, _01337_, _01335_);
  not (_01339_, _33537_);
  and (_01340_, _01152_, _01339_);
  not (_01341_, _33980_);
  and (_01342_, _01156_, _01341_);
  not (_01343_, _33455_);
  and (_01344_, _01163_, _01343_);
  or (_01345_, _01344_, _01342_);
  not (_01346_, _33816_);
  and (_01347_, _01166_, _01346_);
  not (_01348_, _33619_);
  and (_01349_, _01159_, _01348_);
  or (_01350_, _01349_, _01347_);
  or (_01351_, _01350_, _01345_);
  or (_01352_, _01351_, _01340_);
  or (_01353_, _01352_, _01338_);
  or (_01354_, _01353_, _01330_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01354_, _01319_);
  not (_01355_, _33583_);
  and (_01356_, _01125_, _01355_);
  not (_01357_, _33501_);
  and (_01358_, _01104_, _01357_);
  or (_01359_, _01358_, _01356_);
  not (_01360_, _33944_);
  and (_01361_, _01135_, _01360_);
  not (_01362_, _33418_);
  and (_01363_, _01128_, _01362_);
  or (_01364_, _01363_, _01361_);
  or (_01365_, _01364_, _01359_);
  not (_01366_, _33330_);
  and (_01367_, _01132_, _01366_);
  not (_01368_, _33376_);
  and (_01369_, _01111_, _01368_);
  or (_01370_, _01369_, _01367_);
  not (_01371_, _33903_);
  and (_01372_, _01116_, _01371_);
  not (_01373_, _33862_);
  and (_01374_, _01119_, _01373_);
  or (_01375_, _01374_, _01372_);
  or (_01376_, _01375_, _01370_);
  not (_01377_, _33773_);
  and (_01378_, _01147_, _01377_);
  not (_01379_, _33717_);
  and (_01380_, _01144_, _01379_);
  or (_01381_, _01380_, _01378_);
  not (_01382_, _33665_);
  and (_01383_, _01141_, _01382_);
  or (_01384_, _01383_, _01381_);
  not (_01385_, _33542_);
  and (_01386_, _01152_, _01385_);
  not (_01387_, _33821_);
  and (_01388_, _01166_, _01387_);
  not (_01389_, _33460_);
  and (_01390_, _01163_, _01389_);
  or (_01391_, _01390_, _01388_);
  not (_01392_, _33985_);
  and (_01393_, _01156_, _01392_);
  not (_01394_, _33624_);
  and (_01395_, _01159_, _01394_);
  or (_01396_, _01395_, _01393_);
  or (_01397_, _01396_, _01391_);
  or (_01398_, _01397_, _01386_);
  or (_01399_, _01398_, _01384_);
  or (_01400_, _01399_, _01376_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01400_, _01365_);
  not (_01401_, _33547_);
  and (_01402_, _01152_, _01401_);
  not (_01403_, _33381_);
  and (_01404_, _01111_, _01403_);
  or (_01405_, _01404_, _01402_);
  not (_01406_, _33423_);
  and (_01407_, _01128_, _01406_);
  not (_01408_, _33949_);
  and (_01409_, _01135_, _01408_);
  or (_01410_, _01409_, _01407_);
  or (_01411_, _01410_, _01405_);
  not (_01412_, _33506_);
  and (_01413_, _01104_, _01412_);
  not (_01414_, _33867_);
  and (_01415_, _01119_, _01414_);
  or (_01416_, _01415_, _01413_);
  not (_01417_, _33588_);
  and (_01418_, _01125_, _01417_);
  not (_01419_, _33340_);
  and (_01420_, _01132_, _01419_);
  or (_01421_, _01420_, _01418_);
  or (_01422_, _01421_, _01416_);
  not (_01423_, _33724_);
  and (_01424_, _01144_, _01423_);
  not (_01425_, _33780_);
  and (_01426_, _01147_, _01425_);
  not (_01427_, _33671_);
  and (_01428_, _01141_, _01427_);
  or (_01429_, _01428_, _01426_);
  or (_01430_, _01429_, _01424_);
  not (_01431_, _33908_);
  and (_01432_, _01116_, _01431_);
  not (_01433_, _33990_);
  and (_01434_, _01156_, _01433_);
  not (_01435_, _33826_);
  and (_01436_, _01166_, _01435_);
  or (_01437_, _01436_, _01434_);
  not (_01438_, _33465_);
  and (_01439_, _01163_, _01438_);
  not (_01440_, _33629_);
  and (_01441_, _01159_, _01440_);
  or (_01442_, _01441_, _01439_);
  or (_01443_, _01442_, _01437_);
  or (_01444_, _01443_, _01432_);
  or (_01445_, _01444_, _01430_);
  or (_01446_, _01445_, _01422_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01446_, _01411_);
  not (_01447_, _33913_);
  and (_01448_, _01116_, _01447_);
  not (_01449_, _33552_);
  and (_01450_, _01152_, _01449_);
  or (_01451_, _01450_, _01448_);
  not (_01452_, _33593_);
  and (_01453_, _01125_, _01452_);
  not (_01454_, _33345_);
  and (_01455_, _01132_, _01454_);
  or (_01456_, _01455_, _01453_);
  or (_01457_, _01456_, _01451_);
  not (_01458_, _33954_);
  and (_01459_, _01135_, _01458_);
  not (_01460_, _33872_);
  and (_01461_, _01119_, _01460_);
  or (_01462_, _01461_, _01459_);
  not (_01463_, _33511_);
  and (_01464_, _01104_, _01463_);
  not (_01465_, _33429_);
  and (_01466_, _01128_, _01465_);
  or (_01467_, _01466_, _01464_);
  or (_01468_, _01467_, _01462_);
  not (_01469_, _33732_);
  and (_01470_, _01144_, _01469_);
  not (_01471_, _33787_);
  and (_01472_, _01147_, _01471_);
  or (_01473_, _01472_, _01470_);
  not (_01474_, _33678_);
  and (_01475_, _01141_, _01474_);
  or (_01476_, _01475_, _01473_);
  not (_01477_, _33386_);
  and (_01478_, _01111_, _01477_);
  not (_01479_, _33831_);
  and (_01480_, _01166_, _01479_);
  not (_01481_, _33634_);
  and (_01482_, _01159_, _01481_);
  or (_01483_, _01482_, _01480_);
  not (_01484_, _33995_);
  and (_01485_, _01156_, _01484_);
  not (_01486_, _33470_);
  and (_01487_, _01163_, _01486_);
  or (_01488_, _01487_, _01485_);
  or (_01489_, _01488_, _01483_);
  or (_01490_, _01489_, _01478_);
  or (_01491_, _01490_, _01476_);
  or (_01492_, _01491_, _01468_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01492_, _01457_);
  not (_01493_, _33516_);
  and (_01494_, _01104_, _01493_);
  not (_01495_, _33434_);
  and (_01496_, _01128_, _01495_);
  or (_01497_, _01496_, _01494_);
  not (_01498_, _33350_);
  and (_01499_, _01132_, _01498_);
  not (_01500_, _33959_);
  and (_01501_, _01135_, _01500_);
  or (_01502_, _01501_, _01499_);
  or (_01503_, _01502_, _01497_);
  not (_01504_, _33598_);
  and (_01505_, _01125_, _01504_);
  not (_01506_, _33877_);
  and (_01507_, _01119_, _01506_);
  or (_01508_, _01507_, _01505_);
  not (_01509_, _33557_);
  and (_01510_, _01152_, _01509_);
  not (_01511_, _33391_);
  and (_01512_, _01111_, _01511_);
  or (_01513_, _01512_, _01510_);
  or (_01514_, _01513_, _01508_);
  not (_01515_, _33684_);
  and (_01516_, _01141_, _01515_);
  not (_01517_, _33737_);
  and (_01518_, _01144_, _01517_);
  not (_01519_, _33794_);
  and (_01520_, _01147_, _01519_);
  or (_01521_, _01520_, _01518_);
  or (_01522_, _01521_, _01516_);
  not (_01523_, _33918_);
  and (_01524_, _01116_, _01523_);
  not (_01525_, _34000_);
  and (_01526_, _01156_, _01525_);
  not (_01527_, _33836_);
  and (_01528_, _01166_, _01527_);
  or (_01529_, _01528_, _01526_);
  not (_01530_, _33475_);
  and (_01531_, _01163_, _01530_);
  not (_01532_, _33639_);
  and (_01533_, _01159_, _01532_);
  or (_01534_, _01533_, _01531_);
  or (_01535_, _01534_, _01529_);
  or (_01536_, _01535_, _01524_);
  or (_01537_, _01536_, _01522_);
  or (_01538_, _01537_, _01514_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01538_, _01503_);
  not (_01539_, _33355_);
  and (_01540_, _01132_, _01539_);
  not (_01541_, _33439_);
  and (_01542_, _01128_, _01541_);
  or (_01543_, _01542_, _01540_);
  not (_01544_, _33603_);
  and (_01545_, _01125_, _01544_);
  not (_01546_, _33521_);
  and (_01547_, _01104_, _01546_);
  or (_01548_, _01547_, _01545_);
  or (_01549_, _01548_, _01543_);
  not (_01550_, _33923_);
  and (_01551_, _01116_, _01550_);
  not (_01552_, _33882_);
  and (_01553_, _01119_, _01552_);
  or (_01554_, _01553_, _01551_);
  not (_01555_, _33396_);
  and (_01556_, _01111_, _01555_);
  not (_01557_, _33562_);
  and (_01558_, _01152_, _01557_);
  or (_01559_, _01558_, _01556_);
  or (_01560_, _01559_, _01554_);
  not (_01561_, _33800_);
  and (_01562_, _01147_, _01561_);
  not (_01563_, _33744_);
  and (_01564_, _01144_, _01563_);
  or (_01565_, _01564_, _01562_);
  not (_01566_, _33690_);
  and (_01567_, _01141_, _01566_);
  or (_01568_, _01567_, _01565_);
  not (_01569_, _33964_);
  and (_01570_, _01135_, _01569_);
  not (_01571_, _34005_);
  and (_01572_, _01156_, _01571_);
  not (_01573_, _33841_);
  and (_01574_, _01166_, _01573_);
  or (_01575_, _01574_, _01572_);
  not (_01576_, _33644_);
  and (_01577_, _01159_, _01576_);
  not (_01578_, _33480_);
  and (_01579_, _01163_, _01578_);
  or (_01580_, _01579_, _01577_);
  or (_01581_, _01580_, _01575_);
  or (_01582_, _01581_, _01570_);
  or (_01583_, _01582_, _01568_);
  or (_01584_, _01583_, _01560_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01584_, _01549_);
  and (_01585_, _01132_, _01293_);
  and (_01586_, _01135_, _01276_);
  or (_01587_, _01586_, _01585_);
  and (_01588_, _01152_, _01302_);
  and (_01589_, _01104_, _01265_);
  or (_01590_, _01589_, _01588_);
  or (_01591_, _01590_, _01587_);
  and (_01592_, _01128_, _01263_);
  and (_01593_, _01116_, _01297_);
  or (_01594_, _01593_, _01592_);
  and (_01595_, _01111_, _01295_);
  and (_01596_, _01119_, _01285_);
  or (_01597_, _01596_, _01595_);
  or (_01598_, _01597_, _01594_);
  and (_01599_, _01147_, _01290_);
  and (_01600_, _01141_, _01268_);
  and (_01601_, _01144_, _01300_);
  or (_01602_, _01601_, _01600_);
  or (_01603_, _01602_, _01599_);
  and (_01604_, _01125_, _01270_);
  and (_01605_, _01159_, _01281_);
  and (_01606_, _01156_, _01274_);
  or (_01607_, _01606_, _01605_);
  and (_01608_, _01163_, _01279_);
  and (_01609_, _01166_, _01287_);
  or (_01610_, _01609_, _01608_);
  or (_01611_, _01610_, _01607_);
  or (_01612_, _01611_, _01604_);
  or (_01613_, _01612_, _01603_);
  or (_01614_, _01613_, _01598_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01614_, _01591_);
  and (_01615_, _01111_, _01341_);
  and (_01616_, _01116_, _01346_);
  or (_01617_, _01616_, _01615_);
  and (_01618_, _01125_, _01309_);
  and (_01619_, _01135_, _01322_);
  or (_01620_, _01619_, _01618_);
  or (_01621_, _01620_, _01617_);
  and (_01622_, _01152_, _01343_);
  and (_01623_, _01132_, _01320_);
  or (_01624_, _01623_, _01622_);
  and (_01625_, _01104_, _01311_);
  and (_01626_, _01119_, _01333_);
  or (_01627_, _01626_, _01625_);
  or (_01628_, _01627_, _01624_);
  and (_01629_, _01144_, _01348_);
  and (_01630_, _01141_, _01314_);
  and (_01631_, _01147_, _01336_);
  or (_01632_, _01631_, _01630_);
  or (_01633_, _01632_, _01629_);
  and (_01634_, _01128_, _01316_);
  and (_01635_, _01163_, _01327_);
  and (_01636_, _01156_, _01325_);
  or (_01637_, _01636_, _01635_);
  and (_01638_, _01159_, _01339_);
  and (_01639_, _01166_, _01331_);
  or (_01640_, _01639_, _01638_);
  or (_01641_, _01640_, _01637_);
  or (_01642_, _01641_, _01634_);
  or (_01643_, _01642_, _01633_);
  or (_01644_, _01643_, _01628_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01644_, _01621_);
  and (_01645_, _01132_, _01360_);
  and (_01646_, _01135_, _01373_);
  or (_01647_, _01646_, _01645_);
  and (_01648_, _01111_, _01392_);
  and (_01649_, _01128_, _01366_);
  or (_01650_, _01649_, _01648_);
  or (_01651_, _01650_, _01647_);
  and (_01652_, _01119_, _01377_);
  and (_01653_, _01116_, _01387_);
  or (_01654_, _01653_, _01652_);
  and (_01655_, _01125_, _01357_);
  and (_01656_, _01104_, _01362_);
  or (_01657_, _01656_, _01655_);
  or (_01658_, _01657_, _01654_);
  and (_01659_, _01147_, _01382_);
  and (_01660_, _01141_, _01355_);
  and (_01661_, _01144_, _01394_);
  or (_01662_, _01661_, _01660_);
  or (_01663_, _01662_, _01659_);
  and (_01664_, _01152_, _01389_);
  and (_01665_, _01166_, _01379_);
  and (_01666_, _01156_, _01371_);
  or (_01667_, _01666_, _01665_);
  and (_01668_, _01159_, _01385_);
  and (_01669_, _01163_, _01368_);
  or (_01670_, _01669_, _01668_);
  or (_01671_, _01670_, _01667_);
  or (_01672_, _01671_, _01664_);
  or (_01673_, _01672_, _01663_);
  or (_01674_, _01673_, _01658_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01674_, _01651_);
  and (_01675_, _01104_, _01406_);
  and (_01676_, _01125_, _01412_);
  or (_01677_, _01676_, _01675_);
  and (_01678_, _01111_, _01433_);
  and (_01679_, _01128_, _01419_);
  or (_01680_, _01679_, _01678_);
  or (_01681_, _01680_, _01677_);
  and (_01682_, _01119_, _01425_);
  and (_01683_, _01116_, _01435_);
  or (_01684_, _01683_, _01682_);
  and (_01685_, _01152_, _01438_);
  and (_01686_, _01135_, _01414_);
  or (_01687_, _01686_, _01685_);
  or (_01688_, _01687_, _01684_);
  and (_01689_, _01144_, _01440_);
  and (_01690_, _01141_, _01417_);
  and (_01691_, _01147_, _01427_);
  or (_01692_, _01691_, _01690_);
  or (_01693_, _01692_, _01689_);
  and (_01694_, _01132_, _01408_);
  and (_01695_, _01166_, _01423_);
  and (_01696_, _01156_, _01431_);
  or (_01697_, _01696_, _01695_);
  and (_01698_, _01163_, _01403_);
  and (_01699_, _01159_, _01401_);
  or (_01700_, _01699_, _01698_);
  or (_01701_, _01700_, _01697_);
  or (_01702_, _01701_, _01694_);
  or (_01703_, _01702_, _01693_);
  or (_01704_, _01703_, _01688_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _01704_, _01681_);
  and (_01705_, _01132_, _01458_);
  and (_01706_, _01116_, _01479_);
  or (_01707_, _01706_, _01705_);
  and (_01708_, _01111_, _01484_);
  and (_01709_, _01128_, _01454_);
  or (_01710_, _01709_, _01708_);
  or (_01711_, _01710_, _01707_);
  and (_01712_, _01119_, _01471_);
  and (_01713_, _01135_, _01460_);
  or (_01714_, _01713_, _01712_);
  and (_01715_, _01125_, _01463_);
  and (_01716_, _01104_, _01465_);
  or (_01717_, _01716_, _01715_);
  or (_01718_, _01717_, _01714_);
  and (_01719_, _01147_, _01474_);
  and (_01720_, _01141_, _01452_);
  and (_01721_, _01144_, _01481_);
  or (_01722_, _01721_, _01720_);
  or (_01723_, _01722_, _01719_);
  and (_01724_, _01152_, _01486_);
  and (_01725_, _01166_, _01469_);
  and (_01726_, _01156_, _01447_);
  or (_01727_, _01726_, _01725_);
  and (_01728_, _01159_, _01449_);
  and (_01729_, _01163_, _01477_);
  or (_01730_, _01729_, _01728_);
  or (_01731_, _01730_, _01727_);
  or (_01732_, _01731_, _01724_);
  or (_01733_, _01732_, _01723_);
  or (_01734_, _01733_, _01718_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _01734_, _01711_);
  and (_01735_, _01104_, _01495_);
  and (_01736_, _01116_, _01527_);
  or (_01737_, _01736_, _01735_);
  and (_01738_, _01128_, _01498_);
  and (_01739_, _01132_, _01500_);
  or (_01740_, _01739_, _01738_);
  or (_01741_, _01740_, _01737_);
  and (_01742_, _01125_, _01493_);
  and (_01743_, _01152_, _01530_);
  or (_01744_, _01743_, _01742_);
  and (_01745_, _01111_, _01525_);
  and (_01746_, _01119_, _01519_);
  or (_01747_, _01746_, _01745_);
  or (_01748_, _01747_, _01744_);
  and (_01749_, _01147_, _01515_);
  and (_01750_, _01141_, _01504_);
  and (_01751_, _01144_, _01532_);
  or (_01752_, _01751_, _01750_);
  or (_01753_, _01752_, _01749_);
  and (_01754_, _01135_, _01506_);
  and (_01755_, _01163_, _01511_);
  and (_01756_, _01156_, _01523_);
  or (_01757_, _01756_, _01755_);
  and (_01758_, _01159_, _01509_);
  and (_01759_, _01166_, _01517_);
  or (_01760_, _01759_, _01758_);
  or (_01761_, _01760_, _01757_);
  or (_01762_, _01761_, _01754_);
  or (_01763_, _01762_, _01753_);
  or (_01764_, _01763_, _01748_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _01764_, _01741_);
  and (_01765_, _01104_, _01541_);
  and (_01766_, _01116_, _01573_);
  or (_01767_, _01766_, _01765_);
  and (_01768_, _01125_, _01546_);
  and (_01769_, _01135_, _01552_);
  or (_01770_, _01769_, _01768_);
  or (_01771_, _01770_, _01767_);
  and (_01772_, _01128_, _01539_);
  and (_01773_, _01119_, _01561_);
  or (_01774_, _01773_, _01772_);
  and (_01775_, _01111_, _01571_);
  and (_01776_, _01152_, _01578_);
  or (_01777_, _01776_, _01775_);
  or (_01778_, _01777_, _01774_);
  and (_01779_, _01144_, _01576_);
  and (_01780_, _01141_, _01544_);
  and (_01781_, _01147_, _01566_);
  or (_01782_, _01781_, _01780_);
  or (_01783_, _01782_, _01779_);
  and (_01784_, _01132_, _01569_);
  and (_01785_, _01166_, _01563_);
  and (_01786_, _01156_, _01550_);
  or (_01787_, _01786_, _01785_);
  and (_01788_, _01163_, _01555_);
  and (_01789_, _01159_, _01557_);
  or (_01790_, _01789_, _01788_);
  or (_01791_, _01790_, _01787_);
  or (_01792_, _01791_, _01784_);
  or (_01793_, _01792_, _01783_);
  or (_01794_, _01793_, _01778_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _01794_, _01771_);
  and (_01795_, _01116_, _01276_);
  and (_01796_, _01119_, _01297_);
  or (_01797_, _01796_, _01795_);
  and (_01798_, _01132_, _01295_);
  and (_01799_, _01125_, _01281_);
  or (_01800_, _01799_, _01798_);
  or (_01801_, _01800_, _01797_);
  and (_01802_, _01111_, _01263_);
  and (_01803_, _01128_, _01279_);
  or (_01804_, _01803_, _01802_);
  and (_01805_, _01135_, _01274_);
  and (_01806_, _01104_, _01302_);
  or (_01807_, _01806_, _01805_);
  or (_01808_, _01807_, _01804_);
  and (_01809_, _01144_, _01290_);
  and (_01810_, _01147_, _01287_);
  and (_01811_, _01141_, _01300_);
  or (_01812_, _01811_, _01810_);
  or (_01813_, _01812_, _01809_);
  and (_01814_, _01152_, _01270_);
  and (_01815_, _01166_, _01285_);
  and (_01816_, _01156_, _01293_);
  or (_01817_, _01816_, _01815_);
  and (_01818_, _01163_, _01265_);
  and (_01819_, _01159_, _01268_);
  or (_01820_, _01819_, _01818_);
  or (_01821_, _01820_, _01817_);
  or (_01822_, _01821_, _01814_);
  or (_01823_, _01822_, _01813_);
  or (_01824_, _01823_, _01808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _01824_, _01801_);
  and (_01825_, _01119_, _01346_);
  and (_01826_, _01152_, _01309_);
  or (_01827_, _01826_, _01825_);
  and (_01828_, _01104_, _01343_);
  and (_01829_, _01111_, _01316_);
  or (_01830_, _01829_, _01828_);
  or (_01831_, _01830_, _01827_);
  and (_01832_, _01132_, _01341_);
  and (_01833_, _01116_, _01322_);
  or (_01834_, _01833_, _01832_);
  and (_01835_, _01135_, _01325_);
  and (_01836_, _01128_, _01327_);
  or (_01837_, _01836_, _01835_);
  or (_01838_, _01837_, _01834_);
  and (_01839_, _01141_, _01348_);
  and (_01840_, _01147_, _01331_);
  and (_01841_, _01144_, _01336_);
  or (_01842_, _01841_, _01840_);
  or (_01843_, _01842_, _01839_);
  and (_01844_, _01125_, _01339_);
  and (_01845_, _01156_, _01320_);
  and (_01846_, _01159_, _01314_);
  or (_01847_, _01846_, _01845_);
  and (_01848_, _01166_, _01333_);
  and (_01849_, _01163_, _01311_);
  or (_01850_, _01849_, _01848_);
  or (_01851_, _01850_, _01847_);
  or (_01852_, _01851_, _01844_);
  or (_01853_, _01852_, _01843_);
  or (_01854_, _01853_, _01838_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _01854_, _01831_);
  and (_01855_, _01119_, _01387_);
  and (_01856_, _01128_, _01368_);
  or (_01857_, _01856_, _01855_);
  and (_01858_, _01104_, _01389_);
  and (_01859_, _01111_, _01366_);
  or (_01860_, _01859_, _01858_);
  or (_01861_, _01860_, _01857_);
  and (_01862_, _01132_, _01392_);
  and (_01863_, _01116_, _01373_);
  or (_01864_, _01863_, _01862_);
  and (_01865_, _01135_, _01371_);
  and (_01866_, _01152_, _01357_);
  or (_01867_, _01866_, _01865_);
  or (_01868_, _01867_, _01864_);
  and (_01869_, _01141_, _01394_);
  and (_01870_, _01147_, _01379_);
  and (_01871_, _01144_, _01382_);
  or (_01872_, _01871_, _01870_);
  or (_01873_, _01872_, _01869_);
  and (_01874_, _01125_, _01385_);
  and (_01875_, _01156_, _01360_);
  and (_01876_, _01159_, _01355_);
  or (_01877_, _01876_, _01875_);
  and (_01878_, _01166_, _01377_);
  and (_01879_, _01163_, _01362_);
  or (_01880_, _01879_, _01878_);
  or (_01881_, _01880_, _01877_);
  or (_01882_, _01881_, _01874_);
  or (_01883_, _01882_, _01873_);
  or (_01884_, _01883_, _01868_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _01884_, _01861_);
  and (_01885_, _01111_, _01419_);
  and (_01886_, _01104_, _01438_);
  or (_01887_, _01886_, _01885_);
  and (_01888_, _01135_, _01431_);
  and (_01889_, _01116_, _01414_);
  or (_01890_, _01889_, _01888_);
  or (_01891_, _01890_, _01887_);
  and (_01892_, _01132_, _01433_);
  and (_01893_, _01128_, _01403_);
  or (_01894_, _01893_, _01892_);
  and (_01895_, _01125_, _01401_);
  and (_01896_, _01152_, _01412_);
  or (_01897_, _01896_, _01895_);
  or (_01898_, _01897_, _01894_);
  and (_01899_, _01144_, _01427_);
  and (_01900_, _01141_, _01440_);
  or (_01901_, _01900_, _01899_);
  and (_01902_, _01147_, _01423_);
  or (_01903_, _01902_, _01901_);
  and (_01904_, _01119_, _01435_);
  and (_01905_, _01163_, _01406_);
  and (_01906_, _01156_, _01408_);
  or (_01907_, _01906_, _01905_);
  and (_01908_, _01159_, _01417_);
  and (_01909_, _01166_, _01425_);
  or (_01910_, _01909_, _01908_);
  or (_01911_, _01910_, _01907_);
  or (_01912_, _01911_, _01904_);
  or (_01913_, _01912_, _01903_);
  or (_01914_, _01913_, _01898_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _01914_, _01891_);
  and (_01915_, _01128_, _01477_);
  and (_01916_, _01152_, _01463_);
  or (_01917_, _01916_, _01915_);
  and (_01918_, _01135_, _01447_);
  and (_01919_, _01104_, _01486_);
  or (_01920_, _01919_, _01918_);
  or (_01921_, _01920_, _01917_);
  and (_01922_, _01119_, _01479_);
  and (_01923_, _01111_, _01454_);
  or (_01924_, _01923_, _01922_);
  and (_01925_, _01116_, _01460_);
  and (_01926_, _01125_, _01449_);
  or (_01927_, _01926_, _01925_);
  or (_01928_, _01927_, _01924_);
  and (_01929_, _01144_, _01474_);
  and (_01930_, _01141_, _01481_);
  or (_01931_, _01930_, _01929_);
  and (_01932_, _01147_, _01469_);
  or (_01933_, _01932_, _01931_);
  and (_01934_, _01132_, _01484_);
  and (_01935_, _01156_, _01458_);
  and (_01936_, _01163_, _01465_);
  or (_01937_, _01936_, _01935_);
  and (_01938_, _01166_, _01471_);
  and (_01939_, _01159_, _01452_);
  or (_01940_, _01939_, _01938_);
  or (_01941_, _01940_, _01937_);
  or (_01942_, _01941_, _01934_);
  or (_01943_, _01942_, _01933_);
  or (_01944_, _01943_, _01928_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _01944_, _01921_);
  and (_01945_, _01116_, _01506_);
  and (_01946_, _01119_, _01527_);
  or (_01947_, _01946_, _01945_);
  and (_01948_, _01132_, _01525_);
  and (_01949_, _01125_, _01509_);
  or (_01950_, _01949_, _01948_);
  or (_01951_, _01950_, _01947_);
  and (_01952_, _01111_, _01498_);
  and (_01953_, _01128_, _01511_);
  or (_01954_, _01953_, _01952_);
  and (_01955_, _01135_, _01523_);
  and (_01956_, _01104_, _01530_);
  or (_01957_, _01956_, _01955_);
  or (_01958_, _01957_, _01954_);
  and (_01959_, _01144_, _01515_);
  and (_01960_, _01147_, _01517_);
  and (_01961_, _01141_, _01532_);
  or (_01962_, _01961_, _01960_);
  or (_01963_, _01962_, _01959_);
  and (_01964_, _01152_, _01493_);
  and (_01965_, _01166_, _01519_);
  and (_01966_, _01156_, _01500_);
  or (_01967_, _01966_, _01965_);
  and (_01968_, _01163_, _01495_);
  and (_01969_, _01159_, _01504_);
  or (_01970_, _01969_, _01968_);
  or (_01971_, _01970_, _01967_);
  or (_01972_, _01971_, _01964_);
  or (_01973_, _01972_, _01963_);
  or (_01974_, _01973_, _01958_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _01974_, _01951_);
  and (_01975_, _01125_, _01557_);
  and (_01976_, _01128_, _01555_);
  or (_01977_, _01976_, _01975_);
  and (_01978_, _01132_, _01571_);
  and (_01979_, _01111_, _01539_);
  or (_01980_, _01979_, _01978_);
  or (_01981_, _01980_, _01977_);
  and (_01982_, _01104_, _01578_);
  and (_01983_, _01152_, _01546_);
  or (_01984_, _01983_, _01982_);
  and (_01985_, _01119_, _01573_);
  and (_01986_, _01116_, _01552_);
  or (_01987_, _01986_, _01985_);
  or (_01988_, _01987_, _01984_);
  and (_01989_, _01144_, _01566_);
  and (_01990_, _01147_, _01563_);
  and (_01991_, _01141_, _01576_);
  or (_01992_, _01991_, _01990_);
  or (_01993_, _01992_, _01989_);
  and (_01994_, _01135_, _01550_);
  and (_01995_, _01166_, _01561_);
  and (_01996_, _01156_, _01569_);
  or (_01997_, _01996_, _01995_);
  and (_01998_, _01159_, _01544_);
  and (_01999_, _01163_, _01541_);
  or (_02000_, _01999_, _01998_);
  or (_02001_, _02000_, _01997_);
  or (_02002_, _02001_, _01994_);
  or (_02003_, _02002_, _01993_);
  or (_02004_, _02003_, _01988_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02004_, _01981_);
  and (_02005_, _01152_, _01265_);
  and (_02006_, _01116_, _01285_);
  or (_02007_, _02006_, _02005_);
  and (_02008_, _01119_, _01287_);
  and (_02009_, _01111_, _01293_);
  or (_02010_, _02009_, _02008_);
  or (_02011_, _02010_, _02007_);
  and (_02012_, _01125_, _01302_);
  and (_02013_, _01135_, _01297_);
  or (_02014_, _02013_, _02012_);
  and (_02015_, _01104_, _01279_);
  and (_02016_, _01132_, _01274_);
  or (_02017_, _02016_, _02015_);
  or (_02018_, _02017_, _02014_);
  and (_02019_, _01141_, _01281_);
  and (_02020_, _01144_, _01268_);
  or (_02021_, _02020_, _02019_);
  and (_02022_, _01147_, _01300_);
  or (_02023_, _02022_, _02021_);
  and (_02024_, _01128_, _01295_);
  and (_02025_, _01166_, _01290_);
  and (_02026_, _01156_, _01276_);
  or (_02027_, _02026_, _02025_);
  and (_02028_, _01159_, _01270_);
  and (_02029_, _01163_, _01263_);
  or (_02030_, _02029_, _02028_);
  or (_02031_, _02030_, _02027_);
  or (_02032_, _02031_, _02024_);
  or (_02033_, _02032_, _02023_);
  or (_02034_, _02033_, _02018_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02034_, _02011_);
  and (_02035_, _01119_, _01331_);
  and (_02036_, _01111_, _01320_);
  or (_02037_, _02036_, _02035_);
  and (_02038_, _01152_, _01311_);
  and (_02039_, _01135_, _01346_);
  or (_02040_, _02039_, _02038_);
  or (_02041_, _02040_, _02037_);
  and (_02042_, _01125_, _01343_);
  and (_02043_, _01132_, _01325_);
  or (_02044_, _02043_, _02042_);
  and (_02045_, _01128_, _01341_);
  and (_02046_, _01116_, _01333_);
  or (_02047_, _02046_, _02045_);
  or (_02048_, _02047_, _02044_);
  and (_02049_, _01144_, _01314_);
  and (_02050_, _01141_, _01339_);
  or (_02051_, _02050_, _02049_);
  and (_02052_, _01147_, _01348_);
  or (_02053_, _02052_, _02051_);
  and (_02054_, _01104_, _01327_);
  and (_02055_, _01163_, _01316_);
  and (_02056_, _01156_, _01322_);
  or (_02057_, _02056_, _02055_);
  and (_02058_, _01159_, _01309_);
  and (_02059_, _01166_, _01336_);
  or (_02060_, _02059_, _02058_);
  or (_02061_, _02060_, _02057_);
  or (_02062_, _02061_, _02054_);
  or (_02063_, _02062_, _02053_);
  or (_02064_, _02063_, _02048_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02064_, _02041_);
  and (_02065_, _01116_, _01377_);
  and (_02066_, _01111_, _01360_);
  or (_02067_, _02066_, _02065_);
  and (_02068_, _01152_, _01362_);
  and (_02069_, _01135_, _01387_);
  or (_02070_, _02069_, _02068_);
  or (_02071_, _02070_, _02067_);
  and (_02072_, _01125_, _01389_);
  and (_02073_, _01132_, _01371_);
  or (_02074_, _02073_, _02072_);
  and (_02075_, _01128_, _01392_);
  and (_02076_, _01119_, _01379_);
  or (_02077_, _02076_, _02075_);
  or (_02078_, _02077_, _02074_);
  and (_02079_, _01144_, _01355_);
  and (_02080_, _01141_, _01385_);
  or (_02081_, _02080_, _02079_);
  and (_02082_, _01147_, _01394_);
  or (_02083_, _02082_, _02081_);
  and (_02084_, _01104_, _01368_);
  and (_02085_, _01163_, _01366_);
  and (_02086_, _01156_, _01373_);
  or (_02087_, _02086_, _02085_);
  and (_02088_, _01159_, _01357_);
  and (_02089_, _01166_, _01382_);
  or (_02090_, _02089_, _02088_);
  or (_02091_, _02090_, _02087_);
  or (_02092_, _02091_, _02084_);
  or (_02093_, _02092_, _02083_);
  or (_02094_, _02093_, _02078_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02094_, _02071_);
  and (_02095_, _01152_, _01406_);
  and (_02096_, _01119_, _01423_);
  or (_02097_, _02096_, _02095_);
  and (_02098_, _01116_, _01425_);
  and (_02099_, _01111_, _01408_);
  or (_02100_, _02099_, _02098_);
  or (_02101_, _02100_, _02097_);
  and (_02102_, _01128_, _01433_);
  and (_02103_, _01125_, _01438_);
  or (_02104_, _02103_, _02102_);
  and (_02105_, _01104_, _01403_);
  and (_02106_, _01132_, _01431_);
  or (_02107_, _02106_, _02105_);
  or (_02108_, _02107_, _02104_);
  and (_02109_, _01144_, _01417_);
  and (_02110_, _01141_, _01401_);
  and (_02111_, _01147_, _01440_);
  or (_02112_, _02111_, _02110_);
  or (_02113_, _02112_, _02109_);
  and (_02114_, _01135_, _01435_);
  and (_02115_, _01159_, _01412_);
  and (_02116_, _01156_, _01414_);
  or (_02117_, _02116_, _02115_);
  and (_02118_, _01163_, _01419_);
  and (_02119_, _01166_, _01427_);
  or (_02120_, _02119_, _02118_);
  or (_02121_, _02120_, _02117_);
  or (_02122_, _02121_, _02114_);
  or (_02123_, _02122_, _02113_);
  or (_02124_, _02123_, _02108_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02124_, _02101_);
  and (_02125_, _01125_, _01486_);
  and (_02126_, _01132_, _01447_);
  or (_02127_, _02126_, _02125_);
  and (_02128_, _01128_, _01484_);
  and (_02129_, _01152_, _01465_);
  or (_02130_, _02129_, _02128_);
  or (_02131_, _02130_, _02127_);
  and (_02132_, _01116_, _01471_);
  and (_02133_, _01135_, _01479_);
  or (_02134_, _02133_, _02132_);
  and (_02135_, _01104_, _01477_);
  and (_02136_, _01119_, _01469_);
  or (_02137_, _02136_, _02135_);
  or (_02138_, _02137_, _02134_);
  and (_02139_, _01141_, _01449_);
  and (_02140_, _01144_, _01452_);
  and (_02141_, _01147_, _01481_);
  or (_02142_, _02141_, _02140_);
  or (_02143_, _02142_, _02139_);
  and (_02144_, _01111_, _01458_);
  and (_02145_, _01166_, _01474_);
  and (_02146_, _01156_, _01460_);
  or (_02147_, _02146_, _02145_);
  and (_02148_, _01159_, _01463_);
  and (_02149_, _01163_, _01454_);
  or (_02150_, _02149_, _02148_);
  or (_02151_, _02150_, _02147_);
  or (_02152_, _02151_, _02144_);
  or (_02153_, _02152_, _02143_);
  or (_02154_, _02153_, _02138_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02154_, _02131_);
  and (_02155_, _01116_, _01519_);
  and (_02156_, _01132_, _01523_);
  or (_02157_, _02156_, _02155_);
  and (_02158_, _01125_, _01530_);
  and (_02159_, _01135_, _01527_);
  or (_02160_, _02159_, _02158_);
  or (_02161_, _02160_, _02157_);
  and (_02162_, _01152_, _01495_);
  and (_02163_, _01119_, _01517_);
  or (_02164_, _02163_, _02162_);
  and (_02165_, _01128_, _01525_);
  and (_02166_, _01104_, _01511_);
  or (_02167_, _02166_, _02165_);
  or (_02168_, _02167_, _02164_);
  and (_02169_, _01141_, _01509_);
  and (_02170_, _01144_, _01504_);
  and (_02171_, _01147_, _01532_);
  or (_02172_, _02171_, _02170_);
  or (_02173_, _02172_, _02169_);
  and (_02174_, _01111_, _01500_);
  and (_02175_, _01166_, _01515_);
  and (_02176_, _01156_, _01506_);
  or (_02177_, _02176_, _02175_);
  and (_02178_, _01159_, _01493_);
  and (_02179_, _01163_, _01498_);
  or (_02180_, _02179_, _02178_);
  or (_02181_, _02180_, _02177_);
  or (_02182_, _02181_, _02174_);
  or (_02183_, _02182_, _02173_);
  or (_02184_, _02183_, _02168_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02184_, _02161_);
  and (_02185_, _01125_, _01578_);
  and (_02186_, _01132_, _01550_);
  or (_02187_, _02186_, _02185_);
  and (_02188_, _01128_, _01571_);
  and (_02189_, _01152_, _01541_);
  or (_02190_, _02189_, _02188_);
  or (_02191_, _02190_, _02187_);
  and (_02192_, _01116_, _01561_);
  and (_02193_, _01135_, _01573_);
  or (_02194_, _02193_, _02192_);
  and (_02195_, _01104_, _01555_);
  and (_02196_, _01119_, _01563_);
  or (_02197_, _02196_, _02195_);
  or (_02198_, _02197_, _02194_);
  and (_02199_, _01141_, _01557_);
  and (_02200_, _01144_, _01544_);
  and (_02201_, _01147_, _01576_);
  or (_02202_, _02201_, _02200_);
  or (_02203_, _02202_, _02199_);
  and (_02204_, _01111_, _01569_);
  and (_02205_, _01166_, _01566_);
  and (_02206_, _01156_, _01552_);
  or (_02207_, _02206_, _02205_);
  and (_02208_, _01159_, _01546_);
  and (_02209_, _01163_, _01539_);
  or (_02210_, _02209_, _02208_);
  or (_02211_, _02210_, _02207_);
  or (_02212_, _02211_, _02204_);
  or (_02213_, _02212_, _02203_);
  or (_02214_, _02213_, _02198_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02214_, _02191_);
  nand (_02215_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02216_, \oc8051_golden_model_1.PC [3]);
  or (_02217_, \oc8051_golden_model_1.PC [2], _02216_);
  or (_02218_, _02217_, _02215_);
  or (_02219_, _02218_, _33821_);
  not (_02220_, \oc8051_golden_model_1.PC [1]);
  or (_02221_, _02220_, \oc8051_golden_model_1.PC [0]);
  or (_02222_, _02221_, _02217_);
  or (_02223_, _02222_, _33773_);
  and (_02224_, _02223_, _02219_);
  not (_02225_, \oc8051_golden_model_1.PC [2]);
  or (_02226_, _02225_, \oc8051_golden_model_1.PC [3]);
  or (_02227_, _02226_, _02215_);
  or (_02228_, _02227_, _33624_);
  or (_02229_, _02226_, _02221_);
  or (_02230_, _02229_, _33583_);
  and (_02231_, _02230_, _02228_);
  and (_02232_, _02231_, _02224_);
  nand (_02233_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02234_, _02233_, _02215_);
  or (_02235_, _02234_, _33985_);
  or (_02236_, _02233_, _02221_);
  or (_02237_, _02236_, _33944_);
  and (_02238_, _02237_, _02235_);
  or (_02239_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02240_, _02239_, _02215_);
  or (_02241_, _02240_, _33460_);
  or (_02242_, _02239_, _02221_);
  or (_02243_, _02242_, _33418_);
  and (_02244_, _02243_, _02241_);
  and (_02245_, _02244_, _02238_);
  and (_02246_, _02245_, _02232_);
  not (_02247_, \oc8051_golden_model_1.PC [0]);
  or (_02248_, \oc8051_golden_model_1.PC [1], _02247_);
  or (_02249_, _02248_, _02233_);
  or (_02250_, _02249_, _33903_);
  or (_02251_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02252_, _02251_, _02233_);
  or (_02253_, _02252_, _33862_);
  and (_02254_, _02253_, _02250_);
  or (_02255_, _02239_, _02251_);
  or (_02256_, _02255_, _33330_);
  or (_02257_, _02239_, _02248_);
  or (_02258_, _02257_, _33376_);
  and (_02259_, _02258_, _02256_);
  and (_02260_, _02259_, _02254_);
  or (_02261_, _02248_, _02217_);
  or (_02262_, _02261_, _33717_);
  or (_02263_, _02251_, _02217_);
  or (_02264_, _02263_, _33665_);
  and (_02265_, _02264_, _02262_);
  or (_02266_, _02248_, _02226_);
  or (_02267_, _02266_, _33542_);
  or (_02268_, _02251_, _02226_);
  or (_02269_, _02268_, _33501_);
  and (_02270_, _02269_, _02267_);
  and (_02271_, _02270_, _02265_);
  and (_02272_, _02271_, _02260_);
  nand (_02273_, _02272_, _02246_);
  or (_02274_, _02218_, _33826_);
  or (_02275_, _02222_, _33780_);
  and (_02276_, _02275_, _02274_);
  or (_02277_, _02227_, _33629_);
  or (_02278_, _02229_, _33588_);
  and (_02279_, _02278_, _02277_);
  and (_02280_, _02279_, _02276_);
  or (_02281_, _02234_, _33990_);
  or (_02282_, _02236_, _33949_);
  and (_02283_, _02282_, _02281_);
  or (_02284_, _02240_, _33465_);
  or (_02285_, _02242_, _33423_);
  and (_02286_, _02285_, _02284_);
  and (_02287_, _02286_, _02283_);
  and (_02288_, _02287_, _02280_);
  or (_02289_, _02249_, _33908_);
  or (_02290_, _02252_, _33867_);
  and (_02291_, _02290_, _02289_);
  or (_02292_, _02255_, _33340_);
  or (_02293_, _02257_, _33381_);
  and (_02294_, _02293_, _02292_);
  and (_02295_, _02294_, _02291_);
  or (_02296_, _02261_, _33724_);
  or (_02297_, _02263_, _33671_);
  and (_02298_, _02297_, _02296_);
  or (_02299_, _02266_, _33547_);
  or (_02300_, _02268_, _33506_);
  and (_02301_, _02300_, _02299_);
  and (_02302_, _02301_, _02298_);
  and (_02303_, _02302_, _02295_);
  nand (_02304_, _02303_, _02288_);
  or (_02305_, _02304_, _02273_);
  or (_02306_, _02218_, _33811_);
  or (_02307_, _02222_, _33760_);
  and (_02308_, _02307_, _02306_);
  or (_02309_, _02227_, _33614_);
  or (_02310_, _02229_, _33573_);
  and (_02311_, _02310_, _02309_);
  and (_02312_, _02311_, _02308_);
  or (_02313_, _02234_, _33975_);
  or (_02314_, _02236_, _33934_);
  and (_02315_, _02314_, _02313_);
  or (_02316_, _02240_, _33450_);
  or (_02317_, _02242_, _33407_);
  and (_02318_, _02317_, _02316_);
  and (_02319_, _02318_, _02315_);
  and (_02320_, _02319_, _02312_);
  or (_02321_, _02249_, _33893_);
  or (_02322_, _02252_, _33852_);
  and (_02323_, _02322_, _02321_);
  or (_02324_, _02255_, _33308_);
  or (_02325_, _02257_, _33366_);
  and (_02326_, _02325_, _02324_);
  and (_02327_, _02326_, _02323_);
  or (_02328_, _02261_, _33704_);
  or (_02329_, _02263_, _33655_);
  and (_02330_, _02329_, _02328_);
  or (_02331_, _02266_, _33532_);
  or (_02332_, _02268_, _33491_);
  and (_02333_, _02332_, _02331_);
  and (_02334_, _02333_, _02330_);
  and (_02335_, _02334_, _02327_);
  and (_02336_, _02335_, _02320_);
  or (_02337_, _02218_, _33816_);
  or (_02338_, _02222_, _33766_);
  and (_02339_, _02338_, _02337_);
  or (_02340_, _02227_, _33619_);
  or (_02341_, _02229_, _33578_);
  and (_02342_, _02341_, _02340_);
  and (_02343_, _02342_, _02339_);
  or (_02344_, _02234_, _33980_);
  or (_02345_, _02236_, _33939_);
  and (_02346_, _02345_, _02344_);
  or (_02347_, _02240_, _33455_);
  or (_02348_, _02242_, _33412_);
  and (_02349_, _02348_, _02347_);
  and (_02350_, _02349_, _02346_);
  and (_02351_, _02350_, _02343_);
  or (_02352_, _02249_, _33898_);
  or (_02353_, _02252_, _33857_);
  and (_02354_, _02353_, _02352_);
  or (_02355_, _02255_, _33319_);
  or (_02356_, _02257_, _33371_);
  and (_02357_, _02356_, _02355_);
  and (_02358_, _02357_, _02354_);
  or (_02359_, _02261_, _33710_);
  or (_02360_, _02263_, _33660_);
  and (_02361_, _02360_, _02359_);
  or (_02362_, _02266_, _33537_);
  or (_02363_, _02268_, _33496_);
  and (_02364_, _02363_, _02362_);
  and (_02365_, _02364_, _02361_);
  and (_02366_, _02365_, _02358_);
  nand (_02367_, _02366_, _02351_);
  or (_02368_, _02367_, _02336_);
  or (_02369_, _02368_, _02305_);
  not (_02370_, _02369_);
  or (_02371_, _02218_, _33841_);
  or (_02372_, _02222_, _33800_);
  and (_02373_, _02372_, _02371_);
  or (_02374_, _02227_, _33644_);
  or (_02375_, _02229_, _33603_);
  and (_02376_, _02375_, _02374_);
  and (_02377_, _02376_, _02373_);
  or (_02378_, _02234_, _34005_);
  or (_02379_, _02236_, _33964_);
  and (_02380_, _02379_, _02378_);
  or (_02381_, _02240_, _33480_);
  or (_02382_, _02242_, _33439_);
  and (_02383_, _02382_, _02381_);
  and (_02384_, _02383_, _02380_);
  and (_02385_, _02384_, _02377_);
  or (_02386_, _02249_, _33923_);
  or (_02387_, _02252_, _33882_);
  and (_02388_, _02387_, _02386_);
  or (_02389_, _02255_, _33355_);
  or (_02390_, _02257_, _33396_);
  and (_02391_, _02390_, _02389_);
  and (_02392_, _02391_, _02388_);
  or (_02393_, _02261_, _33744_);
  or (_02394_, _02263_, _33690_);
  and (_02395_, _02394_, _02393_);
  or (_02396_, _02266_, _33562_);
  or (_02397_, _02268_, _33521_);
  and (_02398_, _02397_, _02396_);
  and (_02399_, _02398_, _02395_);
  and (_02400_, _02399_, _02392_);
  and (_02401_, _02400_, _02385_);
  or (_02402_, _02218_, _33806_);
  or (_02403_, _02222_, _33753_);
  and (_02404_, _02403_, _02402_);
  or (_02405_, _02227_, _33609_);
  or (_02406_, _02229_, _33568_);
  and (_02407_, _02406_, _02405_);
  and (_02408_, _02407_, _02404_);
  or (_02409_, _02234_, _33970_);
  or (_02410_, _02236_, _33929_);
  and (_02411_, _02410_, _02409_);
  or (_02412_, _02240_, _33445_);
  or (_02413_, _02242_, _33402_);
  and (_02414_, _02413_, _02412_);
  and (_02415_, _02414_, _02411_);
  and (_02416_, _02415_, _02408_);
  or (_02417_, _02249_, _33888_);
  or (_02418_, _02252_, _33847_);
  and (_02419_, _02418_, _02417_);
  or (_02420_, _02255_, _33297_);
  or (_02421_, _02257_, _33361_);
  and (_02422_, _02421_, _02420_);
  and (_02423_, _02422_, _02419_);
  or (_02424_, _02261_, _33697_);
  or (_02425_, _02263_, _33650_);
  and (_02426_, _02425_, _02424_);
  or (_02427_, _02266_, _33527_);
  or (_02428_, _02268_, _33486_);
  and (_02429_, _02428_, _02427_);
  and (_02430_, _02429_, _02426_);
  and (_02431_, _02430_, _02423_);
  and (_02432_, _02431_, _02416_);
  and (_02433_, _02432_, _02401_);
  or (_02434_, _02218_, _33831_);
  or (_02435_, _02222_, _33787_);
  and (_02436_, _02435_, _02434_);
  or (_02437_, _02227_, _33634_);
  or (_02438_, _02229_, _33593_);
  and (_02439_, _02438_, _02437_);
  and (_02440_, _02439_, _02436_);
  or (_02441_, _02234_, _33995_);
  or (_02442_, _02236_, _33954_);
  and (_02443_, _02442_, _02441_);
  or (_02444_, _02240_, _33470_);
  or (_02445_, _02242_, _33429_);
  and (_02446_, _02445_, _02444_);
  and (_02447_, _02446_, _02443_);
  and (_02448_, _02447_, _02440_);
  or (_02449_, _02249_, _33913_);
  or (_02450_, _02252_, _33872_);
  and (_02451_, _02450_, _02449_);
  or (_02452_, _02255_, _33345_);
  or (_02453_, _02257_, _33386_);
  and (_02454_, _02453_, _02452_);
  and (_02455_, _02454_, _02451_);
  or (_02456_, _02261_, _33732_);
  or (_02457_, _02263_, _33678_);
  and (_02458_, _02457_, _02456_);
  or (_02459_, _02266_, _33552_);
  or (_02460_, _02268_, _33511_);
  and (_02461_, _02460_, _02459_);
  and (_02462_, _02461_, _02458_);
  and (_02463_, _02462_, _02455_);
  nand (_02464_, _02463_, _02448_);
  or (_02465_, _02218_, _33836_);
  or (_02466_, _02222_, _33794_);
  and (_02467_, _02466_, _02465_);
  or (_02468_, _02227_, _33639_);
  or (_02469_, _02229_, _33598_);
  and (_02470_, _02469_, _02468_);
  and (_02471_, _02470_, _02467_);
  or (_02472_, _02234_, _34000_);
  or (_02473_, _02236_, _33959_);
  and (_02474_, _02473_, _02472_);
  or (_02475_, _02240_, _33475_);
  or (_02476_, _02242_, _33434_);
  and (_02477_, _02476_, _02475_);
  and (_02478_, _02477_, _02474_);
  and (_02479_, _02478_, _02471_);
  or (_02480_, _02249_, _33918_);
  or (_02481_, _02252_, _33877_);
  and (_02482_, _02481_, _02480_);
  or (_02483_, _02255_, _33350_);
  or (_02484_, _02257_, _33391_);
  and (_02485_, _02484_, _02483_);
  and (_02486_, _02485_, _02482_);
  or (_02487_, _02261_, _33737_);
  or (_02488_, _02263_, _33684_);
  and (_02489_, _02488_, _02487_);
  or (_02490_, _02266_, _33557_);
  or (_02491_, _02268_, _33516_);
  and (_02492_, _02491_, _02490_);
  and (_02493_, _02492_, _02489_);
  and (_02494_, _02493_, _02486_);
  nand (_02495_, _02494_, _02479_);
  or (_02496_, _02495_, _02464_);
  not (_02497_, _02496_);
  and (_02498_, _02497_, _02433_);
  and (_02499_, _02498_, _02370_);
  not (_02500_, _02499_);
  and (_02501_, _02463_, _02448_);
  or (_02502_, _02495_, _02501_);
  not (_02503_, _02502_);
  and (_02504_, _02503_, _02433_);
  and (_02505_, _02504_, _02370_);
  and (_02506_, _02494_, _02479_);
  or (_02507_, _02506_, _02464_);
  not (_02508_, _02507_);
  and (_02509_, _02508_, _02433_);
  and (_02510_, _02509_, _02370_);
  nor (_02511_, _02510_, _02505_);
  and (_02512_, _02511_, _02500_);
  nand (_02513_, _02400_, _02385_);
  or (_02514_, _02432_, _02513_);
  nor (_02515_, _02514_, _02496_);
  and (_02516_, _02515_, _02370_);
  not (_02517_, _02516_);
  or (_02518_, _02506_, _02501_);
  not (_02519_, _02518_);
  and (_02520_, _02432_, _02513_);
  and (_02521_, _02520_, _02519_);
  and (_02522_, _02521_, _02370_);
  and (_02523_, _02508_, _02520_);
  and (_02524_, _02523_, _02370_);
  nor (_02525_, _02524_, _02522_);
  and (_02526_, _02525_, _02517_);
  and (_02527_, _02433_, _02519_);
  and (_02528_, _02527_, _02370_);
  and (_02529_, _02503_, _02520_);
  and (_02530_, _02529_, _02370_);
  nor (_02531_, _02530_, _02528_);
  and (_02532_, _02497_, _02520_);
  and (_02533_, _02532_, _02370_);
  not (_02534_, _02533_);
  and (_02535_, _02534_, _02531_);
  and (_02536_, _02535_, _02526_);
  and (_02537_, _02536_, _02512_);
  and (_02538_, _02366_, _02351_);
  or (_02539_, _02538_, _02336_);
  or (_02540_, _02539_, _02305_);
  not (_02541_, _02540_);
  and (_02542_, _02541_, _02515_);
  not (_02543_, \oc8051_golden_model_1.ACC [1]);
  and (_02544_, _02248_, _02221_);
  nor (_02545_, _02544_, _02543_);
  and (_02546_, \oc8051_golden_model_1.ACC [0], _02247_);
  and (_02547_, _02544_, _02543_);
  nor (_02548_, _02547_, _02545_);
  and (_02549_, _02548_, _02546_);
  nor (_02550_, _02549_, _02545_);
  nor (_02551_, _02215_, _02225_);
  and (_02552_, _02215_, _02225_);
  nor (_02553_, _02552_, _02551_);
  and (_02554_, _02553_, \oc8051_golden_model_1.ACC [2]);
  nor (_02555_, _02553_, \oc8051_golden_model_1.ACC [2]);
  nor (_02557_, _02555_, _02554_);
  not (_02558_, _02557_);
  and (_02559_, _02558_, _02550_);
  nor (_02560_, _02558_, _02550_);
  nor (_02561_, _02560_, _02559_);
  and (_02562_, _02561_, _02542_);
  not (_02563_, _02368_);
  not (_02564_, _02304_);
  and (_02565_, _02564_, _02273_);
  and (_02566_, _02565_, _02563_);
  and (_02567_, _02566_, _02515_);
  or (_02568_, _02514_, _02502_);
  nor (_02569_, _02568_, _02369_);
  nor (_02570_, _02569_, _02567_);
  or (_02571_, _02568_, _02540_);
  and (_02572_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_02573_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02574_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_02575_, _02574_, _02572_);
  and (_02576_, _02575_, _02573_);
  nor (_02577_, _02576_, _02572_);
  and (_02578_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02579_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02580_, _02579_, _02578_);
  not (_02581_, _02580_);
  nor (_02582_, _02581_, _02577_);
  and (_02583_, _02581_, _02577_);
  nor (_02584_, _02583_, _02582_);
  not (_02585_, _02584_);
  or (_02586_, _02585_, _02571_);
  and (_02587_, _02586_, _02570_);
  or (_02588_, _02514_, _02507_);
  or (_02589_, _02588_, _02369_);
  or (_02590_, _02514_, _02518_);
  or (_02591_, _02590_, _02369_);
  and (_02592_, _02591_, _02589_);
  or (_02593_, _02432_, _02401_);
  or (_02594_, _02593_, _02496_);
  or (_02595_, _02594_, _02369_);
  or (_02596_, _02593_, _02502_);
  or (_02597_, _02596_, _02369_);
  and (_02598_, _02597_, _02595_);
  and (_02599_, _02598_, _02592_);
  or (_02600_, _02593_, _02507_);
  or (_02601_, _02600_, _02369_);
  or (_02602_, _02593_, _02518_);
  or (_02603_, _02602_, _02369_);
  and (_02604_, _02603_, _02601_);
  nand (_02605_, _02604_, _02599_);
  or (_02606_, _02553_, _02605_);
  nand (_02607_, _02606_, _02571_);
  nand (_02608_, _02607_, _02587_);
  not (_02609_, _02542_);
  and (_02610_, _02604_, _02599_);
  and (_02611_, _02610_, _02570_);
  and (_02612_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02613_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02614_, _02613_, _02612_);
  or (_02615_, _02614_, _02611_);
  and (_02616_, _02615_, _02609_);
  and (_02617_, _02616_, _02608_);
  or (_02618_, _02617_, _02562_);
  nand (_02619_, _02618_, _02537_);
  not (_02620_, _02614_);
  nor (_02621_, _02620_, _02537_);
  not (_02622_, _02621_);
  and (_02623_, _02622_, _02619_);
  nor (_02624_, _02560_, _02554_);
  not (_02625_, \oc8051_golden_model_1.ACC [3]);
  not (_02626_, _02227_);
  nor (_02627_, _02551_, _02216_);
  nor (_02628_, _02627_, _02626_);
  nor (_02629_, _02628_, _02625_);
  and (_02630_, _02628_, _02625_);
  nor (_02631_, _02630_, _02629_);
  nor (_02632_, _02631_, _02624_);
  and (_02633_, _02631_, _02624_);
  or (_02634_, _02633_, _02632_);
  and (_02635_, _02634_, _02542_);
  not (_02636_, _02628_);
  or (_02637_, _02605_, _02636_);
  nor (_02638_, _02233_, _02220_);
  nor (_02639_, _02612_, \oc8051_golden_model_1.PC [3]);
  nor (_02640_, _02639_, _02638_);
  or (_02641_, _02640_, _02610_);
  and (_02642_, _02641_, _02637_);
  nand (_02643_, _02642_, _02571_);
  nor (_02644_, _02582_, _02578_);
  and (_02645_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02646_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02647_, _02646_, _02645_);
  not (_02648_, _02647_);
  nor (_02649_, _02648_, _02644_);
  and (_02650_, _02648_, _02644_);
  nor (_02651_, _02650_, _02649_);
  not (_02652_, _02651_);
  or (_02653_, _02652_, _02571_);
  and (_02654_, _02653_, _02570_);
  nand (_02655_, _02654_, _02643_);
  or (_02656_, _02640_, _02570_);
  and (_02657_, _02656_, _02609_);
  and (_02658_, _02657_, _02655_);
  or (_02659_, _02658_, _02635_);
  and (_02660_, _02659_, _02537_);
  not (_02661_, _02640_);
  nor (_02662_, _02661_, _02537_);
  or (_02663_, _02662_, _02660_);
  or (_02664_, _02663_, _02623_);
  nor (_02665_, _02537_, _02220_);
  not (_02666_, _02665_);
  nor (_02667_, _02548_, _02546_);
  nor (_02668_, _02667_, _02549_);
  and (_02669_, _02668_, _02542_);
  and (_02670_, _02571_, _02544_);
  and (_02671_, _02670_, _02604_);
  nand (_02672_, _02671_, _02599_);
  nor (_02673_, _02575_, _02573_);
  nor (_02674_, _02673_, _02576_);
  or (_02675_, _02674_, _02571_);
  nand (_02676_, _02675_, _02672_);
  nand (_02677_, _02676_, _02570_);
  or (_02678_, _02611_, _02220_);
  and (_02679_, _02678_, _02677_);
  and (_02680_, _02679_, _02609_);
  nor (_02681_, _02680_, _02669_);
  nand (_02682_, _02681_, _02537_);
  and (_02683_, _02682_, _02666_);
  or (_02684_, _02605_, _02247_);
  or (_02685_, _02610_, \oc8051_golden_model_1.PC [0]);
  nand (_02686_, _02685_, _02684_);
  nand (_02687_, _02686_, _02571_);
  nor (_02688_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02689_, _02688_, _02573_);
  or (_02690_, _02689_, _02571_);
  and (_02691_, _02690_, _02570_);
  and (_02692_, _02691_, _02687_);
  nor (_02693_, _02570_, _02247_);
  or (_02694_, _02693_, _02692_);
  nand (_02695_, _02694_, _02609_);
  not (_02696_, \oc8051_golden_model_1.ACC [0]);
  and (_02697_, _02696_, \oc8051_golden_model_1.PC [0]);
  or (_02698_, _02546_, _02609_);
  or (_02699_, _02698_, _02697_);
  and (_02700_, _02699_, _02537_);
  nand (_02701_, _02700_, _02695_);
  nor (_02702_, _02537_, \oc8051_golden_model_1.PC [0]);
  not (_02703_, _02702_);
  and (_02704_, _02703_, _02701_);
  or (_02705_, _02704_, _02683_);
  or (_02706_, _02705_, _02664_);
  or (_02707_, _02706_, _33486_);
  nand (_02708_, _02682_, _02666_);
  or (_02709_, _02704_, _02708_);
  nand (_02710_, _02622_, _02619_);
  or (_02711_, _02663_, _02710_);
  or (_02712_, _02711_, _02709_);
  or (_02713_, _02712_, _33402_);
  and (_02714_, _02713_, _02707_);
  nand (_02715_, _02703_, _02701_);
  or (_02716_, _02715_, _02683_);
  nor (_02717_, _02662_, _02660_);
  or (_02718_, _02717_, _02623_);
  or (_02719_, _02718_, _02716_);
  or (_02720_, _02719_, _33888_);
  or (_02721_, _02717_, _02710_);
  or (_02722_, _02721_, _02716_);
  or (_02723_, _02722_, _33697_);
  and (_02724_, _02723_, _02720_);
  and (_02725_, _02724_, _02714_);
  or (_02726_, _02664_, _02709_);
  or (_02727_, _02726_, _33568_);
  or (_02728_, _02716_, _02664_);
  or (_02729_, _02728_, _33527_);
  and (_02730_, _02729_, _02727_);
  or (_02731_, _02705_, _02711_);
  or (_02732_, _02731_, _33297_);
  or (_02733_, _02711_, _02716_);
  or (_02734_, _02733_, _33361_);
  and (_02735_, _02734_, _02732_);
  and (_02736_, _02735_, _02730_);
  and (_02737_, _02736_, _02725_);
  or (_02738_, _02718_, _02705_);
  or (_02739_, _02738_, _33847_);
  or (_02740_, _02715_, _02708_);
  or (_02741_, _02721_, _02740_);
  or (_02742_, _02741_, _33806_);
  and (_02743_, _02742_, _02739_);
  or (_02744_, _02718_, _02740_);
  or (_02745_, _02744_, _33970_);
  or (_02746_, _02718_, _02709_);
  or (_02747_, _02746_, _33929_);
  and (_02748_, _02747_, _02745_);
  and (_02749_, _02748_, _02743_);
  or (_02750_, _02740_, _02664_);
  or (_02751_, _02750_, _33609_);
  or (_02752_, _02711_, _02740_);
  or (_02753_, _02752_, _33445_);
  and (_02754_, _02753_, _02751_);
  or (_02755_, _02721_, _02709_);
  or (_02756_, _02755_, _33753_);
  or (_02758_, _02705_, _02721_);
  or (_02759_, _02758_, _33650_);
  and (_02760_, _02759_, _02756_);
  and (_02761_, _02760_, _02754_);
  and (_02762_, _02761_, _02749_);
  and (_02763_, _02762_, _02737_);
  or (_02764_, _02744_, _33990_);
  or (_02765_, _02706_, _33506_);
  and (_02766_, _02765_, _02764_);
  or (_02767_, _02755_, _33780_);
  or (_02768_, _02752_, _33465_);
  and (_02769_, _02768_, _02767_);
  and (_02770_, _02769_, _02766_);
  or (_02771_, _02746_, _33949_);
  or (_02772_, _02719_, _33908_);
  and (_02773_, _02772_, _02771_);
  or (_02774_, _02750_, _33629_);
  or (_02775_, _02726_, _33588_);
  and (_02776_, _02775_, _02774_);
  and (_02777_, _02776_, _02773_);
  and (_02778_, _02777_, _02770_);
  or (_02779_, _02728_, _33547_);
  or (_02780_, _02712_, _33423_);
  and (_02781_, _02780_, _02779_);
  or (_02782_, _02731_, _33340_);
  or (_02783_, _02733_, _33381_);
  and (_02784_, _02783_, _02782_);
  and (_02785_, _02784_, _02781_);
  or (_02786_, _02738_, _33867_);
  or (_02787_, _02758_, _33671_);
  and (_02788_, _02787_, _02786_);
  or (_02789_, _02741_, _33826_);
  or (_02790_, _02722_, _33724_);
  and (_02791_, _02790_, _02789_);
  and (_02792_, _02791_, _02788_);
  and (_02793_, _02792_, _02785_);
  nand (_02794_, _02793_, _02778_);
  and (_02795_, _02794_, _02763_);
  not (_02796_, _02305_);
  and (_02797_, _02538_, _02336_);
  and (_02798_, _02797_, _02796_);
  and (_02799_, _02798_, _02504_);
  and (_02800_, _02799_, _02795_);
  and (_02801_, _02799_, _02763_);
  not (_02802_, _02801_);
  or (_02803_, _02726_, _33573_);
  or (_02804_, _02728_, _33532_);
  and (_02805_, _02804_, _02803_);
  or (_02806_, _02752_, _33450_);
  or (_02807_, _02712_, _33407_);
  and (_02808_, _02807_, _02806_);
  and (_02809_, _02808_, _02805_);
  or (_02810_, _02722_, _33704_);
  or (_02811_, _02758_, _33655_);
  and (_02812_, _02811_, _02810_);
  or (_02813_, _02719_, _33893_);
  or (_02814_, _02738_, _33852_);
  and (_02815_, _02814_, _02813_);
  and (_02816_, _02815_, _02812_);
  and (_02817_, _02816_, _02809_);
  or (_02818_, _02731_, _33308_);
  or (_02819_, _02733_, _33366_);
  and (_02820_, _02819_, _02818_);
  or (_02821_, _02750_, _33614_);
  or (_02822_, _02706_, _33491_);
  and (_02823_, _02822_, _02821_);
  and (_02824_, _02823_, _02820_);
  or (_02825_, _02744_, _33975_);
  or (_02826_, _02746_, _33934_);
  and (_02827_, _02826_, _02825_);
  or (_02828_, _02741_, _33811_);
  or (_02829_, _02755_, _33760_);
  and (_02830_, _02829_, _02828_);
  and (_02831_, _02830_, _02827_);
  and (_02832_, _02831_, _02824_);
  nand (_02833_, _02832_, _02817_);
  and (_02834_, _02566_, _02521_);
  and (_02835_, _02834_, _02763_);
  and (_02836_, _02835_, _02833_);
  and (_02837_, _02832_, _02817_);
  not (_02838_, _02763_);
  not (_02839_, _02567_);
  and (_02840_, _02565_, _02367_);
  and (_02841_, _02840_, _02515_);
  not (_02842_, _02841_);
  not (_02843_, _02273_);
  and (_02844_, _02538_, _02304_);
  and (_02845_, _02844_, _02843_);
  and (_02846_, _02845_, _02515_);
  not (_02847_, _02846_);
  and (_02848_, _02367_, _02336_);
  and (_02849_, _02304_, _02843_);
  and (_02850_, _02849_, _02848_);
  and (_02851_, _02850_, _02515_);
  not (_02852_, _02515_);
  not (_02853_, _02539_);
  and (_02854_, _02849_, _02853_);
  and (_02855_, _02304_, _02273_);
  nor (_02856_, _02855_, _02854_);
  nor (_02857_, _02856_, _02852_);
  nor (_02858_, _02857_, _02851_);
  and (_02859_, _02858_, _02847_);
  and (_02860_, _02859_, _02842_);
  and (_02861_, _02860_, _02839_);
  nor (_02862_, _02861_, _02838_);
  and (_02863_, _02862_, _02837_);
  not (_02864_, _02568_);
  and (_02865_, _02848_, _02796_);
  and (_02866_, _02865_, _02864_);
  and (_02867_, _02795_, _02866_);
  not (_02868_, \oc8051_golden_model_1.SP [0]);
  nor (_02869_, _02591_, _02868_);
  not (_02870_, _02590_);
  and (_02871_, _02865_, _02870_);
  and (_02872_, _02871_, _02795_);
  and (_02873_, _02871_, _02763_);
  not (_02874_, _02873_);
  not (_02875_, _02594_);
  and (_02876_, _02798_, _02875_);
  and (_02877_, _02865_, _02875_);
  and (_02878_, _02877_, _02795_);
  and (_02879_, _02877_, _02763_);
  and (_02880_, _02875_, _02566_);
  and (_02881_, _02880_, _02763_);
  and (_02882_, _02881_, _02833_);
  not (_02883_, _02596_);
  and (_02884_, _02865_, _02883_);
  and (_02885_, _02884_, _02795_);
  and (_02886_, _02884_, _02763_);
  and (_02887_, _02566_, _02498_);
  not (_02888_, _02887_);
  and (_02889_, _02798_, _02509_);
  and (_02890_, _02865_, _02509_);
  not (_02891_, _02890_);
  and (_02892_, _02566_, _02509_);
  nor (_02893_, _02741_, _33841_);
  nor (_02894_, _02750_, _33644_);
  nor (_02895_, _02894_, _02893_);
  nor (_02896_, _02726_, _33603_);
  nor (_02897_, _02731_, _33355_);
  nor (_02898_, _02897_, _02896_);
  and (_02899_, _02898_, _02895_);
  nor (_02900_, _02744_, _34005_);
  nor (_02901_, _02752_, _33480_);
  nor (_02902_, _02901_, _02900_);
  nor (_02903_, _02746_, _33964_);
  nor (_02904_, _02758_, _33690_);
  nor (_02905_, _02904_, _02903_);
  and (_02906_, _02905_, _02902_);
  and (_02907_, _02906_, _02899_);
  nor (_02908_, _02728_, _33562_);
  nor (_02909_, _02706_, _33521_);
  nor (_02910_, _02909_, _02908_);
  nor (_02911_, _02755_, _33800_);
  nor (_02912_, _02733_, _33396_);
  nor (_02913_, _02912_, _02911_);
  and (_02914_, _02913_, _02910_);
  nor (_02915_, _02719_, _33923_);
  nor (_02916_, _02712_, _33439_);
  nor (_02917_, _02916_, _02915_);
  nor (_02919_, _02738_, _33882_);
  nor (_02920_, _02722_, _33744_);
  nor (_02921_, _02920_, _02919_);
  and (_02922_, _02921_, _02917_);
  and (_02923_, _02922_, _02914_);
  and (_02924_, _02923_, _02907_);
  nor (_02925_, _02924_, _02838_);
  and (_02926_, _02794_, _02838_);
  nor (_02927_, _02926_, _02925_);
  and (_02928_, _02865_, _02521_);
  and (_02930_, _02865_, _02515_);
  nor (_02931_, _02930_, _02928_);
  not (_02932_, _02931_);
  and (_02933_, _02932_, _02927_);
  not (_02934_, _02884_);
  nor (_02935_, _02877_, _02866_);
  and (_02936_, _02935_, _02934_);
  and (_02937_, _02798_, _02870_);
  nor (_02938_, _02871_, _02937_);
  not (_02939_, _02588_);
  and (_02940_, _02798_, _02939_);
  and (_02941_, _02865_, _02939_);
  nor (_02942_, _02941_, _02940_);
  and (_02943_, _02942_, _02938_);
  and (_02944_, _02943_, _02936_);
  nor (_02945_, _02944_, _02927_);
  and (_02946_, _02798_, _02883_);
  and (_02947_, _02946_, \oc8051_golden_model_1.SP [3]);
  and (_02948_, _02883_, _02566_);
  not (_02949_, _02600_);
  and (_02951_, _02949_, _02566_);
  nor (_02952_, _02951_, _02948_);
  nor (_02953_, _02952_, _02794_);
  and (_02954_, _02870_, _02566_);
  nor (_02955_, _02954_, _02876_);
  and (_02956_, _02849_, _02367_);
  and (_02957_, _02956_, _02939_);
  not (_02958_, _02957_);
  and (_02959_, _02849_, _02563_);
  and (_02960_, _02959_, _02939_);
  and (_02962_, _02849_, _02797_);
  and (_02963_, _02962_, _02939_);
  nor (_02964_, _02963_, _02960_);
  and (_02965_, _02964_, _02958_);
  and (_02966_, _02855_, _02538_);
  and (_02967_, _02966_, _02939_);
  and (_02968_, _02855_, _02367_);
  and (_02969_, _02968_, _02939_);
  nor (_02970_, _02969_, _02967_);
  and (_02971_, _02970_, _02965_);
  and (_02973_, _02971_, _02955_);
  not (_02974_, \oc8051_golden_model_1.PSW [3]);
  and (_02975_, _02952_, _02974_);
  nor (_02976_, _02946_, _02884_);
  not (_02977_, _02976_);
  or (_02978_, _02977_, _02975_);
  and (_02979_, _02864_, _02566_);
  nor (_02980_, _02979_, _02880_);
  and (_02981_, _02980_, _02978_);
  and (_02982_, _02981_, _02973_);
  nor (_02983_, _02982_, _02953_);
  or (_02984_, _02983_, _02947_);
  or (_02985_, _02984_, _02945_);
  not (_02986_, _02866_);
  not (_02987_, _02877_);
  and (_02988_, _02943_, _02987_);
  nand (_02989_, _02988_, _02986_);
  nand (_02990_, _02989_, _02927_);
  not (_02991_, _02979_);
  not (_02992_, _02880_);
  and (_02994_, _02955_, _02992_);
  and (_02995_, _02994_, _02971_);
  and (_02996_, _02995_, _02991_);
  or (_02997_, _02996_, _02794_);
  and (_02998_, _02997_, _02990_);
  and (_02999_, _02998_, _02985_);
  and (_03000_, _02999_, _02839_);
  and (_03001_, _02854_, _02870_);
  and (_03002_, _02855_, _02797_);
  and (_03003_, _03002_, _02870_);
  nor (_03005_, _03003_, _03001_);
  not (_03006_, _02948_);
  and (_03007_, _02855_, _02853_);
  and (_03008_, _03007_, _02870_);
  and (_03009_, _02855_, _02563_);
  and (_03010_, _03009_, _02870_);
  nor (_03011_, _03010_, _03008_);
  and (_03012_, _03011_, _03006_);
  and (_03013_, _03012_, _03005_);
  and (_03014_, _02565_, _02853_);
  and (_03016_, _03014_, _02870_);
  and (_03017_, _02962_, _02870_);
  or (_03018_, _03017_, _03016_);
  nor (_03019_, _02850_, _02959_);
  nor (_03020_, _03019_, _02590_);
  nor (_03021_, _03020_, _03018_);
  and (_03022_, _02541_, _02529_);
  not (_03023_, _03022_);
  and (_03024_, _02848_, _02565_);
  and (_03025_, _03024_, _02870_);
  not (_03027_, _03025_);
  and (_03028_, _02797_, _02565_);
  and (_03029_, _03028_, _02870_);
  nor (_03030_, _03029_, _02954_);
  and (_03031_, _03030_, _03027_);
  and (_03032_, _03031_, _03023_);
  and (_03033_, _03032_, _03021_);
  and (_03034_, _02865_, _02504_);
  nor (_03035_, _03034_, _02799_);
  and (_03036_, _02865_, _02498_);
  not (_03038_, _03036_);
  and (_03039_, _03038_, _03035_);
  and (_03040_, _02798_, _02527_);
  nor (_03041_, _02889_, _03040_);
  and (_03042_, _02541_, _02532_);
  not (_03043_, _03042_);
  and (_03044_, _03043_, _03041_);
  and (_03045_, _03044_, _03039_);
  and (_03046_, _02798_, _02864_);
  and (_03047_, _02855_, _02848_);
  and (_03049_, _03047_, _02870_);
  nor (_03050_, _03049_, _03046_);
  and (_03051_, _02541_, _02523_);
  nor (_03052_, _03051_, _02834_);
  and (_03053_, _03052_, _03050_);
  and (_03054_, _03053_, _03045_);
  and (_03055_, _03054_, _03033_);
  and (_03056_, _03055_, _03013_);
  and (_03057_, _03056_, _02553_);
  nor (_03058_, _03056_, _02620_);
  nor (_03060_, _03058_, _03057_);
  nor (_03061_, _03056_, _02661_);
  and (_03062_, _03056_, _02636_);
  nor (_03063_, _03062_, _03061_);
  nor (_03064_, _03063_, _03060_);
  nand (_03065_, _03056_, _02247_);
  or (_03066_, _03056_, _02247_);
  nand (_03067_, _03066_, _03065_);
  and (_03068_, _03065_, \oc8051_golden_model_1.PC [1]);
  nor (_03069_, _03065_, \oc8051_golden_model_1.PC [1]);
  nor (_03071_, _03069_, _03068_);
  and (_03072_, _03071_, _03067_);
  and (_03073_, _03072_, _03064_);
  and (_03074_, _03073_, _01433_);
  and (_03075_, _03063_, _03060_);
  and (_03076_, _03075_, _03072_);
  and (_03077_, _03076_, _01438_);
  nor (_03078_, _03077_, _03074_);
  not (_03079_, _03067_);
  and (_03080_, _03071_, _03079_);
  and (_03082_, _03080_, _03064_);
  and (_03083_, _03082_, _01408_);
  not (_03084_, _03060_);
  nor (_03085_, _03063_, _03084_);
  nor (_03086_, _03071_, _03067_);
  and (_03087_, _03086_, _03085_);
  and (_03088_, _03087_, _01427_);
  nor (_03089_, _03088_, _03083_);
  and (_03090_, _03089_, _03078_);
  nor (_03091_, _03071_, _03079_);
  and (_03092_, _03063_, _03084_);
  and (_03093_, _03092_, _03091_);
  and (_03094_, _03093_, _01401_);
  and (_03095_, _03092_, _03080_);
  and (_03096_, _03095_, _01417_);
  nor (_03097_, _03096_, _03094_);
  and (_03098_, _03085_, _03072_);
  and (_03099_, _03098_, _01435_);
  and (_03100_, _03092_, _03072_);
  and (_03101_, _03100_, _01440_);
  nor (_03102_, _03101_, _03099_);
  and (_03103_, _03102_, _03097_);
  and (_03104_, _03103_, _03090_);
  and (_03105_, _03091_, _03064_);
  and (_03106_, _03105_, _01431_);
  and (_03107_, _03086_, _03064_);
  and (_03108_, _03107_, _01414_);
  nor (_03109_, _03108_, _03106_);
  and (_03110_, _03085_, _03091_);
  and (_03111_, _03110_, _01423_);
  and (_03112_, _03075_, _03080_);
  and (_03113_, _03112_, _01406_);
  nor (_03114_, _03113_, _03111_);
  and (_03115_, _03114_, _03109_);
  and (_03116_, _03085_, _03080_);
  and (_03117_, _03116_, _01425_);
  and (_03118_, _03092_, _03086_);
  and (_03119_, _03118_, _01412_);
  nor (_03120_, _03119_, _03117_);
  and (_03121_, _03075_, _03086_);
  and (_03122_, _03121_, _01419_);
  and (_03123_, _03075_, _03091_);
  and (_03124_, _03123_, _01403_);
  nor (_03125_, _03124_, _03122_);
  and (_03126_, _03125_, _03120_);
  and (_03127_, _03126_, _03115_);
  and (_03128_, _03127_, _03104_);
  nor (_03129_, _03128_, _02839_);
  or (_03130_, _03129_, _02932_);
  nor (_03131_, _03130_, _03000_);
  nor (_03132_, _03131_, _02933_);
  and (_03133_, _02566_, _02527_);
  not (_03134_, _03133_);
  and (_03135_, _02566_, _02529_);
  not (_03136_, _03135_);
  and (_03137_, _02865_, _02529_);
  nor (_03138_, _03137_, _03022_);
  and (_03139_, _03138_, _03136_);
  and (_03140_, _03139_, _03134_);
  and (_03141_, _02566_, _02532_);
  not (_03142_, _03141_);
  and (_03143_, _02865_, _02532_);
  nor (_03144_, _03143_, _03042_);
  and (_03145_, _03144_, _03142_);
  and (_03146_, _02566_, _02523_);
  not (_03147_, _03146_);
  and (_03148_, _02865_, _02523_);
  nor (_03149_, _03148_, _03051_);
  and (_03150_, _03149_, _03147_);
  and (_03151_, _03150_, _03145_);
  and (_03152_, _03151_, _03140_);
  not (_03153_, _03152_);
  nor (_03154_, _03153_, _03132_);
  and (_03155_, _02865_, _02527_);
  nor (_03156_, _03152_, _02794_);
  nor (_03157_, _03156_, _03155_);
  not (_03158_, _03157_);
  nor (_03159_, _03158_, _03154_);
  and (_03160_, _03155_, \oc8051_golden_model_1.SP [3]);
  or (_03161_, _03160_, _03040_);
  or (_03162_, _03161_, _03159_);
  nand (_03163_, _02927_, _03040_);
  and (_03164_, _03163_, _03162_);
  nor (_03165_, _03164_, _02892_);
  not (_03166_, _02892_);
  nor (_03167_, _03166_, _02794_);
  nor (_03168_, _03167_, _03165_);
  nand (_03169_, _03168_, _02891_);
  nand (_03170_, _02890_, \oc8051_golden_model_1.SP [3]);
  and (_03171_, _03170_, _03169_);
  or (_03173_, _03171_, _02889_);
  and (_03174_, _02566_, _02504_);
  not (_03175_, _02889_);
  nor (_03176_, _03175_, _02927_);
  nor (_03177_, _03176_, _03174_);
  nand (_03178_, _03177_, _03173_);
  not (_03179_, _03174_);
  nor (_03180_, _03179_, _02794_);
  nor (_03181_, _03180_, _02799_);
  and (_03182_, _03181_, _03178_);
  not (_03183_, _02799_);
  nor (_03184_, _03183_, _02927_);
  or (_03185_, _03184_, _03182_);
  nand (_03186_, _03185_, _02888_);
  and (_03187_, _02887_, _02794_);
  not (_03188_, _03187_);
  and (_03189_, _03188_, _03186_);
  nor (_03190_, _02741_, _33836_);
  nor (_03191_, _02750_, _33639_);
  nor (_03192_, _03191_, _03190_);
  nor (_03193_, _02728_, _33557_);
  nor (_03194_, _02733_, _33391_);
  nor (_03195_, _03194_, _03193_);
  and (_03196_, _03195_, _03192_);
  nor (_03197_, _02744_, _34000_);
  nor (_03198_, _02752_, _33475_);
  nor (_03199_, _03198_, _03197_);
  nor (_03200_, _02746_, _33959_);
  nor (_03201_, _02722_, _33737_);
  nor (_03202_, _03201_, _03200_);
  and (_03203_, _03202_, _03199_);
  and (_03204_, _03203_, _03196_);
  nor (_03205_, _02726_, _33598_);
  nor (_03206_, _02706_, _33516_);
  nor (_03207_, _03206_, _03205_);
  nor (_03208_, _02719_, _33918_);
  nor (_03209_, _02731_, _33350_);
  nor (_03210_, _03209_, _03208_);
  and (_03211_, _03210_, _03207_);
  nor (_03212_, _02755_, _33794_);
  nor (_03213_, _02712_, _33434_);
  nor (_03214_, _03213_, _03212_);
  nor (_03215_, _02738_, _33877_);
  nor (_03216_, _02758_, _33684_);
  nor (_03217_, _03216_, _03215_);
  and (_03218_, _03217_, _03214_);
  and (_03219_, _03218_, _03211_);
  and (_03220_, _03219_, _03204_);
  nor (_03221_, _03220_, _02838_);
  not (_03222_, _03221_);
  not (_03223_, _03040_);
  and (_03224_, _03183_, _02931_);
  and (_03225_, _03224_, _03223_);
  nor (_03226_, _02884_, _02866_);
  and (_03227_, _03226_, _03175_);
  and (_03228_, _03227_, _03225_);
  and (_03229_, _03228_, _02988_);
  nor (_03230_, _03229_, _03222_);
  not (_03231_, _03230_);
  and (_03232_, _03100_, _01394_);
  and (_03233_, _03095_, _01355_);
  nor (_03234_, _03233_, _03232_);
  and (_03235_, _03093_, _01385_);
  and (_03236_, _03076_, _01389_);
  nor (_03237_, _03236_, _03235_);
  and (_03238_, _03237_, _03234_);
  and (_03239_, _03073_, _01392_);
  and (_03240_, _03082_, _01360_);
  nor (_03241_, _03240_, _03239_);
  and (_03242_, _03105_, _01371_);
  and (_03243_, _03116_, _01377_);
  nor (_03244_, _03243_, _03242_);
  and (_03245_, _03244_, _03241_);
  and (_03246_, _03245_, _03238_);
  and (_03247_, _03087_, _01382_);
  and (_03248_, _03123_, _01368_);
  nor (_03249_, _03248_, _03247_);
  and (_03250_, _03098_, _01387_);
  and (_03251_, _03121_, _01366_);
  nor (_03252_, _03251_, _03250_);
  and (_03253_, _03252_, _03249_);
  and (_03254_, _03110_, _01379_);
  and (_03255_, _03118_, _01357_);
  nor (_03256_, _03255_, _03254_);
  and (_03257_, _03107_, _01373_);
  and (_03258_, _03112_, _01362_);
  nor (_03259_, _03258_, _03257_);
  and (_03260_, _03259_, _03256_);
  and (_03261_, _03260_, _03253_);
  and (_03262_, _03261_, _03246_);
  nor (_03263_, _03262_, _02839_);
  not (_03264_, \oc8051_golden_model_1.SP [2]);
  nor (_03265_, _02946_, _03155_);
  and (_03266_, _03265_, _02891_);
  nor (_03267_, _03266_, _03264_);
  not (_03268_, _03267_);
  and (_03269_, _02968_, _02509_);
  not (_03270_, _03269_);
  and (_03271_, _03002_, _02504_);
  and (_03272_, _02855_, _02509_);
  and (_03273_, _03272_, _02797_);
  nor (_03274_, _03273_, _03271_);
  and (_03275_, _03274_, _03270_);
  and (_03276_, _03009_, _02509_);
  and (_03277_, _03002_, _02527_);
  nor (_03278_, _03277_, _03276_);
  and (_03279_, _03009_, _02527_);
  not (_03280_, _03279_);
  and (_03281_, _02968_, _02523_);
  and (_03282_, _02968_, _02527_);
  nor (_03283_, _03282_, _03281_);
  and (_03284_, _03283_, _03280_);
  and (_03285_, _03284_, _03278_);
  and (_03286_, _03285_, _03275_);
  and (_03287_, _03286_, _03268_);
  not (_03288_, _02966_);
  nor (_03289_, _02515_, _02523_);
  nor (_03290_, _03289_, _03288_);
  not (_03291_, _03290_);
  and (_03292_, _02966_, _02498_);
  not (_03293_, _03292_);
  and (_03294_, _02966_, _02875_);
  not (_03295_, _03294_);
  and (_03296_, _02968_, _02498_);
  not (_03297_, _02797_);
  and (_03298_, _02855_, _03297_);
  and (_03299_, _03298_, _02504_);
  nor (_03300_, _03299_, _03296_);
  and (_03301_, _03300_, _03295_);
  and (_03302_, _03301_, _03293_);
  and (_03303_, _03302_, _03291_);
  and (_03304_, _02855_, _02883_);
  nor (_03305_, _02496_, _02432_);
  and (_03306_, _03305_, _02968_);
  nor (_03307_, _03306_, _03304_);
  and (_03308_, _02855_, _02949_);
  and (_03309_, _02520_, _02506_);
  and (_03310_, _03309_, _02855_);
  nor (_03311_, _03310_, _03308_);
  and (_03312_, _03311_, _03307_);
  nor (_03313_, _03010_, _03003_);
  and (_03314_, _03313_, _03312_);
  and (_03315_, _02966_, _02864_);
  not (_03316_, _03315_);
  and (_03317_, _02968_, _02870_);
  and (_03318_, _02968_, _02864_);
  nor (_03319_, _03318_, _03317_);
  and (_03320_, _03319_, _03316_);
  and (_03321_, _03320_, _03314_);
  and (_03322_, _03321_, _03303_);
  and (_03323_, _03322_, _03287_);
  not (_03324_, _03323_);
  nor (_03325_, _03324_, _03263_);
  nor (_03326_, _02744_, _33985_);
  nor (_03327_, _02741_, _33821_);
  nor (_03328_, _03327_, _03326_);
  nor (_03329_, _02728_, _33542_);
  nor (_03330_, _02706_, _33501_);
  nor (_03331_, _03330_, _03329_);
  and (_03332_, _03331_, _03328_);
  nor (_03333_, _02746_, _33944_);
  nor (_03334_, _02719_, _33903_);
  nor (_03335_, _03334_, _03333_);
  nor (_03336_, _02755_, _33773_);
  nor (_03337_, _02722_, _33717_);
  nor (_03338_, _03337_, _03336_);
  and (_03339_, _03338_, _03335_);
  and (_03340_, _03339_, _03332_);
  nor (_03341_, _02752_, _33460_);
  nor (_03342_, _02712_, _33418_);
  nor (_03343_, _03342_, _03341_);
  nor (_03344_, _02750_, _33624_);
  nor (_03345_, _02731_, _33330_);
  nor (_03346_, _03345_, _03344_);
  and (_03347_, _03346_, _03343_);
  nor (_03348_, _02738_, _33862_);
  nor (_03349_, _02758_, _33665_);
  nor (_03350_, _03349_, _03348_);
  nor (_03351_, _02726_, _33583_);
  nor (_03352_, _02733_, _33376_);
  nor (_03353_, _03352_, _03351_);
  and (_03354_, _03353_, _03350_);
  and (_03355_, _03354_, _03347_);
  and (_03356_, _03355_, _03340_);
  and (_03357_, _02980_, _02952_);
  and (_03358_, _02565_, _02509_);
  and (_03359_, _03358_, _02563_);
  nor (_03360_, _03174_, _02887_);
  not (_03361_, _03360_);
  nor (_03362_, _03361_, _03359_);
  and (_03363_, _03362_, _03357_);
  and (_03364_, _03363_, _03152_);
  and (_03365_, _03364_, _02973_);
  nor (_03366_, _03365_, _03356_);
  not (_03367_, _03366_);
  and (_03368_, _03367_, _03325_);
  and (_03369_, _03368_, _03231_);
  not (_03370_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_03371_, _02979_, _02833_);
  not (_03372_, _02795_);
  nor (_03374_, _02942_, _03372_);
  and (_03375_, _02954_, _02833_);
  or (_03376_, _02992_, _02837_);
  and (_03377_, _02948_, _02833_);
  not (_03378_, _02593_);
  and (_03379_, _03024_, _03378_);
  and (_03380_, _03379_, _02495_);
  not (_03381_, _03380_);
  not (_03382_, _02602_);
  and (_03383_, _02865_, _03382_);
  nand (_03384_, _02336_, _02304_);
  nor (_03385_, _03384_, _02600_);
  nor (_03386_, _03385_, _03383_);
  and (_03387_, _03386_, _03381_);
  and (_03388_, _03002_, _02883_);
  nor (_03389_, _03388_, _02948_);
  and (_03390_, _03024_, _02883_);
  and (_03391_, _02849_, _02336_);
  and (_03392_, _03391_, _02883_);
  and (_03393_, _03047_, _02883_);
  and (_03394_, _02865_, _02949_);
  or (_03395_, _03394_, _03393_);
  or (_03396_, _03395_, _03392_);
  nor (_03397_, _03396_, _03390_);
  and (_03398_, _03397_, _03389_);
  and (_03399_, _03398_, _03387_);
  or (_03400_, _03399_, _03377_);
  not (_03401_, _02951_);
  or (_03402_, _03401_, _02833_);
  and (_03403_, _03402_, _02976_);
  nand (_03404_, _03403_, _03400_);
  and (_03405_, _02946_, \oc8051_golden_model_1.SP [0]);
  nor (_03406_, _02885_, _03405_);
  nand (_03407_, _03406_, _03404_);
  or (_03408_, _02850_, _03002_);
  nor (_03409_, _03408_, _03024_);
  or (_03410_, _03409_, _02594_);
  and (_03411_, _02962_, _02875_);
  nor (_03412_, _03411_, _02880_);
  and (_03413_, _02968_, _02875_);
  nand (_03414_, _03413_, _02336_);
  and (_03415_, _03414_, _03412_);
  and (_03416_, _03415_, _03410_);
  nand (_03417_, _03416_, _03407_);
  nand (_03418_, _03417_, _03376_);
  and (_03419_, _03418_, _02987_);
  or (_03420_, _02878_, _03419_);
  and (_03421_, _02876_, _02837_);
  and (_03422_, _03391_, _02870_);
  and (_03423_, _03317_, _02336_);
  or (_03424_, _02954_, _03025_);
  or (_03425_, _03424_, _03003_);
  or (_03426_, _03425_, _03423_);
  nor (_03427_, _03426_, _03422_);
  not (_03428_, _03427_);
  nor (_03429_, _03428_, _03421_);
  and (_03430_, _03429_, _03420_);
  or (_03431_, _03430_, _03375_);
  nand (_03432_, _03431_, _02938_);
  not (_03433_, _02971_);
  not (_03434_, _02938_);
  and (_03435_, _03434_, _02795_);
  nor (_03436_, _03435_, _03433_);
  nand (_03437_, _03436_, _03432_);
  and (_03438_, _03433_, _02837_);
  and (_03439_, _03024_, _02939_);
  not (_03440_, _03439_);
  and (_03441_, _03440_, _02942_);
  not (_03442_, _03441_);
  nor (_03443_, _03442_, _03438_);
  and (_03444_, _03443_, _03437_);
  or (_03445_, _03444_, _03374_);
  and (_03446_, _03318_, _02336_);
  not (_03447_, _03446_);
  and (_03448_, _02845_, _02864_);
  and (_03449_, _03448_, _02336_);
  not (_03450_, _03449_);
  and (_03451_, _03024_, _02864_);
  nor (_03452_, _03451_, _02979_);
  and (_03453_, _03452_, _03450_);
  and (_03454_, _02850_, _02864_);
  and (_03455_, _02855_, _02864_);
  and (_03456_, _03455_, _02797_);
  nor (_03457_, _03456_, _03454_);
  and (_03458_, _03457_, _03453_);
  and (_03459_, _03458_, _03447_);
  and (_03460_, _03459_, _03445_);
  or (_03461_, _03460_, _03371_);
  and (_03462_, _03461_, _02986_);
  or (_03463_, _03462_, _02867_);
  and (_03464_, _02855_, _02336_);
  nor (_03465_, _03464_, _02566_);
  nor (_03466_, _03465_, _02852_);
  not (_03467_, _03466_);
  and (_03468_, _02962_, _02515_);
  not (_03469_, _03468_);
  and (_03470_, _03024_, _02515_);
  nor (_03471_, _03470_, _02851_);
  and (_03472_, _03471_, _03469_);
  and (_03473_, _03472_, _03467_);
  and (_03474_, _03473_, _03463_);
  and (_03475_, _03095_, _01268_);
  and (_03476_, _03093_, _01281_);
  nor (_03477_, _03476_, _03475_);
  and (_03478_, _03105_, _01274_);
  and (_03479_, _03098_, _01297_);
  nor (_03480_, _03479_, _03478_);
  and (_03481_, _03480_, _03477_);
  and (_03482_, _03116_, _01285_);
  and (_03483_, _03110_, _01287_);
  nor (_03484_, _03483_, _03482_);
  and (_03485_, _03073_, _01295_);
  and (_03486_, _03107_, _01276_);
  nor (_03487_, _03486_, _03485_);
  and (_03488_, _03487_, _03484_);
  and (_03489_, _03488_, _03481_);
  and (_03490_, _03121_, _01263_);
  and (_03491_, _03112_, _01265_);
  nor (_03492_, _03491_, _03490_);
  and (_03493_, _03100_, _01300_);
  and (_03494_, _03118_, _01270_);
  nor (_03495_, _03494_, _03493_);
  and (_03496_, _03495_, _03492_);
  and (_03497_, _03082_, _01293_);
  and (_03498_, _03087_, _01290_);
  nor (_03499_, _03498_, _03497_);
  and (_03500_, _03076_, _01302_);
  and (_03501_, _03123_, _01279_);
  nor (_03502_, _03501_, _03500_);
  and (_03503_, _03502_, _03499_);
  and (_03504_, _03503_, _03496_);
  and (_03505_, _03504_, _03489_);
  nor (_03506_, _03505_, _02839_);
  or (_03507_, _03506_, _03474_);
  not (_03508_, _02930_);
  nor (_03509_, _03508_, _02795_);
  and (_03510_, _03024_, _02521_);
  nor (_03511_, _03510_, _02928_);
  not (_03512_, _03511_);
  nor (_03513_, _03512_, _03509_);
  and (_03514_, _03513_, _03507_);
  and (_03515_, _02928_, _02795_);
  or (_03516_, _03515_, _03514_);
  and (_03517_, _03002_, _02523_);
  not (_03518_, _03517_);
  and (_03519_, _03047_, _02523_);
  not (_03520_, _03519_);
  and (_03521_, _03024_, _02523_);
  and (_03522_, _03391_, _02523_);
  nor (_03523_, _03522_, _03521_);
  and (_03524_, _03523_, _03520_);
  and (_03525_, _03524_, _03518_);
  and (_03526_, _03525_, _03516_);
  nor (_03527_, _03150_, _02833_);
  not (_03528_, _02529_);
  nor (_03529_, _03024_, _02850_);
  nor (_03530_, _03529_, _03528_);
  not (_03531_, _03530_);
  and (_03532_, _02962_, _02529_);
  not (_03533_, _03532_);
  and (_03534_, _03002_, _02529_);
  and (_03535_, _03047_, _02529_);
  nor (_03536_, _03535_, _03534_);
  and (_03537_, _03536_, _03533_);
  and (_03538_, _03537_, _03531_);
  not (_03539_, _03538_);
  nor (_03540_, _03539_, _03527_);
  and (_03541_, _03540_, _03526_);
  nor (_03542_, _03139_, _02833_);
  not (_03543_, _02532_);
  nor (_03544_, _02850_, _03464_);
  nor (_03545_, _03024_, _02962_);
  and (_03546_, _03545_, _03544_);
  nor (_03547_, _03546_, _03543_);
  nor (_03548_, _03547_, _03542_);
  and (_03549_, _03548_, _03541_);
  nor (_03550_, _03145_, _02833_);
  not (_03551_, _02527_);
  nor (_03552_, _03544_, _03551_);
  not (_03553_, _03552_);
  and (_03554_, _02962_, _02527_);
  not (_03555_, _03554_);
  and (_03556_, _03024_, _02527_);
  nor (_03557_, _03556_, _03133_);
  and (_03558_, _03557_, _03555_);
  and (_03559_, _03558_, _03553_);
  not (_03560_, _03559_);
  nor (_03561_, _03560_, _03550_);
  and (_03562_, _03561_, _03549_);
  and (_03563_, _03133_, _02833_);
  or (_03564_, _03563_, _03562_);
  and (_03565_, _03155_, _02868_);
  nor (_03566_, _03565_, _03040_);
  and (_03567_, _03566_, _03564_);
  and (_03568_, _03040_, _02795_);
  or (_03569_, _03568_, _03567_);
  and (_03570_, _02850_, _02509_);
  and (_03571_, _03024_, _02509_);
  nor (_03572_, _03571_, _03570_);
  and (_03573_, _02962_, _02509_);
  not (_03575_, _02509_);
  nor (_03576_, _03465_, _03575_);
  nor (_03577_, _03576_, _03573_);
  and (_03578_, _03577_, _03572_);
  and (_03579_, _03578_, _03569_);
  and (_03580_, _02892_, _02833_);
  or (_03581_, _03580_, _03579_);
  and (_03582_, _02890_, _02868_);
  nor (_03583_, _03582_, _02889_);
  and (_03584_, _03583_, _03581_);
  and (_03585_, _02889_, _02795_);
  or (_03586_, _03585_, _03584_);
  and (_03587_, _02962_, _02504_);
  nor (_03588_, _03587_, _03174_);
  and (_03589_, _03024_, _02504_);
  not (_03590_, _03589_);
  and (_03591_, _03047_, _02504_);
  and (_03592_, _02850_, _02504_);
  or (_03593_, _03592_, _03271_);
  nor (_03594_, _03593_, _03591_);
  and (_03595_, _03594_, _03590_);
  and (_03596_, _03595_, _03588_);
  and (_03597_, _03596_, _03586_);
  and (_03598_, _03174_, _02833_);
  or (_03599_, _03598_, _03597_);
  and (_03600_, _03599_, _03183_);
  or (_03601_, _02800_, _03600_);
  and (_03602_, _03047_, _02498_);
  not (_03603_, _03602_);
  and (_03604_, _03024_, _02498_);
  nor (_03605_, _03604_, _02887_);
  and (_03606_, _03605_, _03603_);
  and (_03607_, _03002_, _02498_);
  and (_03608_, _02849_, _02498_);
  and (_03609_, _03608_, _02336_);
  nor (_03610_, _03609_, _03607_);
  and (_03611_, _03610_, _03606_);
  nand (_03612_, _03611_, _03601_);
  and (_03613_, _02887_, _02833_);
  not (_03614_, _03613_);
  nand (_03615_, _03614_, _03612_);
  or (_03616_, _03615_, _03370_);
  nor (_03617_, _02744_, _33995_);
  nor (_03618_, _02758_, _33678_);
  nor (_03619_, _03618_, _03617_);
  nor (_03620_, _02728_, _33552_);
  nor (_03621_, _02731_, _33345_);
  nor (_03622_, _03621_, _03620_);
  and (_03623_, _03622_, _03619_);
  nor (_03624_, _02750_, _33634_);
  nor (_03625_, _02706_, _33511_);
  nor (_03626_, _03625_, _03624_);
  nor (_03627_, _02746_, _33954_);
  nor (_03628_, _02738_, _33872_);
  nor (_03629_, _03628_, _03627_);
  and (_03630_, _03629_, _03626_);
  and (_03631_, _03630_, _03623_);
  nor (_03632_, _02755_, _33787_);
  nor (_03633_, _02722_, _33732_);
  nor (_03634_, _03633_, _03632_);
  nor (_03635_, _02752_, _33470_);
  nor (_03636_, _02733_, _33386_);
  nor (_03637_, _03636_, _03635_);
  and (_03638_, _03637_, _03634_);
  nor (_03639_, _02719_, _33913_);
  nor (_03640_, _02726_, _33593_);
  nor (_03641_, _03640_, _03639_);
  nor (_03642_, _02741_, _33831_);
  nor (_03643_, _02712_, _33429_);
  nor (_03644_, _03643_, _03642_);
  and (_03645_, _03644_, _03641_);
  and (_03646_, _03645_, _03638_);
  and (_03647_, _03646_, _03631_);
  nor (_03648_, _03647_, _02838_);
  and (_03649_, _03648_, _02866_);
  not (_03650_, _03649_);
  nor (_03651_, _02889_, _02884_);
  and (_03652_, _03651_, _03225_);
  and (_03653_, _03652_, _02988_);
  not (_03654_, _03653_);
  and (_03655_, _03654_, _03648_);
  not (_03656_, _03655_);
  nor (_03657_, _02758_, _33660_);
  nor (_03658_, _02706_, _33496_);
  nor (_03659_, _03658_, _03657_);
  nor (_03660_, _02744_, _33980_);
  nor (_03661_, _02750_, _33619_);
  nor (_03662_, _03661_, _03660_);
  and (_03663_, _03662_, _03659_);
  nor (_03664_, _02722_, _33710_);
  nor (_03665_, _02728_, _33537_);
  nor (_03666_, _03665_, _03664_);
  nor (_03667_, _02731_, _33319_);
  nor (_03668_, _02733_, _33371_);
  nor (_03669_, _03668_, _03667_);
  and (_03670_, _03669_, _03666_);
  and (_03671_, _03670_, _03663_);
  nor (_03672_, _02719_, _33898_);
  nor (_03673_, _02755_, _33766_);
  nor (_03674_, _03673_, _03672_);
  nor (_03675_, _02726_, _33578_);
  nor (_03676_, _02712_, _33412_);
  nor (_03677_, _03676_, _03675_);
  and (_03678_, _03677_, _03674_);
  nor (_03679_, _02741_, _33816_);
  nor (_03680_, _02738_, _33857_);
  nor (_03681_, _03680_, _03679_);
  nor (_03682_, _02746_, _33939_);
  nor (_03683_, _02752_, _33455_);
  nor (_03684_, _03683_, _03682_);
  and (_03685_, _03684_, _03681_);
  and (_03686_, _03685_, _03678_);
  and (_03687_, _03686_, _03671_);
  nor (_03688_, _03687_, _03365_);
  not (_03689_, _03688_);
  and (_03690_, _03100_, _01348_);
  and (_03691_, _03076_, _01343_);
  nor (_03692_, _03691_, _03690_);
  and (_03693_, _03073_, _01341_);
  and (_03694_, _03107_, _01322_);
  nor (_03695_, _03694_, _03693_);
  and (_03696_, _03695_, _03692_);
  and (_03697_, _03112_, _01311_);
  and (_03698_, _03123_, _01327_);
  nor (_03699_, _03698_, _03697_);
  and (_03700_, _03093_, _01339_);
  and (_03701_, _03118_, _01309_);
  nor (_03702_, _03701_, _03700_);
  and (_03703_, _03702_, _03699_);
  and (_03704_, _03703_, _03696_);
  and (_03705_, _03082_, _01320_);
  and (_03706_, _03105_, _01325_);
  nor (_03707_, _03706_, _03705_);
  and (_03708_, _03116_, _01333_);
  and (_03709_, _03087_, _01336_);
  nor (_03710_, _03709_, _03708_);
  and (_03711_, _03710_, _03707_);
  and (_03712_, _03095_, _01314_);
  and (_03713_, _03121_, _01316_);
  nor (_03714_, _03713_, _03712_);
  and (_03715_, _03098_, _01346_);
  and (_03716_, _03110_, _01331_);
  nor (_03717_, _03716_, _03715_);
  and (_03718_, _03717_, _03714_);
  and (_03719_, _03718_, _03711_);
  and (_03720_, _03719_, _03704_);
  nor (_03721_, _03720_, _02839_);
  and (_03722_, _02890_, \oc8051_golden_model_1.SP [1]);
  not (_03723_, _03722_);
  and (_03724_, _02968_, _02949_);
  nor (_03725_, _03724_, _03592_);
  and (_03726_, _03725_, _03723_);
  and (_03727_, _02854_, _02504_);
  and (_03728_, _02854_, _02509_);
  nor (_03729_, _03728_, _03727_);
  and (_03730_, _02854_, _02527_);
  and (_03731_, _02854_, _02515_);
  nor (_03732_, _03731_, _03730_);
  and (_03733_, _03732_, _03729_);
  and (_03734_, _02850_, _02527_);
  nor (_03735_, _03734_, _03269_);
  and (_03736_, _02956_, _02498_);
  nor (_03737_, _03736_, _03570_);
  and (_03738_, _03737_, _03735_);
  and (_03739_, _03738_, _03733_);
  and (_03740_, _03739_, _03726_);
  not (_03741_, \oc8051_golden_model_1.SP [1]);
  nor (_03742_, _03265_, _03741_);
  not (_03743_, _03742_);
  nor (_03744_, _02507_, _02401_);
  and (_03745_, _03744_, _02956_);
  not (_03746_, _03745_);
  and (_03747_, _03746_, _03319_);
  and (_03748_, _03747_, _03743_);
  nor (_03749_, _03306_, _03296_);
  and (_03750_, _02968_, _02883_);
  and (_03751_, _02968_, _02532_);
  nor (_03752_, _03751_, _03750_);
  and (_03753_, _03752_, _03749_);
  not (_03754_, _02851_);
  and (_03755_, _03754_, _03283_);
  and (_03756_, _03755_, _03753_);
  and (_03757_, _02956_, _02532_);
  and (_03758_, _02956_, _02529_);
  nor (_03759_, _03758_, _03757_);
  and (_03760_, _02956_, _02883_);
  and (_03761_, _02968_, _02504_);
  nor (_03762_, _03761_, _03760_);
  and (_03763_, _03762_, _03759_);
  and (_03764_, _02968_, _02529_);
  and (_03765_, _02956_, _02875_);
  nor (_03766_, _03765_, _03764_);
  and (_03767_, _02956_, _02864_);
  and (_03768_, _02956_, _02870_);
  nor (_03769_, _03768_, _03767_);
  and (_03770_, _03769_, _03766_);
  and (_03771_, _03770_, _03763_);
  and (_03772_, _03771_, _03756_);
  and (_03773_, _03772_, _03748_);
  and (_03774_, _03773_, _03740_);
  not (_03776_, _03774_);
  nor (_03777_, _03776_, _03721_);
  and (_03778_, _03777_, _03689_);
  and (_03779_, _03778_, _03656_);
  and (_03780_, _03779_, _03650_);
  nand (_03781_, _03615_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_03782_, _03781_, _03780_);
  nand (_03783_, _03782_, _03616_);
  not (_03784_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_03785_, _03614_, _03612_);
  or (_03786_, _03785_, _03784_);
  not (_03787_, _03780_);
  nand (_03788_, _03785_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_03789_, _03788_, _03787_);
  nand (_03790_, _03789_, _03786_);
  nand (_03791_, _03790_, _03783_);
  nand (_03792_, _03791_, _03369_);
  not (_03793_, _03369_);
  not (_03794_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_03795_, _03785_, _03794_);
  not (_03796_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_03797_, _03615_, _03796_);
  and (_03798_, _03797_, _03787_);
  nand (_03799_, _03798_, _03795_);
  not (_03800_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_03801_, _03615_, _03800_);
  not (_03802_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_03803_, _03785_, _03802_);
  and (_03804_, _03803_, _03780_);
  nand (_03805_, _03804_, _03801_);
  nand (_03806_, _03805_, _03799_);
  nand (_03807_, _03806_, _03793_);
  nand (_03808_, _03807_, _03792_);
  nand (_03809_, _03808_, _03189_);
  not (_03810_, _03189_);
  not (_03811_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_03812_, _03785_, _03811_);
  not (_03813_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_03814_, _03615_, _03813_);
  and (_03815_, _03814_, _03787_);
  nand (_03816_, _03815_, _03812_);
  not (_03817_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03818_, _03615_, _03817_);
  nand (_03819_, _03615_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_03820_, _03819_, _03780_);
  nand (_03821_, _03820_, _03818_);
  nand (_03822_, _03821_, _03816_);
  nand (_03823_, _03822_, _03369_);
  not (_03824_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_03825_, _03785_, _03824_);
  nand (_03826_, _03785_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_03827_, _03826_, _03787_);
  nand (_03828_, _03827_, _03825_);
  not (_03829_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_03830_, _03615_, _03829_);
  nand (_03831_, _03615_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_03832_, _03831_, _03780_);
  nand (_03833_, _03832_, _03830_);
  nand (_03834_, _03833_, _03828_);
  nand (_03835_, _03834_, _03793_);
  nand (_03836_, _03835_, _03823_);
  nand (_03837_, _03836_, _03810_);
  and (_03838_, _03837_, _03809_);
  and (_03839_, _02840_, _03382_);
  and (_03840_, _02840_, _02883_);
  nor (_03841_, _03840_, _03839_);
  or (_03842_, _03841_, _03838_);
  and (_03843_, _02948_, _02763_);
  not (_03844_, _03843_);
  and (_03845_, _03382_, _02566_);
  and (_03846_, _03845_, _02763_);
  nor (_03847_, _03384_, _02602_);
  nor (_03848_, _03847_, _03846_);
  not (_03849_, _02603_);
  and (_03850_, _03846_, _02833_);
  or (_03851_, _03850_, _03849_);
  or (_03852_, _03851_, _03848_);
  nor (_03853_, _02603_, _02868_);
  not (_03854_, _03853_);
  and (_03855_, _03464_, _02883_);
  nor (_03856_, _03392_, _03855_);
  and (_03857_, _03856_, _03854_);
  and (_03858_, _03857_, _03852_);
  and (_03859_, _03858_, _03844_);
  and (_03860_, _03859_, _03842_);
  and (_03861_, _03843_, _02833_);
  nor (_03862_, _03861_, _03860_);
  nor (_03863_, _03862_, _02886_);
  nor (_03864_, _03863_, _02885_);
  nor (_03865_, _02597_, _02868_);
  nor (_03866_, _03865_, _03864_);
  nor (_03867_, _03384_, _02594_);
  and (_03868_, _02946_, _02763_);
  and (_03869_, _03868_, _02837_);
  nor (_03870_, _03869_, _03867_);
  and (_03871_, _03870_, _03866_);
  nand (_03872_, _03837_, _03809_);
  and (_03873_, _02840_, _02875_);
  and (_03874_, _03873_, _03872_);
  nor (_03875_, _03874_, _02881_);
  and (_03876_, _03875_, _03871_);
  nor (_03877_, _03876_, _02882_);
  nor (_03878_, _03877_, _02879_);
  nor (_03879_, _03878_, _02878_);
  or (_03880_, _03879_, _02876_);
  nand (_03881_, _02876_, _02868_);
  nand (_03882_, _03881_, _03880_);
  and (_03883_, _03882_, _02874_);
  nor (_03884_, _03883_, _02872_);
  nor (_03885_, _03384_, _02588_);
  or (_03886_, _03885_, _03884_);
  nor (_03887_, _03886_, _02869_);
  and (_03888_, _02866_, _02763_);
  and (_03889_, _02840_, _02939_);
  and (_03890_, _03889_, _03872_);
  nor (_03891_, _03890_, _03888_);
  and (_03892_, _03891_, _03887_);
  nor (_03893_, _03892_, _02867_);
  nor (_03894_, _03893_, _02569_);
  and (_03895_, _02569_, _02868_);
  nor (_03896_, _03895_, _03894_);
  not (_03897_, _03384_);
  and (_03898_, _03897_, _02521_);
  or (_03899_, _03898_, _03896_);
  nor (_03900_, _03899_, _02863_);
  and (_03901_, _02840_, _02521_);
  and (_03902_, _03901_, _03872_);
  nor (_03903_, _03902_, _02835_);
  and (_03904_, _03903_, _03900_);
  nor (_03905_, _03904_, _02836_);
  nor (_03906_, _03905_, _02522_);
  and (_03907_, _02522_, _02868_);
  nor (_03908_, _03907_, _03906_);
  and (_03909_, _03137_, _02763_);
  and (_03910_, _03149_, _03023_);
  nor (_03911_, _03910_, _02838_);
  nor (_03912_, _03911_, _03909_);
  nor (_03913_, _03912_, _02833_);
  nor (_03914_, _03913_, _02530_);
  not (_03915_, _03914_);
  nor (_03916_, _03915_, _03908_);
  and (_03917_, _02530_, _02868_);
  nor (_03918_, _03917_, _03916_);
  not (_03919_, _03144_);
  and (_03920_, _03919_, _02763_);
  and (_03921_, _03920_, _02837_);
  nor (_03922_, _03921_, _02528_);
  not (_03923_, _03922_);
  nor (_03924_, _03923_, _03918_);
  and (_03925_, _02528_, _02868_);
  nor (_03926_, _03925_, _03924_);
  and (_03927_, _02840_, _02504_);
  and (_03928_, _03927_, _03872_);
  and (_03929_, _03174_, _02763_);
  and (_03930_, _03897_, _02504_);
  or (_03931_, _03930_, _03929_);
  or (_03932_, _03931_, _03928_);
  nor (_03933_, _03932_, _03926_);
  and (_03934_, _03929_, _02833_);
  nor (_03935_, _03934_, _03933_);
  nor (_03936_, _03034_, _02505_);
  nor (_03937_, _03936_, _02868_);
  nor (_03938_, _03937_, _03935_);
  and (_03939_, _03938_, _02802_);
  nor (_03940_, _03939_, _02800_);
  and (_03941_, _02840_, _02498_);
  and (_03942_, _03941_, _03872_);
  and (_03943_, _02887_, _02763_);
  and (_03944_, _03897_, _02498_);
  or (_03945_, _03944_, _03943_);
  or (_03946_, _03945_, _03942_);
  nor (_03947_, _03946_, _03940_);
  and (_03948_, _03943_, _02833_);
  nor (_03949_, _03948_, _03947_);
  not (_03950_, _03949_);
  not (_03951_, _03687_);
  and (_03952_, _03943_, _03951_);
  and (_03953_, _03648_, _02799_);
  and (_03954_, _03741_, \oc8051_golden_model_1.SP [0]);
  and (_03955_, \oc8051_golden_model_1.SP [1], _02868_);
  nor (_03956_, _03955_, _03954_);
  not (_03957_, _03956_);
  and (_03958_, _03957_, _02528_);
  and (_03959_, _03951_, _02835_);
  nor (_03960_, _03957_, _02591_);
  and (_03961_, _03957_, _02876_);
  not (_03962_, _02876_);
  and (_03963_, _03648_, _02884_);
  and (_03964_, _03843_, _03951_);
  not (_03965_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03966_, _03615_, _03965_);
  nand (_03967_, _03615_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_03968_, _03967_, _03780_);
  nand (_03969_, _03968_, _03966_);
  not (_03970_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_03971_, _03785_, _03970_);
  nand (_03972_, _03785_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_03973_, _03972_, _03787_);
  nand (_03974_, _03973_, _03971_);
  nand (_03975_, _03974_, _03969_);
  nand (_03977_, _03975_, _03369_);
  not (_03978_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_03979_, _03785_, _03978_);
  not (_03980_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03981_, _03615_, _03980_);
  and (_03982_, _03981_, _03787_);
  nand (_03983_, _03982_, _03979_);
  not (_03984_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_03985_, _03615_, _03984_);
  not (_03986_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_03987_, _03785_, _03986_);
  and (_03988_, _03987_, _03780_);
  nand (_03989_, _03988_, _03985_);
  nand (_03990_, _03989_, _03983_);
  nand (_03991_, _03990_, _03793_);
  nand (_03992_, _03991_, _03977_);
  nand (_03993_, _03992_, _03189_);
  not (_03994_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_03995_, _03785_, _03994_);
  nand (_03996_, _03785_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03997_, _03996_, _03787_);
  nand (_03998_, _03997_, _03995_);
  not (_03999_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_04000_, _03615_, _03999_);
  nand (_04001_, _03615_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_04002_, _04001_, _03780_);
  nand (_04003_, _04002_, _04000_);
  nand (_04004_, _04003_, _03998_);
  nand (_04005_, _04004_, _03369_);
  not (_04006_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_04007_, _03785_, _04006_);
  nand (_04008_, _03785_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_04009_, _04008_, _03787_);
  nand (_04010_, _04009_, _04007_);
  not (_04011_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_04012_, _03615_, _04011_);
  nand (_04013_, _03615_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_04014_, _04013_, _03780_);
  nand (_04015_, _04014_, _04012_);
  nand (_04016_, _04015_, _04010_);
  nand (_04017_, _04016_, _03793_);
  nand (_04018_, _04017_, _04005_);
  nand (_04019_, _04018_, _03810_);
  nand (_04020_, _04019_, _03993_);
  not (_04021_, _04020_);
  or (_04022_, _04021_, _03841_);
  and (_04023_, _02844_, _03382_);
  nor (_04024_, _04023_, _03846_);
  and (_04025_, _03846_, _03951_);
  or (_04026_, _04025_, _03849_);
  or (_04027_, _04026_, _04024_);
  and (_04028_, _02962_, _02883_);
  and (_04029_, _02959_, _02883_);
  nor (_04030_, _04029_, _04028_);
  nor (_04031_, _03957_, _02603_);
  and (_04032_, _02966_, _02883_);
  nor (_04033_, _04032_, _04031_);
  and (_04034_, _04033_, _04030_);
  and (_04035_, _04034_, _04027_);
  and (_04036_, _04035_, _03844_);
  and (_04037_, _04036_, _04022_);
  nor (_04038_, _04037_, _03964_);
  nor (_04039_, _04038_, _02886_);
  nor (_04040_, _04039_, _03963_);
  nor (_04041_, _03957_, _02597_);
  or (_04042_, _04041_, _04040_);
  and (_04043_, _02959_, _02875_);
  not (_04044_, _04043_);
  nor (_04045_, _03411_, _03294_);
  and (_04046_, _04045_, _04044_);
  not (_04047_, _04046_);
  and (_04048_, _03868_, _03687_);
  nor (_04049_, _04048_, _04047_);
  not (_04050_, _04049_);
  nor (_04051_, _04050_, _04042_);
  and (_04052_, _04020_, _03873_);
  nor (_04053_, _04052_, _02881_);
  and (_04054_, _04053_, _04051_);
  and (_04055_, _03951_, _02881_);
  nor (_04056_, _04055_, _04054_);
  and (_04057_, _03647_, _02879_);
  nor (_04058_, _04057_, _04056_);
  and (_04059_, _04058_, _03962_);
  nor (_04060_, _04059_, _03961_);
  and (_04061_, _03647_, _02873_);
  or (_04062_, _04061_, _04060_);
  not (_04063_, _02967_);
  nand (_04064_, _02964_, _04063_);
  or (_04065_, _04064_, _04062_);
  nor (_04066_, _04065_, _03960_);
  and (_04067_, _04020_, _03889_);
  nor (_04068_, _04067_, _03888_);
  and (_04069_, _04068_, _04066_);
  nor (_04070_, _04069_, _03649_);
  nor (_04071_, _04070_, _02569_);
  and (_04072_, _03957_, _02569_);
  nor (_04073_, _04072_, _04071_);
  and (_04074_, _02862_, _03687_);
  and (_04075_, _03009_, _02521_);
  and (_04076_, _02959_, _02521_);
  nor (_04077_, _04076_, _04075_);
  and (_04078_, _02962_, _02521_);
  and (_04079_, _03002_, _02521_);
  nor (_04080_, _04079_, _04078_);
  and (_04081_, _04080_, _04077_);
  not (_04082_, _04081_);
  nor (_04083_, _04082_, _04074_);
  not (_04084_, _04083_);
  nor (_04085_, _04084_, _04073_);
  and (_04086_, _04020_, _03901_);
  nor (_04087_, _04086_, _02835_);
  and (_04088_, _04087_, _04085_);
  nor (_04089_, _04088_, _03959_);
  nor (_04090_, _04089_, _02522_);
  and (_04091_, _03957_, _02522_);
  nor (_04092_, _04091_, _04090_);
  nor (_04093_, _03912_, _03951_);
  nor (_04094_, _04093_, _02530_);
  not (_04095_, _04094_);
  nor (_04096_, _04095_, _04092_);
  and (_04097_, _03957_, _02530_);
  nor (_04098_, _04097_, _04096_);
  and (_04099_, _03920_, _03687_);
  nor (_04100_, _04099_, _02528_);
  not (_04101_, _04100_);
  nor (_04102_, _04101_, _04098_);
  nor (_04103_, _04102_, _03958_);
  and (_04104_, _02959_, _02504_);
  nor (_04105_, _04104_, _03587_);
  and (_04106_, _02966_, _02504_);
  not (_04107_, _04106_);
  and (_04108_, _04107_, _04105_);
  not (_04109_, _04108_);
  nor (_04110_, _04109_, _04103_);
  and (_04111_, _04020_, _03927_);
  nor (_04112_, _04111_, _03929_);
  and (_04113_, _04112_, _04110_);
  and (_04114_, _03929_, _03951_);
  nor (_04115_, _04114_, _04113_);
  nor (_04116_, _03957_, _03936_);
  nor (_04117_, _04116_, _02801_);
  not (_04118_, _04117_);
  nor (_04119_, _04118_, _04115_);
  nor (_04120_, _04119_, _03953_);
  and (_04121_, _03608_, _02538_);
  nor (_04122_, _04121_, _04120_);
  and (_04123_, _04122_, _03293_);
  and (_04124_, _04020_, _03941_);
  nor (_04125_, _04124_, _03943_);
  and (_04126_, _04125_, _04123_);
  nor (_04127_, _04126_, _03952_);
  not (_04128_, _00000_);
  not (_04129_, _03909_);
  nor (_04130_, _03727_, _03593_);
  not (_04131_, _02522_);
  and (_04132_, _02531_, _04131_);
  and (_04133_, _02603_, _02597_);
  not (_04134_, _02569_);
  and (_04135_, _02591_, _04134_);
  and (_04136_, _04135_, _04133_);
  and (_04137_, _04136_, _04132_);
  not (_04138_, _02336_);
  and (_04139_, _03941_, _04138_);
  not (_04140_, _04139_);
  and (_04141_, _02850_, _02939_);
  nor (_04142_, _04043_, _04141_);
  and (_04143_, _04142_, _04140_);
  and (_04144_, _04143_, _04137_);
  and (_04145_, _04144_, _04130_);
  nor (_04146_, _03901_, _03889_);
  nor (_04147_, _03873_, _02876_);
  and (_04148_, _04147_, _04146_);
  and (_04149_, _02854_, _02939_);
  not (_04150_, _03936_);
  nor (_04151_, _04150_, _04149_);
  and (_04152_, _04151_, _04148_);
  nor (_04153_, _03604_, _03413_);
  and (_04154_, _04153_, _03841_);
  nor (_04155_, _03304_, _02969_);
  nor (_04156_, _03765_, _03760_);
  and (_04157_, _04156_, _04155_);
  and (_04158_, _04157_, _04154_);
  and (_04159_, _04158_, _04152_);
  and (_04160_, _02854_, _02498_);
  nor (_04161_, _04121_, _04160_);
  and (_04162_, _04161_, _04063_);
  nor (_04163_, _03609_, _03411_);
  nand (_04164_, _03391_, _02521_);
  and (_04165_, _04164_, _04163_);
  and (_04166_, _04165_, _04162_);
  and (_04167_, _04166_, _04159_);
  and (_04168_, _03298_, _02521_);
  nor (_04169_, _04168_, _04076_);
  and (_04170_, _04169_, _04030_);
  and (_04171_, _02854_, _02521_);
  nor (_04172_, _04171_, _04079_);
  and (_04173_, _04172_, _04105_);
  and (_04174_, _04173_, _04170_);
  and (_04175_, _02849_, _03382_);
  not (_04176_, _04175_);
  and (_04178_, _02855_, _03382_);
  nor (_04179_, _04178_, _03927_);
  and (_04180_, _04179_, _04176_);
  and (_04181_, _04180_, _03301_);
  and (_04182_, _03293_, _02964_);
  and (_04183_, _04182_, _04181_);
  and (_04184_, _04183_, _04174_);
  and (_04185_, _04184_, _04167_);
  and (_04186_, _04185_, _04145_);
  and (_04187_, _04186_, _04129_);
  nor (_04188_, _03911_, _02835_);
  nor (_04189_, _03868_, _02881_);
  and (_04190_, _04189_, _04188_);
  and (_04191_, _04190_, _04187_);
  and (_04192_, _02763_, _02567_);
  not (_04193_, _04192_);
  not (_04194_, _03845_);
  nor (_04195_, _02841_, _02846_);
  and (_04196_, _04195_, _04194_);
  and (_04197_, _04196_, _02858_);
  nor (_04198_, _04197_, _02838_);
  nor (_04199_, _02799_, _02877_);
  and (_04200_, _04199_, _02888_);
  and (_04201_, _04200_, _03226_);
  nor (_04202_, _04201_, _02838_);
  nor (_04203_, _04202_, _04198_);
  and (_04204_, _04203_, _04193_);
  nor (_04205_, _03843_, _02873_);
  nor (_04206_, _03929_, _03920_);
  and (_04207_, _04206_, _04205_);
  and (_04208_, _04207_, _04204_);
  and (_04209_, _04208_, _04191_);
  nor (_04210_, _04209_, _04128_);
  not (_04211_, _04210_);
  nor (_04212_, _04211_, _04127_);
  and (_04213_, _04212_, _03950_);
  and (_04214_, _02887_, _02795_);
  and (_04215_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04216_, _04215_, \oc8051_golden_model_1.SP [2]);
  or (_04217_, _04216_, \oc8051_golden_model_1.SP [3]);
  and (_04218_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04219_, _04218_, \oc8051_golden_model_1.SP [3]);
  nand (_04220_, _04219_, \oc8051_golden_model_1.SP [0]);
  and (_04221_, _04220_, _04217_);
  and (_04222_, _04221_, _02569_);
  not (_04223_, _04221_);
  nor (_04224_, _04223_, _02591_);
  not (_04225_, _02597_);
  and (_04226_, _02924_, _02886_);
  nand (_04227_, _03785_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand (_04228_, _03615_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_04229_, _04228_, _03780_);
  nand (_04230_, _04229_, _04227_);
  nand (_04231_, _03615_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand (_04232_, _03785_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_04233_, _04232_, _03787_);
  nand (_04234_, _04233_, _04231_);
  nand (_04235_, _04234_, _04230_);
  nand (_04236_, _04235_, _03369_);
  not (_04237_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_04238_, _03785_, _04237_);
  not (_04239_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04240_, _03615_, _04239_);
  and (_04241_, _04240_, _03787_);
  nand (_04242_, _04241_, _04238_);
  not (_04243_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04244_, _03615_, _04243_);
  not (_04245_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_04246_, _03785_, _04245_);
  and (_04247_, _04246_, _03780_);
  nand (_04248_, _04247_, _04244_);
  nand (_04249_, _04248_, _04242_);
  nand (_04250_, _04249_, _03793_);
  nand (_04251_, _04250_, _04236_);
  nand (_04252_, _04251_, _03189_);
  nand (_04253_, _03615_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_04254_, _03785_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_04255_, _04254_, _03787_);
  nand (_04256_, _04255_, _04253_);
  nand (_04257_, _03785_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_04258_, _03615_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_04259_, _04258_, _03780_);
  nand (_04260_, _04259_, _04257_);
  nand (_04261_, _04260_, _04256_);
  nand (_04262_, _04261_, _03369_);
  nand (_04263_, _03615_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_04264_, _03785_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_04265_, _04264_, _03787_);
  nand (_04266_, _04265_, _04263_);
  nand (_04267_, _03785_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_04268_, _03615_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_04269_, _04268_, _03780_);
  nand (_04270_, _04269_, _04267_);
  nand (_04271_, _04270_, _04266_);
  nand (_04272_, _04271_, _03793_);
  nand (_04273_, _04272_, _04262_);
  nand (_04274_, _04273_, _03810_);
  nand (_04275_, _04274_, _04252_);
  and (_04276_, _04275_, _03840_);
  nor (_04277_, _04223_, _02603_);
  nor (_04279_, _03839_, \oc8051_golden_model_1.PSW [3]);
  and (_04280_, _04275_, _03839_);
  or (_04281_, _04280_, _03846_);
  nor (_04282_, _04281_, _04279_);
  and (_04283_, _03845_, _02795_);
  nor (_04284_, _04283_, _04282_);
  nor (_04285_, _04284_, _03849_);
  or (_04286_, _04285_, _03840_);
  nor (_04287_, _04286_, _04277_);
  or (_04288_, _04287_, _03843_);
  nor (_04289_, _04288_, _04276_);
  and (_04290_, _03843_, _02794_);
  or (_04291_, _04290_, _02886_);
  nor (_04292_, _04291_, _04289_);
  nor (_04293_, _04292_, _04226_);
  nor (_04294_, _04293_, _04225_);
  nor (_04295_, _04221_, _02597_);
  nor (_04296_, _04295_, _03868_);
  not (_04297_, _04296_);
  nor (_04298_, _04297_, _04294_);
  and (_04299_, _03868_, _02794_);
  nor (_04300_, _04299_, _03873_);
  not (_04301_, _04300_);
  nor (_04302_, _04301_, _04298_);
  and (_04303_, _04275_, _03873_);
  nor (_04304_, _04303_, _02881_);
  not (_04305_, _04304_);
  nor (_04306_, _04305_, _04302_);
  and (_04307_, _02881_, _02794_);
  or (_04308_, _04307_, _02879_);
  nor (_04309_, _04308_, _04306_);
  and (_04310_, _02924_, _02879_);
  nor (_04311_, _04310_, _04309_);
  and (_04312_, _04311_, _03962_);
  and (_04313_, _04221_, _02876_);
  nor (_04314_, _04313_, _04312_);
  nor (_04315_, _04314_, _02873_);
  nor (_04316_, _02874_, _02927_);
  or (_04317_, _04316_, _04315_);
  and (_04318_, _04317_, _02591_);
  or (_04319_, _04318_, _03889_);
  nor (_04320_, _04319_, _04224_);
  and (_04321_, _04275_, _03889_);
  nor (_04322_, _04321_, _03888_);
  not (_04323_, _04322_);
  nor (_04324_, _04323_, _04320_);
  not (_04325_, _03888_);
  nor (_04326_, _04325_, _02927_);
  nor (_04327_, _04326_, _04324_);
  nor (_04328_, _04327_, _02569_);
  nor (_04329_, _04328_, _04222_);
  or (_04330_, _04329_, _02862_);
  and (_04331_, _02862_, _02794_);
  nor (_04332_, _04331_, _03901_);
  and (_04333_, _04332_, _04330_);
  and (_04334_, _04275_, _03901_);
  nor (_04335_, _04334_, _02835_);
  not (_04336_, _04335_);
  nor (_04337_, _04336_, _04333_);
  and (_04338_, _02795_, _02834_);
  nor (_04339_, _04338_, _04337_);
  nor (_04340_, _04339_, _02522_);
  and (_04341_, _04221_, _02522_);
  not (_04342_, _04341_);
  and (_04343_, _04342_, _03912_);
  not (_04344_, _04343_);
  nor (_04345_, _04344_, _04340_);
  nor (_04346_, _03912_, _02794_);
  nor (_04347_, _04346_, _02530_);
  not (_04348_, _04347_);
  nor (_04349_, _04348_, _04345_);
  and (_04350_, _04221_, _02530_);
  or (_04351_, _04350_, _03920_);
  nor (_04352_, _04351_, _04349_);
  not (_04353_, _02794_);
  and (_04354_, _03920_, _04353_);
  nor (_04355_, _04354_, _02528_);
  not (_04356_, _04355_);
  nor (_04357_, _04356_, _04352_);
  and (_04358_, _04221_, _02528_);
  nor (_04359_, _04358_, _03927_);
  not (_04360_, _04359_);
  nor (_04361_, _04360_, _04357_);
  and (_04362_, _04275_, _03927_);
  nor (_04363_, _04362_, _03929_);
  not (_04364_, _04363_);
  nor (_04365_, _04364_, _04361_);
  and (_04366_, _03174_, _02795_);
  nor (_04367_, _04366_, _04150_);
  not (_04368_, _04367_);
  nor (_04369_, _04368_, _04365_);
  nor (_04370_, _04221_, _03936_);
  nor (_04371_, _04370_, _02801_);
  not (_04372_, _04371_);
  nor (_04373_, _04372_, _04369_);
  not (_04374_, _02924_);
  and (_04375_, _02801_, _04374_);
  nor (_04376_, _04375_, _03941_);
  not (_04377_, _04376_);
  nor (_04378_, _04377_, _04373_);
  and (_04380_, _04275_, _03941_);
  nor (_04381_, _04380_, _03943_);
  not (_04382_, _04381_);
  nor (_04383_, _04382_, _04378_);
  nor (_04384_, _04383_, _04214_);
  not (_04385_, _03356_);
  and (_04386_, _03943_, _04385_);
  and (_04387_, _03221_, _02799_);
  nor (_04388_, _04215_, \oc8051_golden_model_1.SP [2]);
  nor (_04389_, _04388_, _04216_);
  and (_04390_, _04389_, _02528_);
  and (_04391_, _04385_, _02835_);
  and (_04392_, _02862_, _03356_);
  and (_04393_, _02849_, _02521_);
  and (_04394_, _04389_, _02876_);
  nand (_04395_, _03785_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand (_04396_, _03615_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_04397_, _04396_, _03780_);
  nand (_04398_, _04397_, _04395_);
  not (_04399_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_04400_, _03785_, _04399_);
  not (_04401_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_04402_, _03615_, _04401_);
  and (_04403_, _04402_, _03787_);
  nand (_04404_, _04403_, _04400_);
  nand (_04405_, _04404_, _04398_);
  nand (_04406_, _04405_, _03369_);
  not (_04407_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_04408_, _03785_, _04407_);
  not (_04409_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_04410_, _03615_, _04409_);
  and (_04411_, _04410_, _03787_);
  nand (_04412_, _04411_, _04408_);
  not (_04413_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_04414_, _03615_, _04413_);
  not (_04415_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_04416_, _03785_, _04415_);
  and (_04417_, _04416_, _03780_);
  nand (_04418_, _04417_, _04414_);
  nand (_04419_, _04418_, _04412_);
  nand (_04420_, _04419_, _03793_);
  nand (_04421_, _04420_, _04406_);
  nand (_04422_, _04421_, _03189_);
  not (_04423_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_04424_, _03785_, _04423_);
  not (_04425_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_04426_, _03615_, _04425_);
  and (_04427_, _04426_, _03787_);
  nand (_04428_, _04427_, _04424_);
  nand (_04429_, _03785_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_04430_, _03615_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_04431_, _04430_, _03780_);
  nand (_04432_, _04431_, _04429_);
  nand (_04433_, _04432_, _04428_);
  nand (_04434_, _04433_, _03369_);
  not (_04435_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_04436_, _03785_, _04435_);
  not (_04437_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_04438_, _03615_, _04437_);
  and (_04439_, _04438_, _03787_);
  nand (_04440_, _04439_, _04436_);
  nand (_04441_, _03785_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_04442_, _03615_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_04443_, _04442_, _03780_);
  nand (_04444_, _04443_, _04441_);
  nand (_04445_, _04444_, _04440_);
  nand (_04446_, _04445_, _03793_);
  nand (_04447_, _04446_, _04434_);
  nand (_04448_, _04447_, _03810_);
  nand (_04449_, _04448_, _04422_);
  not (_04450_, _04449_);
  or (_04451_, _04450_, _03841_);
  nor (_04452_, _04175_, _03846_);
  and (_04453_, _03846_, _04385_);
  or (_04454_, _04453_, _03849_);
  or (_04455_, _04454_, _04452_);
  nor (_04456_, _04389_, _02603_);
  not (_04457_, _04456_);
  not (_04458_, _03760_);
  and (_04459_, _04030_, _04458_);
  and (_04460_, _04459_, _04457_);
  and (_04461_, _04460_, _04455_);
  and (_04462_, _04461_, _03844_);
  and (_04463_, _04462_, _04451_);
  and (_04464_, _03843_, _04385_);
  nor (_04465_, _04464_, _04463_);
  and (_04466_, _03220_, _02886_);
  nor (_04467_, _04466_, _04465_);
  or (_04468_, _04389_, _02597_);
  nand (_04469_, _04468_, _04467_);
  and (_04470_, _03868_, _03356_);
  and (_04471_, _02849_, _02875_);
  nor (_04472_, _04471_, _04470_);
  not (_04473_, _04472_);
  nor (_04474_, _04473_, _04469_);
  and (_04475_, _04449_, _03873_);
  nor (_04476_, _04475_, _02881_);
  and (_04477_, _04476_, _04474_);
  and (_04478_, _04385_, _02881_);
  nor (_04479_, _04478_, _04477_);
  and (_04481_, _03220_, _02879_);
  nor (_04482_, _04481_, _04479_);
  and (_04483_, _04482_, _03962_);
  nor (_04484_, _04483_, _04394_);
  and (_04485_, _02873_, _03220_);
  or (_04486_, _04485_, _04484_);
  nor (_04487_, _04389_, _02591_);
  not (_04488_, _04487_);
  and (_04489_, _04488_, _02965_);
  not (_04490_, _04489_);
  nor (_04491_, _04490_, _04486_);
  and (_04492_, _04449_, _03889_);
  not (_04493_, _04492_);
  and (_04494_, _04493_, _04491_);
  and (_04495_, _03888_, _03220_);
  nor (_04496_, _04495_, _02569_);
  and (_04497_, _04496_, _04494_);
  and (_04498_, _04389_, _02569_);
  nor (_04499_, _04498_, _04497_);
  or (_04500_, _04499_, _04393_);
  nor (_04501_, _04500_, _04392_);
  and (_04502_, _04449_, _03901_);
  nor (_04503_, _04502_, _02835_);
  and (_04504_, _04503_, _04501_);
  nor (_04505_, _04504_, _04391_);
  nor (_04506_, _04505_, _02522_);
  and (_04507_, _04389_, _02522_);
  nor (_04508_, _04507_, _04506_);
  nor (_04509_, _03912_, _04385_);
  nor (_04510_, _04509_, _02530_);
  not (_04511_, _04510_);
  nor (_04512_, _04511_, _04508_);
  and (_04513_, _04389_, _02530_);
  nor (_04514_, _04513_, _04512_);
  and (_04515_, _03920_, _03356_);
  nor (_04516_, _04515_, _02528_);
  not (_04517_, _04516_);
  nor (_04518_, _04517_, _04514_);
  nor (_04519_, _04518_, _04390_);
  not (_04520_, _03727_);
  not (_04521_, _03592_);
  and (_04522_, _04105_, _04521_);
  and (_04523_, _04522_, _04520_);
  not (_04524_, _04523_);
  nor (_04525_, _04524_, _04519_);
  and (_04526_, _04449_, _03927_);
  nor (_04527_, _04526_, _03929_);
  and (_04528_, _04527_, _04525_);
  and (_04529_, _03929_, _04385_);
  nor (_04530_, _04529_, _04528_);
  nor (_04531_, _04389_, _03936_);
  nor (_04532_, _04531_, _02801_);
  not (_04533_, _04532_);
  nor (_04534_, _04533_, _04530_);
  nor (_04535_, _04534_, _04387_);
  nor (_04536_, _04535_, _03608_);
  and (_04537_, _04449_, _03941_);
  nor (_04538_, _04537_, _03943_);
  and (_04539_, _04538_, _04536_);
  nor (_04540_, _04539_, _04386_);
  nor (_04541_, _04540_, _04211_);
  not (_04542_, _04541_);
  nor (_04543_, _04542_, _04384_);
  and (_04544_, _04543_, _04213_);
  or (_04545_, _04544_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_04546_, _04218_, _02868_);
  nor (_04547_, _04389_, _03955_);
  nor (_04548_, _04547_, _04546_);
  and (_04549_, _04219_, _02868_);
  nor (_04550_, _04546_, _04221_);
  nor (_04551_, _04550_, _04549_);
  and (_04552_, _35182_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_04553_, _04552_);
  and (_04554_, _04137_, _03936_);
  nor (_04555_, _04554_, _04553_);
  and (_04556_, _04555_, _04551_);
  and (_04557_, _04556_, _04548_);
  and (_04558_, _04557_, _03954_);
  not (_04559_, _04558_);
  and (_04560_, _04559_, _04545_);
  not (_04561_, _04127_);
  nor (_04562_, _04553_, _04209_);
  not (_04563_, _04562_);
  nor (_04564_, _04563_, _03949_);
  and (_04565_, _04564_, _04561_);
  not (_04566_, _04540_);
  nor (_04567_, _04563_, _04384_);
  and (_04568_, _04567_, _04566_);
  and (_04569_, _04568_, _04565_);
  not (_04570_, _04569_);
  not (_04571_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_04572_, _03615_, _04571_);
  not (_04573_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_04574_, _03785_, _04573_);
  and (_04575_, _04574_, _03780_);
  nand (_04576_, _04575_, _04572_);
  not (_04577_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_04578_, _03785_, _04577_);
  not (_04579_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_04580_, _03615_, _04579_);
  and (_04582_, _04580_, _03787_);
  nand (_04583_, _04582_, _04578_);
  nand (_04584_, _04583_, _04576_);
  nand (_04585_, _04584_, _03369_);
  not (_04586_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_04587_, _03785_, _04586_);
  not (_04588_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_04589_, _03615_, _04588_);
  and (_04590_, _04589_, _03787_);
  nand (_04591_, _04590_, _04587_);
  not (_04592_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_04593_, _03615_, _04592_);
  not (_04594_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_04595_, _03785_, _04594_);
  and (_04596_, _04595_, _03780_);
  nand (_04597_, _04596_, _04593_);
  nand (_04598_, _04597_, _04591_);
  nand (_04599_, _04598_, _03793_);
  nand (_04600_, _04599_, _04585_);
  nand (_04601_, _04600_, _03189_);
  not (_04602_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_04603_, _03785_, _04602_);
  not (_04604_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_04605_, _03615_, _04604_);
  and (_04606_, _04605_, _03787_);
  nand (_04607_, _04606_, _04603_);
  nand (_04608_, _03785_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_04609_, _03615_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_04610_, _04609_, _03780_);
  nand (_04611_, _04610_, _04608_);
  nand (_04612_, _04611_, _04607_);
  nand (_04613_, _04612_, _03369_);
  not (_04614_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_04615_, _03785_, _04614_);
  not (_04616_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_04617_, _03615_, _04616_);
  and (_04618_, _04617_, _03787_);
  nand (_04619_, _04618_, _04615_);
  not (_04620_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_04621_, _03615_, _04620_);
  not (_04622_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_04623_, _03785_, _04622_);
  and (_04624_, _04623_, _03780_);
  nand (_04625_, _04624_, _04621_);
  nand (_04626_, _04625_, _04619_);
  nand (_04627_, _04626_, _03793_);
  nand (_04628_, _04627_, _04613_);
  nand (_04629_, _04628_, _03810_);
  nand (_04630_, _04629_, _04601_);
  or (_04631_, _04630_, _02838_);
  and (_04632_, _02924_, _02838_);
  and (_04633_, _04632_, _03220_);
  and (_04634_, _04633_, _03647_);
  and (_04635_, _04634_, _04353_);
  and (_04636_, _03687_, _02833_);
  and (_04637_, _04636_, _03356_);
  and (_04638_, _04637_, _04635_);
  and (_04639_, _04638_, \oc8051_golden_model_1.SP [7]);
  not (_04640_, _04639_);
  nor (_04641_, _03687_, _02833_);
  and (_04642_, _04641_, _03356_);
  and (_04643_, _04642_, _04635_);
  and (_04644_, _04643_, \oc8051_golden_model_1.DPL [7]);
  and (_04645_, _03687_, _02837_);
  and (_04646_, _04645_, _03356_);
  and (_04647_, _04646_, _02794_);
  and (_04648_, _04647_, _04634_);
  and (_04649_, _04648_, \oc8051_golden_model_1.TCON [7]);
  nor (_04650_, _04649_, _04644_);
  and (_04651_, _04650_, _04640_);
  and (_04652_, _03356_, _04353_);
  and (_04653_, _04645_, _04652_);
  and (_04654_, _04653_, _04634_);
  and (_04655_, _04654_, \oc8051_golden_model_1.P0 [7]);
  not (_04656_, _04655_);
  not (_04657_, _03647_);
  and (_04658_, _04657_, _03220_);
  and (_04659_, _04658_, _04632_);
  and (_04660_, _04659_, _04653_);
  and (_04661_, _04660_, \oc8051_golden_model_1.P1 [7]);
  not (_04662_, _04661_);
  not (_04663_, _03220_);
  and (_04664_, _03647_, _04663_);
  and (_04665_, _04664_, _04632_);
  and (_04666_, _04665_, _04653_);
  and (_04667_, _04666_, \oc8051_golden_model_1.P2 [7]);
  nor (_04668_, _03647_, _03220_);
  and (_04669_, _04668_, _04632_);
  and (_04670_, _04669_, _04653_);
  and (_04671_, _04670_, \oc8051_golden_model_1.P3 [7]);
  nor (_04672_, _04671_, _04667_);
  and (_04673_, _04672_, _04662_);
  and (_04674_, _04673_, _04656_);
  and (_04675_, _04674_, _04651_);
  nand (_04676_, _03356_, _02794_);
  nor (_04677_, _03687_, _02837_);
  not (_04678_, _04677_);
  nor (_04679_, _04678_, _04676_);
  and (_04680_, _04679_, _04634_);
  and (_04681_, _04680_, \oc8051_golden_model_1.TL1 [7]);
  nor (_04683_, _03356_, _04353_);
  and (_04684_, _04683_, _04636_);
  and (_04685_, _04684_, _04634_);
  and (_04686_, _04685_, \oc8051_golden_model_1.TH1 [7]);
  nor (_04687_, _04686_, _04681_);
  and (_04688_, _04637_, _02794_);
  and (_04689_, _04688_, _04634_);
  and (_04690_, _04689_, \oc8051_golden_model_1.TMOD [7]);
  and (_04691_, _04659_, _04647_);
  and (_04692_, _04691_, \oc8051_golden_model_1.SCON [7]);
  nor (_04693_, _04692_, _04690_);
  and (_04694_, _04693_, _04687_);
  and (_04695_, _04677_, _03356_);
  and (_04696_, _04695_, _04635_);
  and (_04697_, _04696_, \oc8051_golden_model_1.DPH [7]);
  not (_04698_, _04697_);
  not (_04699_, _04641_);
  nor (_04700_, _04676_, _04699_);
  and (_04701_, _04700_, _04634_);
  and (_04702_, _04701_, \oc8051_golden_model_1.TL0 [7]);
  and (_04703_, _04683_, _04645_);
  and (_04704_, _04703_, _04634_);
  and (_04705_, _04704_, \oc8051_golden_model_1.TH0 [7]);
  nor (_04706_, _04705_, _04702_);
  and (_04707_, _04706_, _04698_);
  and (_04708_, _04707_, _04694_);
  and (_04709_, _04677_, _04385_);
  and (_04710_, _04709_, _04635_);
  and (_04711_, _04710_, \oc8051_golden_model_1.PCON [7]);
  not (_04712_, _04711_);
  and (_04713_, _04669_, _04647_);
  and (_04714_, _04713_, \oc8051_golden_model_1.IP [7]);
  not (_04715_, _04714_);
  nor (_04716_, _02924_, _02763_);
  and (_04717_, _04716_, _04658_);
  and (_04718_, _04717_, _04653_);
  and (_04719_, _04718_, \oc8051_golden_model_1.PSW [7]);
  and (_04720_, _04716_, _04668_);
  and (_04721_, _04720_, _04653_);
  and (_04722_, _04721_, \oc8051_golden_model_1.B [7]);
  nor (_04723_, _04722_, _04719_);
  and (_04724_, _04723_, _04715_);
  and (_04725_, _04688_, _04659_);
  and (_04726_, _04725_, \oc8051_golden_model_1.SBUF [7]);
  not (_04727_, _04726_);
  and (_04728_, _04665_, _04647_);
  and (_04729_, _04728_, \oc8051_golden_model_1.IE [7]);
  and (_04730_, _04716_, _04664_);
  and (_04731_, _04730_, _04653_);
  and (_04732_, _04731_, \oc8051_golden_model_1.ACC [7]);
  nor (_04733_, _04732_, _04729_);
  and (_04734_, _04733_, _04727_);
  and (_04735_, _04734_, _04724_);
  and (_04736_, _04735_, _04712_);
  and (_04737_, _04736_, _04708_);
  and (_04738_, _04737_, _04675_);
  and (_04739_, _04738_, _04631_);
  not (_04740_, _04739_);
  nand (_04741_, _03785_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand (_04742_, _03615_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_04743_, _04742_, _03780_);
  nand (_04744_, _04743_, _04741_);
  nand (_04745_, _03615_, \oc8051_golden_model_1.IRAM[3] [6]);
  nand (_04746_, _03785_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_04747_, _04746_, _03787_);
  nand (_04748_, _04747_, _04745_);
  nand (_04749_, _04748_, _04744_);
  nand (_04750_, _04749_, _03369_);
  not (_04751_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_04752_, _03785_, _04751_);
  not (_04753_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_04754_, _03615_, _04753_);
  and (_04755_, _04754_, _03787_);
  nand (_04756_, _04755_, _04752_);
  not (_04757_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_04758_, _03615_, _04757_);
  not (_04759_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_04760_, _03785_, _04759_);
  and (_04761_, _04760_, _03780_);
  nand (_04762_, _04761_, _04758_);
  nand (_04763_, _04762_, _04756_);
  nand (_04764_, _04763_, _03793_);
  nand (_04765_, _04764_, _04750_);
  nand (_04766_, _04765_, _03189_);
  nand (_04767_, _03615_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_04768_, _03785_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_04769_, _04768_, _03787_);
  nand (_04770_, _04769_, _04767_);
  nand (_04771_, _03785_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_04772_, _03615_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_04773_, _04772_, _03780_);
  nand (_04774_, _04773_, _04771_);
  nand (_04775_, _04774_, _04770_);
  nand (_04776_, _04775_, _03369_);
  nand (_04777_, _03615_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_04778_, _03785_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_04779_, _04778_, _03787_);
  nand (_04780_, _04779_, _04777_);
  nand (_04781_, _03785_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_04782_, _03615_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_04784_, _04782_, _03780_);
  nand (_04785_, _04784_, _04781_);
  nand (_04786_, _04785_, _04780_);
  nand (_04787_, _04786_, _03793_);
  nand (_04788_, _04787_, _04776_);
  nand (_04789_, _04788_, _03810_);
  nand (_04790_, _04789_, _04766_);
  or (_04791_, _04790_, _02838_);
  and (_04792_, _04638_, \oc8051_golden_model_1.SP [6]);
  and (_04793_, _04643_, \oc8051_golden_model_1.DPL [6]);
  nor (_04794_, _04793_, _04792_);
  nand (_04795_, _04696_, \oc8051_golden_model_1.DPH [6]);
  and (_04796_, _04795_, _04794_);
  and (_04797_, _04648_, \oc8051_golden_model_1.TCON [6]);
  not (_04798_, _04797_);
  and (_04799_, _04701_, \oc8051_golden_model_1.TL0 [6]);
  and (_04800_, _04691_, \oc8051_golden_model_1.SCON [6]);
  nor (_04801_, _04800_, _04799_);
  and (_04802_, _04801_, _04798_);
  and (_04803_, _04704_, \oc8051_golden_model_1.TH0 [6]);
  and (_04804_, _04685_, \oc8051_golden_model_1.TH1 [6]);
  nor (_04805_, _04804_, _04803_);
  and (_04806_, _04689_, \oc8051_golden_model_1.TMOD [6]);
  and (_04807_, _04680_, \oc8051_golden_model_1.TL1 [6]);
  nor (_04808_, _04807_, _04806_);
  and (_04809_, _04808_, _04805_);
  and (_04810_, _04809_, _04802_);
  and (_04811_, _04810_, _04796_);
  and (_04812_, _04725_, \oc8051_golden_model_1.SBUF [6]);
  and (_04813_, _04728_, \oc8051_golden_model_1.IE [6]);
  nor (_04814_, _04813_, _04812_);
  not (_04815_, _04814_);
  and (_04816_, _04710_, \oc8051_golden_model_1.PCON [6]);
  nor (_04817_, _04816_, _04815_);
  and (_04818_, _04654_, \oc8051_golden_model_1.P0 [6]);
  not (_04819_, _04818_);
  and (_04820_, _04713_, \oc8051_golden_model_1.IP [6]);
  and (_04821_, _04721_, \oc8051_golden_model_1.B [6]);
  nor (_04822_, _04821_, _04820_);
  and (_04823_, _04718_, \oc8051_golden_model_1.PSW [6]);
  and (_04824_, _04731_, \oc8051_golden_model_1.ACC [6]);
  nor (_04825_, _04824_, _04823_);
  and (_04826_, _04825_, _04822_);
  and (_04827_, _04660_, \oc8051_golden_model_1.P1 [6]);
  not (_04828_, _04827_);
  and (_04829_, _04666_, \oc8051_golden_model_1.P2 [6]);
  and (_04830_, _04670_, \oc8051_golden_model_1.P3 [6]);
  nor (_04831_, _04830_, _04829_);
  and (_04832_, _04831_, _04828_);
  and (_04833_, _04832_, _04826_);
  and (_04834_, _04833_, _04819_);
  and (_04835_, _04834_, _04817_);
  and (_04836_, _04835_, _04811_);
  and (_04837_, _04836_, _04791_);
  not (_04838_, _04837_);
  nand (_04839_, _03785_, \oc8051_golden_model_1.IRAM[0] [5]);
  not (_04840_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_04841_, _03785_, _04840_);
  and (_04842_, _04841_, _03780_);
  nand (_04843_, _04842_, _04839_);
  nand (_04844_, _03615_, \oc8051_golden_model_1.IRAM[3] [5]);
  not (_04845_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_04846_, _03615_, _04845_);
  and (_04847_, _04846_, _03787_);
  nand (_04848_, _04847_, _04844_);
  nand (_04849_, _04848_, _04843_);
  nand (_04850_, _04849_, _03369_);
  not (_04851_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_04852_, _03785_, _04851_);
  not (_04853_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_04854_, _03615_, _04853_);
  and (_04855_, _04854_, _03787_);
  nand (_04856_, _04855_, _04852_);
  not (_04857_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_04858_, _03615_, _04857_);
  not (_04859_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_04860_, _03785_, _04859_);
  and (_04861_, _04860_, _03780_);
  nand (_04862_, _04861_, _04858_);
  nand (_04863_, _04862_, _04856_);
  nand (_04864_, _04863_, _03793_);
  nand (_04865_, _04864_, _04850_);
  nand (_04866_, _04865_, _03189_);
  nand (_04867_, _03615_, \oc8051_golden_model_1.IRAM[11] [5]);
  not (_04868_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_04869_, _03615_, _04868_);
  and (_04870_, _04869_, _03787_);
  nand (_04871_, _04870_, _04867_);
  nand (_04872_, _03785_, \oc8051_golden_model_1.IRAM[8] [5]);
  not (_04873_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_04874_, _03785_, _04873_);
  and (_04875_, _04874_, _03780_);
  nand (_04876_, _04875_, _04872_);
  nand (_04877_, _04876_, _04871_);
  nand (_04878_, _04877_, _03369_);
  nand (_04879_, _03615_, \oc8051_golden_model_1.IRAM[15] [5]);
  not (_04880_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_04881_, _03615_, _04880_);
  and (_04882_, _04881_, _03787_);
  nand (_04883_, _04882_, _04879_);
  nand (_04885_, _03785_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_04886_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_04887_, _03785_, _04886_);
  and (_04888_, _04887_, _03780_);
  nand (_04889_, _04888_, _04885_);
  nand (_04890_, _04889_, _04883_);
  nand (_04891_, _04890_, _03793_);
  nand (_04892_, _04891_, _04878_);
  nand (_04893_, _04892_, _03810_);
  nand (_04894_, _04893_, _04866_);
  or (_04895_, _04894_, _02838_);
  and (_04896_, _04638_, \oc8051_golden_model_1.SP [5]);
  not (_04897_, _04896_);
  and (_04898_, _04643_, \oc8051_golden_model_1.DPL [5]);
  and (_04899_, _04648_, \oc8051_golden_model_1.TCON [5]);
  nor (_04900_, _04899_, _04898_);
  and (_04901_, _04900_, _04897_);
  and (_04902_, _04654_, \oc8051_golden_model_1.P0 [5]);
  not (_04903_, _04902_);
  and (_04904_, _04660_, \oc8051_golden_model_1.P1 [5]);
  not (_04905_, _04904_);
  and (_04906_, _04666_, \oc8051_golden_model_1.P2 [5]);
  and (_04907_, _04670_, \oc8051_golden_model_1.P3 [5]);
  nor (_04908_, _04907_, _04906_);
  and (_04909_, _04908_, _04905_);
  and (_04910_, _04909_, _04903_);
  and (_04911_, _04910_, _04901_);
  and (_04912_, _04689_, \oc8051_golden_model_1.TMOD [5]);
  and (_04913_, _04685_, \oc8051_golden_model_1.TH1 [5]);
  nor (_04914_, _04913_, _04912_);
  and (_04915_, _04701_, \oc8051_golden_model_1.TL0 [5]);
  and (_04916_, _04680_, \oc8051_golden_model_1.TL1 [5]);
  nor (_04917_, _04916_, _04915_);
  and (_04918_, _04917_, _04914_);
  and (_04919_, _04696_, \oc8051_golden_model_1.DPH [5]);
  not (_04920_, _04919_);
  and (_04921_, _04704_, \oc8051_golden_model_1.TH0 [5]);
  and (_04922_, _04691_, \oc8051_golden_model_1.SCON [5]);
  nor (_04923_, _04922_, _04921_);
  and (_04924_, _04923_, _04920_);
  and (_04925_, _04924_, _04918_);
  and (_04926_, _04710_, \oc8051_golden_model_1.PCON [5]);
  not (_04927_, _04926_);
  and (_04928_, _04718_, \oc8051_golden_model_1.PSW [5]);
  not (_04929_, _04928_);
  and (_04930_, _04713_, \oc8051_golden_model_1.IP [5]);
  and (_04931_, _04731_, \oc8051_golden_model_1.ACC [5]);
  nor (_04932_, _04931_, _04930_);
  and (_04933_, _04932_, _04929_);
  and (_04934_, _04725_, \oc8051_golden_model_1.SBUF [5]);
  not (_04935_, _04934_);
  and (_04936_, _04728_, \oc8051_golden_model_1.IE [5]);
  and (_04937_, _04721_, \oc8051_golden_model_1.B [5]);
  nor (_04938_, _04937_, _04936_);
  and (_04939_, _04938_, _04935_);
  and (_04940_, _04939_, _04933_);
  and (_04941_, _04940_, _04927_);
  and (_04942_, _04941_, _04925_);
  and (_04943_, _04942_, _04911_);
  and (_04944_, _04943_, _04895_);
  not (_04945_, _04944_);
  or (_04946_, _04275_, _02838_);
  and (_04947_, _04638_, \oc8051_golden_model_1.SP [3]);
  and (_04948_, _04643_, \oc8051_golden_model_1.DPL [3]);
  nor (_04949_, _04948_, _04947_);
  nand (_04950_, _04696_, \oc8051_golden_model_1.DPH [3]);
  and (_04951_, _04950_, _04949_);
  and (_04952_, _04648_, \oc8051_golden_model_1.TCON [3]);
  not (_04953_, _04952_);
  and (_04954_, _04701_, \oc8051_golden_model_1.TL0 [3]);
  and (_04955_, _04691_, \oc8051_golden_model_1.SCON [3]);
  nor (_04956_, _04955_, _04954_);
  and (_04957_, _04956_, _04953_);
  and (_04958_, _04704_, \oc8051_golden_model_1.TH0 [3]);
  and (_04959_, _04685_, \oc8051_golden_model_1.TH1 [3]);
  nor (_04960_, _04959_, _04958_);
  and (_04961_, _04689_, \oc8051_golden_model_1.TMOD [3]);
  and (_04962_, _04680_, \oc8051_golden_model_1.TL1 [3]);
  nor (_04963_, _04962_, _04961_);
  and (_04964_, _04963_, _04960_);
  and (_04965_, _04964_, _04957_);
  and (_04966_, _04965_, _04951_);
  and (_04967_, _04725_, \oc8051_golden_model_1.SBUF [3]);
  and (_04968_, _04728_, \oc8051_golden_model_1.IE [3]);
  nor (_04969_, _04968_, _04967_);
  not (_04970_, _04969_);
  and (_04971_, _04710_, \oc8051_golden_model_1.PCON [3]);
  nor (_04972_, _04971_, _04970_);
  and (_04973_, _04654_, \oc8051_golden_model_1.P0 [3]);
  not (_04974_, _04973_);
  and (_04975_, _04713_, \oc8051_golden_model_1.IP [3]);
  and (_04976_, _04721_, \oc8051_golden_model_1.B [3]);
  nor (_04977_, _04976_, _04975_);
  and (_04978_, _04718_, \oc8051_golden_model_1.PSW [3]);
  and (_04979_, _04731_, \oc8051_golden_model_1.ACC [3]);
  nor (_04980_, _04979_, _04978_);
  and (_04981_, _04980_, _04977_);
  and (_04982_, _04660_, \oc8051_golden_model_1.P1 [3]);
  not (_04983_, _04982_);
  and (_04984_, _04666_, \oc8051_golden_model_1.P2 [3]);
  and (_04985_, _04670_, \oc8051_golden_model_1.P3 [3]);
  nor (_04986_, _04985_, _04984_);
  and (_04987_, _04986_, _04983_);
  and (_04988_, _04987_, _04981_);
  and (_04989_, _04988_, _04974_);
  and (_04990_, _04989_, _04972_);
  and (_04991_, _04990_, _04966_);
  and (_04992_, _04991_, _04946_);
  not (_04993_, _04992_);
  or (_04994_, _04020_, _02838_);
  and (_04995_, _04725_, \oc8051_golden_model_1.SBUF [1]);
  and (_04996_, _04728_, \oc8051_golden_model_1.IE [1]);
  nor (_04997_, _04996_, _04995_);
  nand (_04998_, _04710_, \oc8051_golden_model_1.PCON [1]);
  and (_04999_, _04998_, _04997_);
  and (_05000_, _04666_, \oc8051_golden_model_1.P2 [1]);
  and (_05001_, _04670_, \oc8051_golden_model_1.P3 [1]);
  nor (_05002_, _05001_, _05000_);
  and (_05003_, _05002_, _04999_);
  and (_05004_, _04718_, \oc8051_golden_model_1.PSW [1]);
  and (_05005_, _04721_, \oc8051_golden_model_1.B [1]);
  nor (_05006_, _05005_, _05004_);
  and (_05007_, _04713_, \oc8051_golden_model_1.IP [1]);
  and (_05008_, _04731_, \oc8051_golden_model_1.ACC [1]);
  nor (_05009_, _05008_, _05007_);
  and (_05010_, _05009_, _05006_);
  and (_05011_, _04648_, \oc8051_golden_model_1.TCON [1]);
  and (_05012_, _04704_, \oc8051_golden_model_1.TH0 [1]);
  nor (_05013_, _05012_, _05011_);
  and (_05014_, _04660_, \oc8051_golden_model_1.P1 [1]);
  and (_05015_, _04680_, \oc8051_golden_model_1.TL1 [1]);
  nor (_05016_, _05015_, _05014_);
  and (_05017_, _05016_, _05013_);
  and (_05018_, _04691_, \oc8051_golden_model_1.SCON [1]);
  and (_05019_, _04685_, \oc8051_golden_model_1.TH1 [1]);
  nor (_05020_, _05019_, _05018_);
  and (_05021_, _04701_, \oc8051_golden_model_1.TL0 [1]);
  and (_05022_, _04689_, \oc8051_golden_model_1.TMOD [1]);
  nor (_05023_, _05022_, _05021_);
  and (_05024_, _05023_, _05020_);
  and (_05025_, _05024_, _05017_);
  and (_05026_, _05025_, _05010_);
  and (_05027_, _05026_, _05003_);
  and (_05028_, _04654_, \oc8051_golden_model_1.P0 [1]);
  not (_05029_, _05028_);
  and (_05030_, _04638_, \oc8051_golden_model_1.SP [1]);
  and (_05031_, _04643_, \oc8051_golden_model_1.DPL [1]);
  nor (_05032_, _05031_, _05030_);
  nand (_05033_, _04696_, \oc8051_golden_model_1.DPH [1]);
  and (_05034_, _05033_, _05032_);
  and (_05035_, _05034_, _05029_);
  and (_05036_, _05035_, _05027_);
  and (_05037_, _05036_, _04994_);
  not (_05038_, _05037_);
  or (_05039_, _03872_, _02838_);
  and (_05040_, _04638_, \oc8051_golden_model_1.SP [0]);
  and (_05041_, _04643_, \oc8051_golden_model_1.DPL [0]);
  nor (_05042_, _05041_, _05040_);
  nand (_05043_, _04696_, \oc8051_golden_model_1.DPH [0]);
  and (_05044_, _05043_, _05042_);
  and (_05045_, _04648_, \oc8051_golden_model_1.TCON [0]);
  not (_05046_, _05045_);
  and (_05047_, _04701_, \oc8051_golden_model_1.TL0 [0]);
  and (_05048_, _04691_, \oc8051_golden_model_1.SCON [0]);
  nor (_05049_, _05048_, _05047_);
  and (_05050_, _05049_, _05046_);
  and (_05051_, _04704_, \oc8051_golden_model_1.TH0 [0]);
  and (_05052_, _04685_, \oc8051_golden_model_1.TH1 [0]);
  nor (_05053_, _05052_, _05051_);
  and (_05054_, _04689_, \oc8051_golden_model_1.TMOD [0]);
  and (_05055_, _04680_, \oc8051_golden_model_1.TL1 [0]);
  nor (_05056_, _05055_, _05054_);
  and (_05057_, _05056_, _05053_);
  and (_05058_, _05057_, _05050_);
  and (_05059_, _05058_, _05044_);
  and (_05060_, _04725_, \oc8051_golden_model_1.SBUF [0]);
  and (_05061_, _04728_, \oc8051_golden_model_1.IE [0]);
  nor (_05062_, _05061_, _05060_);
  not (_05063_, _05062_);
  and (_05064_, _04710_, \oc8051_golden_model_1.PCON [0]);
  nor (_05065_, _05064_, _05063_);
  and (_05066_, _04654_, \oc8051_golden_model_1.P0 [0]);
  not (_05067_, _05066_);
  and (_05068_, _04713_, \oc8051_golden_model_1.IP [0]);
  and (_05069_, _04721_, \oc8051_golden_model_1.B [0]);
  nor (_05070_, _05069_, _05068_);
  and (_05071_, _04718_, \oc8051_golden_model_1.PSW [0]);
  and (_05072_, _04731_, \oc8051_golden_model_1.ACC [0]);
  nor (_05073_, _05072_, _05071_);
  and (_05074_, _05073_, _05070_);
  and (_05075_, _04660_, \oc8051_golden_model_1.P1 [0]);
  not (_05076_, _05075_);
  and (_05077_, _04666_, \oc8051_golden_model_1.P2 [0]);
  and (_05078_, _04670_, \oc8051_golden_model_1.P3 [0]);
  nor (_05079_, _05078_, _05077_);
  and (_05080_, _05079_, _05076_);
  and (_05081_, _05080_, _05074_);
  and (_05082_, _05081_, _05067_);
  and (_05083_, _05082_, _05065_);
  and (_05084_, _05083_, _05059_);
  nand (_05085_, _05084_, _05039_);
  and (_05086_, _05085_, _05038_);
  or (_05087_, _04449_, _02838_);
  and (_05088_, _04638_, \oc8051_golden_model_1.SP [2]);
  not (_05089_, _05088_);
  and (_05090_, _04689_, \oc8051_golden_model_1.TMOD [2]);
  and (_05091_, _04728_, \oc8051_golden_model_1.IE [2]);
  nor (_05092_, _05091_, _05090_);
  and (_05093_, _05092_, _05089_);
  and (_05094_, _04643_, \oc8051_golden_model_1.DPL [2]);
  and (_05095_, _04696_, \oc8051_golden_model_1.DPH [2]);
  nor (_05096_, _05095_, _05094_);
  and (_05097_, _05096_, _05093_);
  and (_05098_, _04648_, \oc8051_golden_model_1.TCON [2]);
  not (_05099_, _05098_);
  and (_05100_, _04701_, \oc8051_golden_model_1.TL0 [2]);
  and (_05101_, _04680_, \oc8051_golden_model_1.TL1 [2]);
  nor (_05102_, _05101_, _05100_);
  and (_05103_, _05102_, _05099_);
  and (_05104_, _04685_, \oc8051_golden_model_1.TH1 [2]);
  and (_05105_, _04691_, \oc8051_golden_model_1.SCON [2]);
  nor (_05106_, _05105_, _05104_);
  and (_05107_, _04704_, \oc8051_golden_model_1.TH0 [2]);
  and (_05108_, _04725_, \oc8051_golden_model_1.SBUF [2]);
  nor (_05109_, _05108_, _05107_);
  and (_05110_, _05109_, _05106_);
  and (_05111_, _05110_, _05103_);
  and (_05112_, _05111_, _05097_);
  and (_05113_, _04718_, \oc8051_golden_model_1.PSW [2]);
  and (_05114_, _04721_, \oc8051_golden_model_1.B [2]);
  nor (_05115_, _05114_, _05113_);
  and (_05116_, _04713_, \oc8051_golden_model_1.IP [2]);
  and (_05117_, _04731_, \oc8051_golden_model_1.ACC [2]);
  nor (_05118_, _05117_, _05116_);
  and (_05119_, _05118_, _05115_);
  and (_05120_, _04710_, \oc8051_golden_model_1.PCON [2]);
  not (_05121_, _05120_);
  and (_05122_, _05121_, _05119_);
  and (_05123_, _04654_, \oc8051_golden_model_1.P0 [2]);
  not (_05124_, _05123_);
  and (_05125_, _04660_, \oc8051_golden_model_1.P1 [2]);
  not (_05126_, _05125_);
  and (_05127_, _04666_, \oc8051_golden_model_1.P2 [2]);
  and (_05128_, _04670_, \oc8051_golden_model_1.P3 [2]);
  nor (_05129_, _05128_, _05127_);
  and (_05130_, _05129_, _05126_);
  and (_05131_, _05130_, _05124_);
  and (_05132_, _05131_, _05122_);
  and (_05133_, _05132_, _05112_);
  and (_05134_, _05133_, _05087_);
  not (_05135_, _05134_);
  and (_05136_, _05135_, _05086_);
  and (_05137_, _05136_, _04993_);
  nand (_05138_, _03785_, \oc8051_golden_model_1.IRAM[0] [4]);
  not (_05139_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05140_, _03785_, _05139_);
  and (_05141_, _05140_, _03780_);
  nand (_05142_, _05141_, _05138_);
  nand (_05143_, _03615_, \oc8051_golden_model_1.IRAM[3] [4]);
  not (_05144_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05145_, _03615_, _05144_);
  and (_05146_, _05145_, _03787_);
  nand (_05147_, _05146_, _05143_);
  nand (_05148_, _05147_, _05142_);
  nand (_05149_, _05148_, _03369_);
  not (_05150_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_05151_, _03785_, _05150_);
  not (_05152_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05153_, _03615_, _05152_);
  and (_05154_, _05153_, _03787_);
  nand (_05155_, _05154_, _05151_);
  not (_05156_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_05157_, _03615_, _05156_);
  not (_05158_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05159_, _03785_, _05158_);
  and (_05160_, _05159_, _03780_);
  nand (_05161_, _05160_, _05157_);
  nand (_05162_, _05161_, _05155_);
  nand (_05163_, _05162_, _03793_);
  nand (_05164_, _05163_, _05149_);
  nand (_05165_, _05164_, _03189_);
  nand (_05166_, _03615_, \oc8051_golden_model_1.IRAM[11] [4]);
  not (_05167_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05168_, _03615_, _05167_);
  and (_05169_, _05168_, _03787_);
  nand (_05170_, _05169_, _05166_);
  nand (_05171_, _03785_, \oc8051_golden_model_1.IRAM[8] [4]);
  not (_05172_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_05173_, _03785_, _05172_);
  and (_05174_, _05173_, _03780_);
  nand (_05175_, _05174_, _05171_);
  nand (_05176_, _05175_, _05170_);
  nand (_05177_, _05176_, _03369_);
  nand (_05178_, _03615_, \oc8051_golden_model_1.IRAM[15] [4]);
  not (_05179_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05180_, _03615_, _05179_);
  and (_05181_, _05180_, _03787_);
  nand (_05182_, _05181_, _05178_);
  nand (_05183_, _03785_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_05184_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_05185_, _03785_, _05184_);
  and (_05186_, _05185_, _03780_);
  nand (_05187_, _05186_, _05183_);
  nand (_05188_, _05187_, _05182_);
  nand (_05189_, _05188_, _03793_);
  nand (_05190_, _05189_, _05177_);
  nand (_05191_, _05190_, _03810_);
  nand (_05192_, _05191_, _05165_);
  or (_05193_, _05192_, _02838_);
  and (_05194_, _04666_, \oc8051_golden_model_1.P2 [4]);
  and (_05195_, _04670_, \oc8051_golden_model_1.P3 [4]);
  nor (_05196_, _05195_, _05194_);
  and (_05197_, _04725_, \oc8051_golden_model_1.SBUF [4]);
  and (_05198_, _04728_, \oc8051_golden_model_1.IE [4]);
  nor (_05199_, _05198_, _05197_);
  and (_05200_, _04709_, _04353_);
  and (_05201_, _05200_, _04634_);
  and (_05202_, _05201_, \oc8051_golden_model_1.PCON [4]);
  not (_05203_, _05202_);
  and (_05204_, _05203_, _05199_);
  and (_05205_, _05204_, _05196_);
  and (_05206_, _04713_, \oc8051_golden_model_1.IP [4]);
  and (_05207_, _04721_, \oc8051_golden_model_1.B [4]);
  nor (_05208_, _05207_, _05206_);
  and (_05209_, _04718_, \oc8051_golden_model_1.PSW [4]);
  and (_05210_, _04731_, \oc8051_golden_model_1.ACC [4]);
  nor (_05211_, _05210_, _05209_);
  and (_05212_, _05211_, _05208_);
  and (_05213_, _04648_, \oc8051_golden_model_1.TCON [4]);
  and (_05214_, _04704_, \oc8051_golden_model_1.TH0 [4]);
  nor (_05215_, _05214_, _05213_);
  and (_05216_, _04660_, \oc8051_golden_model_1.P1 [4]);
  and (_05217_, _04680_, \oc8051_golden_model_1.TL1 [4]);
  nor (_05218_, _05217_, _05216_);
  and (_05219_, _05218_, _05215_);
  and (_05220_, _04691_, \oc8051_golden_model_1.SCON [4]);
  and (_05221_, _04685_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05222_, _05221_, _05220_);
  and (_05223_, _04701_, \oc8051_golden_model_1.TL0 [4]);
  and (_05224_, _04689_, \oc8051_golden_model_1.TMOD [4]);
  nor (_05225_, _05224_, _05223_);
  and (_05226_, _05225_, _05222_);
  and (_05227_, _05226_, _05219_);
  and (_05228_, _05227_, _05212_);
  and (_05229_, _05228_, _05205_);
  and (_05230_, _04654_, \oc8051_golden_model_1.P0 [4]);
  not (_05231_, _05230_);
  and (_05232_, _04638_, \oc8051_golden_model_1.SP [4]);
  and (_05233_, _04643_, \oc8051_golden_model_1.DPL [4]);
  nor (_05234_, _05233_, _05232_);
  nand (_05235_, _04696_, \oc8051_golden_model_1.DPH [4]);
  and (_05236_, _05235_, _05234_);
  and (_05237_, _05236_, _05231_);
  and (_05238_, _05237_, _05229_);
  and (_05239_, _05238_, _05193_);
  not (_05240_, _05239_);
  and (_05241_, _05240_, _05137_);
  and (_05242_, _05241_, _04945_);
  and (_05243_, _05242_, _04838_);
  nor (_05244_, _05243_, _04740_);
  and (_05245_, _05243_, _04740_);
  nor (_05246_, _05245_, _05244_);
  and (_05247_, _05246_, _03943_);
  not (_05248_, _04894_);
  not (_05249_, _05192_);
  nor (_05250_, _04020_, _03872_);
  nor (_05251_, _04449_, _04275_);
  and (_05252_, _05251_, _05250_);
  and (_05253_, _05252_, _05249_);
  and (_05254_, _05253_, _05248_);
  nor (_05255_, _05254_, _04630_);
  and (_05256_, _02855_, _02498_);
  nor (_05257_, _05256_, _03608_);
  nor (_05258_, _04790_, _04630_);
  and (_05259_, _04790_, _04630_);
  nor (_05260_, _05259_, _05258_);
  and (_05261_, _05260_, _05254_);
  or (_05262_, _05261_, _05257_);
  or (_05263_, _05262_, _05255_);
  and (_05264_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_05265_, _05264_, \oc8051_golden_model_1.PC [6]);
  and (_05266_, _05265_, _02638_);
  and (_05267_, _05266_, \oc8051_golden_model_1.PC [7]);
  nor (_05268_, _05266_, \oc8051_golden_model_1.PC [7]);
  nor (_05269_, _05268_, _05267_);
  and (_05270_, _05269_, _02528_);
  and (_05271_, _03022_, _02763_);
  and (_05272_, _03098_, _01165_);
  and (_05273_, _03121_, _01131_);
  nor (_05274_, _05273_, _05272_);
  and (_05275_, _03073_, _01154_);
  and (_05276_, _03095_, _01123_);
  nor (_05277_, _05276_, _05275_);
  and (_05278_, _05277_, _05274_);
  and (_05279_, _03116_, _01146_);
  and (_05280_, _03110_, _01143_);
  nor (_05281_, _05280_, _05279_);
  and (_05282_, _03082_, _01134_);
  and (_05283_, _03076_, _01162_);
  nor (_05284_, _05283_, _05282_);
  and (_05285_, _05284_, _05281_);
  and (_05286_, _05285_, _05278_);
  and (_05287_, _03118_, _01081_);
  and (_05288_, _03123_, _01106_);
  nor (_05289_, _05288_, _05287_);
  and (_05290_, _03100_, _01158_);
  and (_05291_, _03093_, _01151_);
  nor (_05292_, _05291_, _05290_);
  and (_05293_, _05292_, _05289_);
  and (_05294_, _03087_, _01139_);
  and (_05295_, _03112_, _01127_);
  nor (_05296_, _05295_, _05294_);
  and (_05297_, _03105_, _01114_);
  and (_05298_, _03107_, _01118_);
  nor (_05299_, _05298_, _05297_);
  and (_05300_, _05299_, _05296_);
  and (_05301_, _05300_, _05293_);
  and (_05302_, _05301_, _05286_);
  nor (_05303_, _05302_, _04739_);
  and (_05304_, _05303_, _05271_);
  not (_05305_, _02879_);
  not (_05306_, _02927_);
  nor (_05307_, _03648_, _02795_);
  and (_05308_, _05307_, _03222_);
  and (_05309_, _05308_, _05306_);
  and (_05310_, _05309_, _04634_);
  and (_05311_, _05310_, \oc8051_golden_model_1.TCON [7]);
  and (_05312_, _05308_, _02927_);
  and (_05313_, _04730_, _05312_);
  and (_05314_, _05313_, \oc8051_golden_model_1.ACC [7]);
  nor (_05315_, _05314_, _05311_);
  and (_05316_, _04717_, _05312_);
  and (_05317_, _05316_, \oc8051_golden_model_1.PSW [7]);
  not (_05318_, _05317_);
  and (_05319_, _05309_, _04669_);
  and (_05320_, _05319_, \oc8051_golden_model_1.IP [7]);
  and (_05321_, _04720_, _05312_);
  and (_05322_, _05321_, \oc8051_golden_model_1.B [7]);
  nor (_05323_, _05322_, _05320_);
  and (_05324_, _05323_, _05318_);
  and (_05325_, _05324_, _05315_);
  and (_05326_, _05309_, _04659_);
  and (_05327_, _05326_, \oc8051_golden_model_1.SCON [7]);
  and (_05328_, _05309_, _04665_);
  and (_05329_, _05328_, \oc8051_golden_model_1.IE [7]);
  nor (_05330_, _05329_, _05327_);
  and (_05331_, _04635_, \oc8051_golden_model_1.P0 [7]);
  and (_05332_, _04659_, _05312_);
  and (_05333_, _05332_, \oc8051_golden_model_1.P1 [7]);
  nor (_05334_, _05333_, _05331_);
  and (_05335_, _04665_, _05312_);
  and (_05336_, _05335_, \oc8051_golden_model_1.P2 [7]);
  and (_05337_, _04669_, _05312_);
  and (_05338_, _05337_, \oc8051_golden_model_1.P3 [7]);
  nor (_05339_, _05338_, _05336_);
  and (_05340_, _05339_, _05334_);
  and (_05341_, _05340_, _05330_);
  and (_05342_, _05341_, _05325_);
  and (_05343_, _05342_, _04631_);
  nor (_05344_, _05343_, _04709_);
  or (_05345_, _05344_, _05305_);
  not (_05346_, _02886_);
  not (_05347_, _04709_);
  nand (_05348_, _05343_, _05347_);
  or (_05349_, _05348_, _05346_);
  not (_05350_, _04630_);
  and (_05351_, _05192_, _04894_);
  and (_05352_, _04020_, _03872_);
  and (_05353_, _04449_, _04275_);
  and (_05354_, _05353_, _05352_);
  and (_05355_, _05354_, _05351_);
  and (_05356_, _05355_, _04790_);
  or (_05357_, _05356_, _05350_);
  nand (_05358_, _05356_, _05350_);
  and (_05359_, _05358_, _05357_);
  nor (_05360_, _03760_, _03304_);
  and (_05361_, _05360_, _04030_);
  or (_05362_, _05361_, _05359_);
  or (_05363_, _05269_, _02603_);
  not (_05364_, \oc8051_golden_model_1.ACC [7]);
  nand (_05365_, _02603_, _05364_);
  and (_05366_, _05365_, _05363_);
  nor (_05367_, _05366_, _03304_);
  nand (_05368_, _05367_, _04459_);
  and (_05369_, _05368_, _05362_);
  or (_05370_, _05369_, _03840_);
  not (_05371_, _03840_);
  nor (_05372_, _03155_, _02890_);
  nor (_05373_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_05374_, _05373_, _03264_);
  nor (_05375_, _05373_, _03264_);
  nor (_05376_, _05375_, _05374_);
  nor (_05377_, _05376_, _05372_);
  not (_05378_, _05377_);
  not (_05379_, _03889_);
  nand (_05380_, _04449_, _05379_);
  not (_05381_, _05372_);
  and (_05382_, _03889_, _03356_);
  nor (_05383_, _05382_, _05381_);
  nand (_05384_, _05383_, _05380_);
  and (_05385_, _05384_, _05378_);
  or (_05386_, _03889_, _03838_);
  and (_05387_, _03889_, _02837_);
  nor (_05388_, _05387_, _05381_);
  nand (_05389_, _05388_, _05386_);
  nor (_05390_, _05372_, \oc8051_golden_model_1.SP [0]);
  not (_05391_, _05390_);
  and (_05392_, _05391_, _05389_);
  or (_05393_, _05392_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor (_05394_, _05379_, _03687_);
  nor (_05395_, _04020_, _03889_);
  or (_05396_, _05395_, _05394_);
  nand (_05397_, _05396_, _05372_);
  nor (_05398_, _05372_, _03957_);
  not (_05399_, _05398_);
  and (_05400_, _05399_, _05397_);
  nand (_05401_, _05391_, _05389_);
  or (_05402_, _05401_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_05403_, _05402_, _05400_);
  and (_05404_, _05403_, _05393_);
  or (_05405_, _05401_, \oc8051_golden_model_1.IRAM[10] [7]);
  nand (_05406_, _05399_, _05397_);
  or (_05407_, _05392_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_05408_, _05407_, _05406_);
  and (_05409_, _05408_, _05405_);
  nor (_05410_, _05409_, _05404_);
  nand (_05411_, _05410_, _05385_);
  not (_05412_, \oc8051_golden_model_1.SP [3]);
  nor (_05413_, _05374_, _05412_);
  nor (_05414_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05415_, _05414_, _05412_);
  and (_05416_, _05415_, _02868_);
  nor (_05417_, _05416_, _05413_);
  nor (_05418_, _05417_, _05372_);
  not (_05419_, _05418_);
  nand (_05420_, _04275_, _05379_);
  nor (_05421_, _05379_, _02794_);
  nor (_05422_, _05421_, _05381_);
  nand (_05423_, _05422_, _05420_);
  and (_05424_, _05423_, _05419_);
  not (_05425_, _05424_);
  not (_05426_, _05385_);
  or (_05427_, _05392_, _04614_);
  or (_05428_, _05401_, _04616_);
  nand (_05429_, _05428_, _05427_);
  nand (_05430_, _05429_, _05406_);
  or (_05431_, _05392_, _04622_);
  or (_05432_, _05401_, _04620_);
  nand (_05433_, _05432_, _05431_);
  nand (_05434_, _05433_, _05400_);
  and (_05435_, _05434_, _05430_);
  nand (_05436_, _05435_, _05426_);
  and (_05437_, _05436_, _05425_);
  nand (_05438_, _05437_, _05411_);
  or (_05439_, _05392_, _04573_);
  or (_05440_, _05401_, _04571_);
  nand (_05441_, _05440_, _05439_);
  nand (_05442_, _05441_, _05400_);
  or (_05443_, _05392_, _04577_);
  or (_05444_, _05401_, _04579_);
  nand (_05445_, _05444_, _05443_);
  nand (_05446_, _05445_, _05406_);
  nand (_05447_, _05446_, _05442_);
  nand (_05448_, _05447_, _05385_);
  or (_05449_, _05392_, _04594_);
  or (_05450_, _05401_, _04592_);
  nand (_05451_, _05450_, _05449_);
  nand (_05452_, _05451_, _05400_);
  or (_05453_, _05392_, _04586_);
  or (_05454_, _05401_, _04588_);
  nand (_05455_, _05454_, _05453_);
  nand (_05456_, _05455_, _05406_);
  nand (_05457_, _05456_, _05452_);
  nand (_05458_, _05457_, _05426_);
  nand (_05459_, _05458_, _05448_);
  nand (_05460_, _05459_, _05424_);
  nand (_05461_, _05460_, _05438_);
  or (_05462_, _05461_, _05371_);
  and (_05463_, _05462_, _05370_);
  or (_05464_, _05463_, _03843_);
  and (_05465_, _05239_, _04944_);
  not (_05466_, _05085_);
  and (_05467_, _05466_, _05037_);
  and (_05468_, _05134_, _04992_);
  and (_05469_, _05468_, _05467_);
  and (_05470_, _05469_, _05465_);
  and (_05471_, _05470_, _04837_);
  nor (_05472_, _05471_, _04740_);
  and (_05473_, _05471_, _04740_);
  nor (_05474_, _05473_, _05472_);
  or (_05475_, _05474_, _03844_);
  and (_05476_, _05475_, _05464_);
  or (_05477_, _05476_, _02886_);
  and (_05478_, _05477_, _05349_);
  or (_05479_, _05478_, _04225_);
  nor (_05480_, _05269_, _02597_);
  nor (_05481_, _05480_, _03868_);
  and (_05482_, _05481_, _05479_);
  and (_05483_, _05350_, _03868_);
  or (_05484_, _05483_, _02879_);
  or (_05485_, _05484_, _05482_);
  and (_05486_, _05485_, _05345_);
  or (_05487_, _05486_, _02876_);
  and (_05488_, _04666_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05489_, _04670_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05490_, _05489_, _05488_);
  and (_05491_, _04654_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05492_, _04660_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_05493_, _05492_, _05491_);
  and (_05494_, _05493_, _05490_);
  and (_05495_, _05494_, _04651_);
  and (_05496_, _05495_, _04737_);
  and (_05497_, _05496_, _04631_);
  nand (_05498_, _05497_, _02876_);
  and (_05499_, _05498_, _02874_);
  and (_05500_, _05499_, _05487_);
  nor (_05501_, _05343_, _05347_);
  not (_05502_, _05501_);
  and (_05503_, _05502_, _05348_);
  and (_05504_, _05503_, _02873_);
  or (_05505_, _05504_, _05500_);
  and (_05506_, _05505_, _02591_);
  not (_05507_, _05269_);
  or (_05508_, _05507_, _02591_);
  nand (_05509_, _05508_, _02971_);
  or (_05510_, _05509_, _05506_);
  nand (_05511_, _05497_, _03433_);
  and (_05512_, _05511_, _05510_);
  or (_05513_, _05512_, _03889_);
  and (_05514_, _05461_, _02763_);
  nand (_05515_, _05496_, _03889_);
  or (_05516_, _05515_, _05514_);
  and (_05517_, _05516_, _04325_);
  and (_05518_, _05517_, _05513_);
  and (_05519_, _04635_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05520_, _05335_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_05521_, _05520_, _05519_);
  and (_05522_, _05332_, \oc8051_golden_model_1.P1INREG [7]);
  and (_05523_, _05337_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05524_, _05523_, _05522_);
  and (_05525_, _05524_, _05521_);
  and (_05526_, _05525_, _05330_);
  and (_05527_, _05526_, _05325_);
  and (_05528_, _05527_, _04631_);
  nor (_05529_, _05528_, _04709_);
  and (_05530_, _04709_, \oc8051_golden_model_1.PSW [7]);
  nor (_05531_, _05530_, _05529_);
  nor (_05532_, _05531_, _04325_);
  or (_05533_, _05532_, _02569_);
  or (_05534_, _05533_, _05518_);
  not (_05535_, _02859_);
  and (_05536_, _05535_, _02763_);
  and (_05537_, _05507_, _02569_);
  nor (_05538_, _05537_, _05536_);
  and (_05539_, _05538_, _05534_);
  and (_05540_, _02841_, _02763_);
  not (_05541_, _05536_);
  nor (_05542_, _04630_, _05541_);
  or (_05543_, _05542_, _05540_);
  or (_05544_, _05543_, _05539_);
  not (_05545_, _05540_);
  or (_05546_, _05461_, _05545_);
  and (_05547_, _05546_, _04193_);
  and (_05548_, _05547_, _05544_);
  not (_05549_, _05302_);
  nor (_05550_, _05549_, _04630_);
  not (_05551_, _05550_);
  and (_05552_, _03262_, _03128_);
  and (_05553_, _03720_, _03505_);
  and (_05554_, _05553_, _05552_);
  and (_05555_, _03076_, _01578_);
  and (_05556_, _03112_, _01541_);
  nor (_05557_, _05556_, _05555_);
  and (_05558_, _03118_, _01546_);
  and (_05559_, _03123_, _01555_);
  nor (_05560_, _05559_, _05558_);
  and (_05561_, _05560_, _05557_);
  and (_05562_, _03107_, _01552_);
  and (_05563_, _03116_, _01561_);
  nor (_05564_, _05563_, _05562_);
  and (_05565_, _03073_, _01571_);
  and (_05566_, _03105_, _01550_);
  nor (_05567_, _05566_, _05565_);
  and (_05568_, _05567_, _05564_);
  and (_05569_, _05568_, _05561_);
  and (_05570_, _03110_, _01563_);
  and (_05571_, _03093_, _01557_);
  nor (_05572_, _05571_, _05570_);
  and (_05573_, _03098_, _01573_);
  and (_05574_, _03121_, _01539_);
  nor (_05575_, _05574_, _05573_);
  and (_05576_, _05575_, _05572_);
  and (_05577_, _03087_, _01566_);
  and (_05578_, _03100_, _01576_);
  nor (_05579_, _05578_, _05577_);
  and (_05580_, _03082_, _01569_);
  and (_05581_, _03095_, _01544_);
  nor (_05582_, _05581_, _05580_);
  and (_05583_, _05582_, _05579_);
  and (_05584_, _05583_, _05576_);
  and (_05585_, _05584_, _05569_);
  and (_05586_, _05585_, _05549_);
  and (_05587_, _03087_, _01474_);
  and (_05588_, _03118_, _01463_);
  nor (_05589_, _05588_, _05587_);
  and (_05590_, _03073_, _01484_);
  and (_05591_, _03100_, _01481_);
  nor (_05592_, _05591_, _05590_);
  and (_05593_, _05592_, _05589_);
  and (_05594_, _03110_, _01469_);
  and (_05595_, _03093_, _01449_);
  nor (_05596_, _05595_, _05594_);
  and (_05597_, _03121_, _01454_);
  and (_05598_, _03123_, _01477_);
  nor (_05599_, _05598_, _05597_);
  and (_05600_, _05599_, _05596_);
  and (_05601_, _05600_, _05593_);
  and (_05602_, _03105_, _01447_);
  and (_05603_, _03116_, _01471_);
  nor (_05604_, _05603_, _05602_);
  and (_05605_, _03095_, _01452_);
  and (_05606_, _03112_, _01465_);
  nor (_05607_, _05606_, _05605_);
  and (_05608_, _05607_, _05604_);
  and (_05609_, _03098_, _01479_);
  and (_05610_, _03107_, _01460_);
  nor (_05611_, _05610_, _05609_);
  and (_05612_, _03082_, _01458_);
  and (_05613_, _03076_, _01486_);
  nor (_05614_, _05613_, _05612_);
  and (_05615_, _05614_, _05611_);
  and (_05616_, _05615_, _05608_);
  and (_05617_, _05616_, _05601_);
  not (_05618_, _05617_);
  and (_05619_, _03073_, _01525_);
  and (_05620_, _03118_, _01493_);
  nor (_05621_, _05620_, _05619_);
  and (_05622_, _03105_, _01523_);
  and (_05623_, _03110_, _01517_);
  nor (_05624_, _05623_, _05622_);
  and (_05625_, _05624_, _05621_);
  and (_05626_, _03123_, _01511_);
  and (_05627_, _03112_, _01495_);
  nor (_05628_, _05627_, _05626_);
  and (_05629_, _03098_, _01527_);
  and (_05630_, _03076_, _01530_);
  nor (_05631_, _05630_, _05629_);
  and (_05632_, _05631_, _05628_);
  and (_05633_, _05632_, _05625_);
  and (_05634_, _03100_, _01532_);
  and (_05635_, _03087_, _01515_);
  nor (_05636_, _05635_, _05634_);
  and (_05637_, _03082_, _01500_);
  and (_05638_, _03107_, _01506_);
  nor (_05639_, _05638_, _05637_);
  and (_05640_, _05639_, _05636_);
  and (_05641_, _03116_, _01519_);
  and (_05642_, _03095_, _01504_);
  nor (_05643_, _05642_, _05641_);
  and (_05644_, _03093_, _01509_);
  and (_05645_, _03121_, _01498_);
  nor (_05646_, _05645_, _05644_);
  and (_05647_, _05646_, _05643_);
  and (_05648_, _05647_, _05640_);
  and (_05649_, _05648_, _05633_);
  and (_05650_, _05649_, _05618_);
  and (_05651_, _05650_, _05586_);
  and (_05652_, _05651_, _05554_);
  and (_05653_, _05652_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05654_, _03128_);
  and (_05655_, _03262_, _05654_);
  and (_05656_, _05655_, _05553_);
  and (_05657_, _05656_, _05651_);
  and (_05658_, _05657_, \oc8051_golden_model_1.SCON [7]);
  nor (_05659_, _05658_, _05653_);
  not (_05660_, _03505_);
  and (_05661_, _03720_, _05660_);
  and (_05662_, _05661_, _05655_);
  and (_05663_, _05662_, _05651_);
  and (_05664_, _05663_, \oc8051_golden_model_1.SBUF [7]);
  nor (_05665_, _05585_, _05302_);
  and (_05666_, _05665_, _05554_);
  and (_05667_, _05666_, _05650_);
  and (_05668_, _05667_, \oc8051_golden_model_1.PSW [7]);
  nor (_05669_, _05668_, _05664_);
  and (_05670_, _05669_, _05659_);
  not (_05671_, _05649_);
  and (_05672_, _05671_, _05617_);
  and (_05673_, _05672_, _05666_);
  and (_05674_, _05673_, \oc8051_golden_model_1.ACC [7]);
  nor (_05675_, _05649_, _05617_);
  and (_05676_, _05675_, _05666_);
  and (_05677_, _05676_, \oc8051_golden_model_1.B [7]);
  nor (_05678_, _05677_, _05674_);
  and (_05679_, _05649_, _05617_);
  and (_05680_, _05679_, _05586_);
  and (_05681_, _05680_, _05554_);
  and (_05682_, _05681_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05683_, _05680_, _05656_);
  and (_05684_, _05683_, \oc8051_golden_model_1.TCON [7]);
  nor (_05685_, _05684_, _05682_);
  and (_05686_, _05685_, _05678_);
  and (_05687_, _05686_, _05670_);
  nor (_05688_, _03720_, _03505_);
  and (_05689_, _05688_, _05680_);
  and (_05690_, _05689_, _03128_);
  and (_05691_, _05690_, _03262_);
  and (_05692_, _05691_, \oc8051_golden_model_1.DPH [7]);
  not (_05693_, _03262_);
  and (_05694_, _05690_, _05693_);
  and (_05695_, _05694_, \oc8051_golden_model_1.PCON [7]);
  nor (_05696_, _05695_, _05692_);
  and (_05697_, _05696_, _05687_);
  nor (_05698_, _03262_, _03128_);
  and (_05699_, _05698_, _05680_);
  and (_05700_, _05699_, _05553_);
  and (_05701_, _05700_, \oc8051_golden_model_1.TH0 [7]);
  and (_05702_, _05680_, _05655_);
  not (_05703_, _03720_);
  and (_05704_, _05703_, _03505_);
  and (_05705_, _05704_, _05702_);
  and (_05706_, _05705_, \oc8051_golden_model_1.TL0 [7]);
  nor (_05707_, _05706_, _05701_);
  and (_05708_, _05680_, _05552_);
  and (_05709_, _05708_, _05661_);
  and (_05710_, _05709_, \oc8051_golden_model_1.SP [7]);
  and (_05711_, _05708_, _05704_);
  and (_05712_, _05711_, \oc8051_golden_model_1.DPL [7]);
  nor (_05713_, _05712_, _05710_);
  and (_05714_, _05713_, _05707_);
  and (_05715_, _05689_, _05655_);
  and (_05716_, _05715_, \oc8051_golden_model_1.TL1 [7]);
  and (_05717_, _05699_, _05661_);
  and (_05718_, _05717_, \oc8051_golden_model_1.TH1 [7]);
  nor (_05719_, _05718_, _05716_);
  and (_05720_, _05702_, _05661_);
  and (_05721_, _05720_, \oc8051_golden_model_1.TMOD [7]);
  not (_05722_, _05721_);
  and (_05723_, _05672_, _05586_);
  and (_05724_, _05723_, _05554_);
  and (_05725_, _05724_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05726_, _05675_, _05586_);
  and (_05727_, _05726_, _05554_);
  and (_05728_, _05727_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05729_, _05728_, _05725_);
  and (_05730_, _05723_, _05656_);
  and (_05731_, _05730_, \oc8051_golden_model_1.IE [7]);
  and (_05732_, _05726_, _05656_);
  and (_05733_, _05732_, \oc8051_golden_model_1.IP [7]);
  nor (_05734_, _05733_, _05731_);
  and (_05735_, _05734_, _05729_);
  and (_05736_, _05735_, _05722_);
  and (_05737_, _05736_, _05719_);
  and (_05738_, _05737_, _05714_);
  and (_05739_, _05738_, _05697_);
  and (_05740_, _05739_, _05551_);
  nor (_05741_, _05740_, _04193_);
  not (_05742_, _03510_);
  and (_05743_, _03901_, _04138_);
  not (_05744_, _05743_);
  and (_05745_, _05744_, _04164_);
  and (_05746_, _05745_, _04169_);
  and (_05747_, _05746_, _04172_);
  and (_05748_, _05747_, _05742_);
  not (_05749_, _05748_);
  or (_05750_, _05749_, _05741_);
  or (_05751_, _05750_, _05548_);
  and (_05752_, _05749_, _02763_);
  nor (_05753_, _05752_, _02835_);
  and (_05754_, _05753_, _05751_);
  and (_05755_, _05549_, _02835_);
  or (_05756_, _05755_, _02522_);
  or (_05757_, _05756_, _05754_);
  and (_05758_, _03051_, _02763_);
  and (_05759_, _05507_, _02522_);
  nor (_05760_, _05759_, _05758_);
  and (_05761_, _05760_, _05757_);
  and (_05762_, _03148_, _02763_);
  and (_05763_, _05302_, _04739_);
  nor (_05764_, _05763_, _05303_);
  and (_05765_, _05764_, _05758_);
  or (_05766_, _05765_, _05762_);
  or (_05767_, _05766_, _05761_);
  not (_05768_, _05271_);
  not (_05769_, _05762_);
  nor (_05770_, _04739_, _05364_);
  and (_05771_, _04739_, _05364_);
  nor (_05772_, _05771_, _05770_);
  or (_05773_, _05772_, _05769_);
  and (_05774_, _05773_, _05768_);
  and (_05775_, _05774_, _05767_);
  or (_05776_, _05775_, _05304_);
  and (_05777_, _05776_, _04129_);
  and (_05778_, _05770_, _03909_);
  or (_05779_, _05778_, _02530_);
  or (_05780_, _05779_, _05777_);
  and (_05781_, _03042_, _02763_);
  and (_05782_, _05507_, _02530_);
  nor (_05783_, _05782_, _05781_);
  and (_05784_, _05783_, _05780_);
  and (_05785_, _03143_, _02763_);
  not (_05786_, _05781_);
  nor (_05787_, _05763_, _05786_);
  or (_05788_, _05787_, _05785_);
  or (_05789_, _05788_, _05784_);
  not (_05790_, _02528_);
  nand (_05791_, _05771_, _05785_);
  and (_05792_, _05791_, _05790_);
  and (_05793_, _05792_, _05789_);
  nor (_05794_, _05793_, _05270_);
  nor (_05795_, _05794_, _03299_);
  not (_05796_, _04104_);
  and (_05797_, _04130_, _05796_);
  nand (_05798_, _05359_, _03299_);
  nand (_05799_, _05798_, _05797_);
  or (_05800_, _05799_, _05795_);
  not (_05801_, _03587_);
  or (_05802_, _05797_, _05359_);
  and (_05803_, _05802_, _05801_);
  and (_05804_, _05803_, _05800_);
  and (_05805_, _05359_, _03587_);
  or (_05806_, _05805_, _03927_);
  or (_05807_, _05806_, _05804_);
  not (_05808_, _03929_);
  not (_05809_, _03927_);
  and (_05810_, _05460_, _05438_);
  or (_05811_, _05392_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_05812_, _05401_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_05813_, _05812_, _05400_);
  and (_05814_, _05813_, _05811_);
  or (_05815_, _05401_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_05816_, _05392_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_05817_, _05816_, _05406_);
  and (_05818_, _05817_, _05815_);
  nor (_05819_, _05818_, _05814_);
  nand (_05820_, _05819_, _05385_);
  or (_05821_, _05392_, _04751_);
  or (_05822_, _05401_, _04753_);
  nand (_05823_, _05822_, _05821_);
  nand (_05824_, _05823_, _05406_);
  or (_05825_, _05392_, _04759_);
  or (_05826_, _05401_, _04757_);
  nand (_05827_, _05826_, _05825_);
  nand (_05828_, _05827_, _05400_);
  and (_05829_, _05828_, _05824_);
  nand (_05830_, _05829_, _05426_);
  and (_05831_, _05830_, _05424_);
  nand (_05832_, _05831_, _05820_);
  or (_05833_, _05401_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_05834_, _05392_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_05835_, _05834_, _05833_);
  nand (_05836_, _05835_, _05400_);
  or (_05837_, _05401_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_05838_, _05392_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_05839_, _05838_, _05837_);
  nand (_05840_, _05839_, _05406_);
  nand (_05841_, _05840_, _05836_);
  nand (_05842_, _05841_, _05426_);
  or (_05843_, _05401_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_05844_, _05392_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_05845_, _05844_, _05843_);
  nand (_05846_, _05845_, _05400_);
  or (_05847_, _05401_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_05848_, _05392_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_05849_, _05848_, _05847_);
  nand (_05850_, _05849_, _05406_);
  nand (_05851_, _05850_, _05846_);
  nand (_05852_, _05851_, _05385_);
  and (_05853_, _05852_, _05425_);
  nand (_05854_, _05853_, _05842_);
  and (_05855_, _05854_, _05832_);
  or (_05856_, _05392_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_05857_, _05401_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_05858_, _05857_, _05400_);
  and (_05859_, _05858_, _05856_);
  or (_05860_, _05401_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_05861_, _05392_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_05862_, _05861_, _05406_);
  and (_05863_, _05862_, _05860_);
  nor (_05864_, _05863_, _05859_);
  nand (_05865_, _05864_, _05385_);
  or (_05866_, _05392_, _03978_);
  or (_05867_, _05401_, _03980_);
  nand (_05868_, _05867_, _05866_);
  nand (_05869_, _05868_, _05406_);
  or (_05870_, _05392_, _03986_);
  or (_05871_, _05401_, _03984_);
  nand (_05872_, _05871_, _05870_);
  nand (_05873_, _05872_, _05400_);
  and (_05874_, _05873_, _05869_);
  nand (_05875_, _05874_, _05426_);
  and (_05876_, _05875_, _05424_);
  nand (_05877_, _05876_, _05865_);
  or (_05878_, _05401_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_05879_, _05392_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_05880_, _05879_, _05878_);
  nand (_05881_, _05880_, _05400_);
  or (_05882_, _05401_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_05883_, _05392_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_05884_, _05883_, _05882_);
  nand (_05885_, _05884_, _05406_);
  nand (_05886_, _05885_, _05881_);
  nand (_05887_, _05886_, _05426_);
  or (_05888_, _05401_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_05889_, _05392_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_05890_, _05889_, _05888_);
  nand (_05891_, _05890_, _05400_);
  or (_05892_, _05401_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_05893_, _05392_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_05894_, _05893_, _05892_);
  nand (_05895_, _05894_, _05406_);
  nand (_05896_, _05895_, _05891_);
  nand (_05897_, _05896_, _05385_);
  and (_05898_, _05897_, _05425_);
  nand (_05899_, _05898_, _05887_);
  and (_05900_, _05899_, _05877_);
  or (_05901_, _05392_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_05902_, _05401_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_05903_, _05902_, _05400_);
  and (_05904_, _05903_, _05901_);
  or (_05905_, _05401_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_05906_, _05392_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_05907_, _05906_, _05406_);
  and (_05908_, _05907_, _05905_);
  nor (_05909_, _05908_, _05904_);
  nand (_05910_, _05909_, _05385_);
  or (_05911_, _05392_, _03794_);
  or (_05912_, _05401_, _03796_);
  nand (_05913_, _05912_, _05911_);
  nand (_05914_, _05913_, _05406_);
  or (_05915_, _05392_, _03802_);
  or (_05916_, _05401_, _03800_);
  nand (_05917_, _05916_, _05915_);
  nand (_05918_, _05917_, _05400_);
  and (_05919_, _05918_, _05914_);
  nand (_05920_, _05919_, _05426_);
  and (_05921_, _05920_, _05424_);
  nand (_05922_, _05921_, _05910_);
  or (_05923_, _05401_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_05924_, _05392_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_05925_, _05924_, _05923_);
  nand (_05926_, _05925_, _05400_);
  or (_05927_, _05401_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_05928_, _05392_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_05929_, _05928_, _05927_);
  nand (_05930_, _05929_, _05406_);
  nand (_05931_, _05930_, _05926_);
  nand (_05932_, _05931_, _05426_);
  or (_05933_, _05401_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_05934_, _05392_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_05935_, _05934_, _05933_);
  nand (_05936_, _05935_, _05400_);
  or (_05937_, _05401_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_05938_, _05392_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_05939_, _05938_, _05937_);
  nand (_05940_, _05939_, _05406_);
  nand (_05941_, _05940_, _05936_);
  nand (_05942_, _05941_, _05385_);
  and (_05943_, _05942_, _05425_);
  nand (_05944_, _05943_, _05932_);
  and (_05945_, _05944_, _05922_);
  and (_05946_, _05945_, _05900_);
  or (_05947_, _05392_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_05948_, _05401_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_05949_, _05948_, _05400_);
  and (_05950_, _05949_, _05947_);
  or (_05951_, _05401_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_05952_, _05392_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_05953_, _05952_, _05406_);
  and (_05954_, _05953_, _05951_);
  nor (_05955_, _05954_, _05950_);
  nand (_05956_, _05955_, _05385_);
  or (_05957_, _05392_, _04237_);
  or (_05958_, _05401_, _04239_);
  nand (_05959_, _05958_, _05957_);
  nand (_05960_, _05959_, _05406_);
  or (_05961_, _05392_, _04245_);
  or (_05962_, _05401_, _04243_);
  nand (_05963_, _05962_, _05961_);
  nand (_05964_, _05963_, _05400_);
  and (_05965_, _05964_, _05960_);
  nand (_05966_, _05965_, _05426_);
  and (_05967_, _05966_, _05424_);
  nand (_05968_, _05967_, _05956_);
  or (_05969_, _05401_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_05970_, _05392_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_05971_, _05970_, _05969_);
  nand (_05972_, _05971_, _05400_);
  or (_05973_, _05401_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_05974_, _05392_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_05975_, _05974_, _05973_);
  nand (_05976_, _05975_, _05406_);
  nand (_05977_, _05976_, _05972_);
  nand (_05978_, _05977_, _05426_);
  or (_05979_, _05401_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_05980_, _05392_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_05981_, _05980_, _05979_);
  nand (_05982_, _05981_, _05400_);
  or (_05983_, _05401_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_05984_, _05392_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_05985_, _05984_, _05983_);
  nand (_05986_, _05985_, _05406_);
  nand (_05987_, _05986_, _05982_);
  nand (_05988_, _05987_, _05385_);
  and (_05989_, _05988_, _05425_);
  nand (_05990_, _05989_, _05978_);
  and (_05991_, _05990_, _05968_);
  or (_05992_, _05392_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_05993_, _05401_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_05994_, _05993_, _05400_);
  and (_05995_, _05994_, _05992_);
  or (_05996_, _05401_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_05997_, _05392_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_05998_, _05997_, _05406_);
  and (_05999_, _05998_, _05996_);
  nor (_06000_, _05999_, _05995_);
  nand (_06001_, _06000_, _05385_);
  or (_06002_, _05392_, _04407_);
  or (_06003_, _05401_, _04409_);
  nand (_06004_, _06003_, _06002_);
  nand (_06005_, _06004_, _05406_);
  or (_06006_, _05392_, _04415_);
  or (_06007_, _05401_, _04413_);
  nand (_06008_, _06007_, _06006_);
  nand (_06009_, _06008_, _05400_);
  and (_06010_, _06009_, _06005_);
  nand (_06011_, _06010_, _05426_);
  and (_06012_, _06011_, _05424_);
  nand (_06013_, _06012_, _06001_);
  or (_06014_, _05401_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_06015_, _05392_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_06016_, _06015_, _06014_);
  nand (_06017_, _06016_, _05400_);
  or (_06018_, _05401_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_06019_, _05392_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_06020_, _06019_, _06018_);
  nand (_06021_, _06020_, _05406_);
  nand (_06022_, _06021_, _06017_);
  nand (_06023_, _06022_, _05426_);
  or (_06024_, _05401_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_06025_, _05392_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_06026_, _06025_, _06024_);
  nand (_06027_, _06026_, _05400_);
  or (_06028_, _05401_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_06029_, _05392_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_06030_, _06029_, _06028_);
  nand (_06031_, _06030_, _05406_);
  nand (_06032_, _06031_, _06027_);
  nand (_06033_, _06032_, _05385_);
  and (_06034_, _06033_, _05425_);
  nand (_06035_, _06034_, _06023_);
  and (_06036_, _06035_, _06013_);
  and (_06037_, _06036_, _05991_);
  and (_06038_, _06037_, _05946_);
  or (_06039_, _05392_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_06040_, _05401_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_06041_, _06040_, _05400_);
  and (_06042_, _06041_, _06039_);
  or (_06043_, _05401_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_06044_, _05392_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_06045_, _06044_, _05406_);
  and (_06046_, _06045_, _06043_);
  nor (_06047_, _06046_, _06042_);
  nand (_06048_, _06047_, _05385_);
  or (_06049_, _05392_, _04851_);
  or (_06050_, _05401_, _04853_);
  nand (_06051_, _06050_, _06049_);
  nand (_06052_, _06051_, _05406_);
  or (_06053_, _05392_, _04859_);
  or (_06054_, _05401_, _04857_);
  nand (_06055_, _06054_, _06053_);
  nand (_06056_, _06055_, _05400_);
  and (_06057_, _06056_, _06052_);
  nand (_06058_, _06057_, _05426_);
  and (_06059_, _06058_, _05424_);
  nand (_06060_, _06059_, _06048_);
  or (_06061_, _05401_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_06062_, _05392_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_06063_, _06062_, _06061_);
  nand (_06064_, _06063_, _05400_);
  or (_06065_, _05401_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06066_, _05392_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_06067_, _06066_, _06065_);
  nand (_06068_, _06067_, _05406_);
  nand (_06069_, _06068_, _06064_);
  nand (_06070_, _06069_, _05426_);
  or (_06071_, _05401_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_06072_, _05392_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_06073_, _06072_, _06071_);
  nand (_06074_, _06073_, _05400_);
  or (_06075_, _05401_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06076_, _05392_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_06077_, _06076_, _06075_);
  nand (_06078_, _06077_, _05406_);
  nand (_06079_, _06078_, _06074_);
  nand (_06080_, _06079_, _05385_);
  and (_06081_, _06080_, _05425_);
  nand (_06082_, _06081_, _06070_);
  and (_06083_, _06082_, _06060_);
  or (_06084_, _05392_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_06085_, _05401_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_06086_, _06085_, _05400_);
  and (_06087_, _06086_, _06084_);
  or (_06088_, _05401_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_06089_, _05392_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_06090_, _06089_, _05406_);
  and (_06091_, _06090_, _06088_);
  nor (_06092_, _06091_, _06087_);
  nand (_06093_, _06092_, _05385_);
  or (_06094_, _05392_, _05150_);
  or (_06095_, _05401_, _05152_);
  nand (_06096_, _06095_, _06094_);
  nand (_06097_, _06096_, _05406_);
  or (_06098_, _05392_, _05158_);
  or (_06099_, _05401_, _05156_);
  nand (_06100_, _06099_, _06098_);
  nand (_06101_, _06100_, _05400_);
  and (_06102_, _06101_, _06097_);
  nand (_06103_, _06102_, _05426_);
  and (_06104_, _06103_, _05424_);
  nand (_06105_, _06104_, _06093_);
  or (_06106_, _05401_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_06107_, _05392_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_06108_, _06107_, _06106_);
  nand (_06109_, _06108_, _05400_);
  or (_06110_, _05401_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06111_, _05392_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_06112_, _06111_, _06110_);
  nand (_06113_, _06112_, _05406_);
  nand (_06114_, _06113_, _06109_);
  nand (_06115_, _06114_, _05426_);
  or (_06116_, _05401_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_06117_, _05392_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_06118_, _06117_, _06116_);
  nand (_06119_, _06118_, _05400_);
  or (_06120_, _05401_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06121_, _05392_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_06122_, _06121_, _06120_);
  nand (_06123_, _06122_, _05406_);
  nand (_06124_, _06123_, _06119_);
  nand (_06125_, _06124_, _05385_);
  and (_06126_, _06125_, _05425_);
  nand (_06127_, _06126_, _06115_);
  and (_06128_, _06127_, _06105_);
  and (_06129_, _06128_, _06083_);
  and (_06130_, _06129_, _06038_);
  and (_06131_, _06130_, _05855_);
  and (_06132_, _06131_, _05810_);
  nor (_06133_, _06131_, _05810_);
  or (_06134_, _06133_, _06132_);
  or (_06135_, _06134_, _05809_);
  and (_06136_, _06135_, _05808_);
  and (_06137_, _06136_, _05807_);
  and (_06138_, _05474_, _03929_);
  or (_06139_, _06138_, _03034_);
  or (_06140_, _06139_, _06137_);
  and (_06141_, _02251_, \oc8051_golden_model_1.PC [2]);
  and (_06142_, _06141_, \oc8051_golden_model_1.PC [3]);
  and (_06143_, _06142_, _05265_);
  and (_06144_, _06143_, \oc8051_golden_model_1.PC [7]);
  nor (_06145_, _06143_, \oc8051_golden_model_1.PC [7]);
  nor (_06146_, _06145_, _06144_);
  not (_06147_, _06146_);
  nand (_06148_, _06147_, _03034_);
  and (_06149_, _06148_, _06140_);
  or (_06150_, _06149_, _02505_);
  and (_06151_, _05507_, _02505_);
  nor (_06152_, _06151_, _02801_);
  and (_06153_, _06152_, _06150_);
  not (_06154_, _05257_);
  and (_06155_, _05529_, _02801_);
  or (_06156_, _06155_, _06154_);
  or (_06157_, _06156_, _06153_);
  and (_06158_, _06157_, _05263_);
  or (_06159_, _06158_, _03941_);
  not (_06160_, _03943_);
  not (_06161_, _03941_);
  nand (_06162_, _05854_, _05832_);
  nand (_06163_, _05899_, _05877_);
  nand (_06164_, _05944_, _05922_);
  and (_06165_, _06164_, _06163_);
  nand (_06166_, _05990_, _05968_);
  nand (_06167_, _06035_, _06013_);
  and (_06168_, _06167_, _06166_);
  and (_06169_, _06168_, _06165_);
  nand (_06170_, _06082_, _06060_);
  nand (_06171_, _06127_, _06105_);
  and (_06172_, _06171_, _06170_);
  and (_06173_, _06172_, _06169_);
  and (_06174_, _06173_, _06162_);
  nand (_06175_, _06174_, _05461_);
  or (_06176_, _06174_, _05461_);
  and (_06177_, _06176_, _06175_);
  or (_06178_, _06177_, _06161_);
  and (_06179_, _06178_, _06160_);
  and (_06180_, _06179_, _06159_);
  or (_06181_, _06180_, _05247_);
  and (_06182_, _06181_, _04562_);
  or (_06183_, _06182_, _04570_);
  and (_06184_, _06183_, _04560_);
  not (_06185_, _03034_);
  and (_06186_, _06144_, \oc8051_golden_model_1.PC [8]);
  and (_06187_, _06186_, \oc8051_golden_model_1.PC [9]);
  and (_06188_, _06187_, \oc8051_golden_model_1.PC [10]);
  and (_06189_, _06188_, \oc8051_golden_model_1.PC [11]);
  and (_06190_, _06189_, \oc8051_golden_model_1.PC [12]);
  and (_06191_, _06190_, \oc8051_golden_model_1.PC [13]);
  and (_06192_, _06191_, \oc8051_golden_model_1.PC [14]);
  nor (_06193_, _06192_, \oc8051_golden_model_1.PC [15]);
  and (_06194_, _06192_, \oc8051_golden_model_1.PC [15]);
  nor (_06195_, _06194_, _06193_);
  or (_06196_, _06195_, _06185_);
  and (_06197_, _05267_, \oc8051_golden_model_1.PC [8]);
  and (_06198_, _06197_, \oc8051_golden_model_1.PC [9]);
  and (_06199_, _06198_, \oc8051_golden_model_1.PC [10]);
  and (_06200_, _06199_, \oc8051_golden_model_1.PC [11]);
  and (_06201_, _06200_, \oc8051_golden_model_1.PC [12]);
  and (_06202_, _06201_, \oc8051_golden_model_1.PC [13]);
  and (_06203_, _06202_, \oc8051_golden_model_1.PC [14]);
  nor (_06204_, _06203_, \oc8051_golden_model_1.PC [15]);
  and (_06205_, _06203_, \oc8051_golden_model_1.PC [15]);
  nor (_06206_, _06205_, _06204_);
  or (_06207_, _06206_, _03034_);
  and (_06208_, _06207_, _06196_);
  and (_06209_, _06208_, _04555_);
  and (_06210_, _06209_, _04558_);
  or (_35910_, _06210_, _06184_);
  not (_06211_, \oc8051_golden_model_1.B [7]);
  nor (_06212_, _34655_, _06211_);
  not (_06213_, _03137_);
  nor (_06214_, _04721_, _06211_);
  or (_06215_, _06214_, _04740_);
  and (_06216_, _05549_, _04721_);
  or (_06217_, _06216_, _06214_);
  and (_06218_, _06217_, _03022_);
  and (_06219_, _06218_, _06215_);
  not (_06220_, _04721_);
  nor (_06221_, _06220_, _04630_);
  or (_06222_, _06221_, _06214_);
  or (_06223_, _06222_, _02859_);
  and (_06224_, _05474_, _04721_);
  or (_06225_, _06224_, _06214_);
  or (_06226_, _06225_, _03006_);
  and (_06227_, _04721_, \oc8051_golden_model_1.ACC [7]);
  or (_06228_, _06227_, _06214_);
  and (_06229_, _06228_, _03845_);
  nor (_06230_, _03845_, _06211_);
  or (_06231_, _06230_, _02948_);
  or (_06232_, _06231_, _06229_);
  and (_06233_, _06232_, _02976_);
  and (_06234_, _06233_, _06226_);
  and (_06235_, _06222_, _02946_);
  nor (_06236_, _05321_, _06211_);
  and (_06237_, _05348_, _05321_);
  or (_06238_, _06237_, _06236_);
  and (_06239_, _06238_, _02884_);
  or (_06240_, _06239_, _06235_);
  or (_06241_, _06240_, _02880_);
  or (_06242_, _06241_, _06234_);
  or (_06243_, _06228_, _02992_);
  and (_06244_, _06243_, _06242_);
  or (_06245_, _06244_, _02877_);
  not (_06246_, _02871_);
  and (_06247_, _05344_, _05321_);
  or (_06248_, _06247_, _06236_);
  or (_06249_, _06248_, _02987_);
  and (_06250_, _06249_, _06246_);
  and (_06251_, _06250_, _06245_);
  and (_06252_, _03028_, _02939_);
  or (_06253_, _06236_, _05502_);
  and (_06254_, _06253_, _02871_);
  and (_06255_, _06254_, _06238_);
  or (_06256_, _06255_, _06252_);
  or (_06257_, _06256_, _06251_);
  not (_06258_, _06252_);
  and (_06259_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_06260_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_06261_, _06260_, _06259_);
  and (_06262_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_06263_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_06264_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_06265_, _06264_, _06263_);
  nor (_06266_, _06265_, _06261_);
  and (_06267_, _06266_, _06262_);
  nor (_06268_, _06267_, _06261_);
  and (_06269_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_06270_, _06269_, _06264_);
  and (_06271_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_06272_, _06271_, _06259_);
  nor (_06273_, _06272_, _06270_);
  not (_06274_, _06273_);
  nor (_06275_, _06274_, _06268_);
  and (_06276_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_06277_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_06278_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_06279_, _06278_, _06277_);
  nor (_06280_, _06278_, _06277_);
  nor (_06281_, _06280_, _06279_);
  and (_06282_, _06281_, _06276_);
  nor (_06283_, _06281_, _06276_);
  nor (_06284_, _06283_, _06282_);
  and (_06285_, _06274_, _06268_);
  nor (_06286_, _06285_, _06275_);
  and (_06287_, _06286_, _06284_);
  nor (_06288_, _06287_, _06275_);
  not (_06289_, _06264_);
  and (_06290_, _06269_, _06289_);
  and (_06291_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_06292_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_06293_, _06292_, _06277_);
  and (_06294_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_06295_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_06296_, _06295_, _06294_);
  nor (_06297_, _06296_, _06293_);
  and (_06298_, _06297_, _06291_);
  nor (_06299_, _06297_, _06291_);
  nor (_06300_, _06299_, _06298_);
  and (_06301_, _06300_, _06290_);
  nor (_06302_, _06300_, _06290_);
  nor (_06303_, _06302_, _06301_);
  not (_06304_, _06303_);
  nor (_06305_, _06304_, _06288_);
  and (_06306_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_06307_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_06308_, _06307_, _06306_);
  nor (_06309_, _06282_, _06279_);
  and (_06310_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_06311_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_06312_, _06311_, _06310_);
  nor (_06313_, _06311_, _06310_);
  nor (_06314_, _06313_, _06312_);
  not (_06315_, _06314_);
  nor (_06316_, _06315_, _06309_);
  and (_06317_, _06315_, _06309_);
  nor (_06318_, _06317_, _06316_);
  and (_06319_, _06318_, _06308_);
  nor (_06320_, _06318_, _06308_);
  nor (_06321_, _06320_, _06319_);
  and (_06322_, _06304_, _06288_);
  nor (_06323_, _06322_, _06305_);
  and (_06324_, _06323_, _06321_);
  nor (_06325_, _06324_, _06305_);
  nor (_06326_, _06298_, _06293_);
  and (_06327_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_06328_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_06329_, _06328_, _06327_);
  nor (_06330_, _06328_, _06327_);
  nor (_06331_, _06330_, _06329_);
  not (_06332_, _06331_);
  nor (_06333_, _06332_, _06326_);
  and (_06334_, _06332_, _06326_);
  nor (_06335_, _06334_, _06333_);
  and (_06336_, _06335_, _06312_);
  nor (_06337_, _06335_, _06312_);
  nor (_06338_, _06337_, _06336_);
  nor (_06339_, _06301_, _06270_);
  and (_06340_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_06341_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_06342_, _06341_, _06292_);
  nor (_06343_, _06341_, _06292_);
  nor (_06344_, _06343_, _06342_);
  and (_06345_, _06344_, _06340_);
  nor (_06346_, _06344_, _06340_);
  nor (_06347_, _06346_, _06345_);
  not (_06348_, _06347_);
  nor (_06349_, _06348_, _06339_);
  and (_06350_, _06348_, _06339_);
  nor (_06351_, _06350_, _06349_);
  and (_06352_, _06351_, _06338_);
  nor (_06353_, _06351_, _06338_);
  nor (_06354_, _06353_, _06352_);
  not (_06355_, _06354_);
  nor (_06356_, _06355_, _06325_);
  nor (_06357_, _06319_, _06316_);
  not (_06358_, _06357_);
  and (_06359_, _06355_, _06325_);
  nor (_06360_, _06359_, _06356_);
  and (_06361_, _06360_, _06358_);
  nor (_06362_, _06361_, _06356_);
  nor (_06363_, _06336_, _06333_);
  not (_06364_, _06363_);
  nor (_06365_, _06352_, _06349_);
  not (_06366_, _06365_);
  and (_06367_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_06368_, _06367_, _06292_);
  and (_06369_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_06370_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_06371_, _06370_, _06369_);
  nor (_06372_, _06371_, _06368_);
  nor (_06373_, _06345_, _06342_);
  and (_06374_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_06375_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_06376_, _06375_, _06374_);
  nor (_06377_, _06375_, _06374_);
  nor (_06378_, _06377_, _06376_);
  not (_06379_, _06378_);
  nor (_06380_, _06379_, _06373_);
  and (_06381_, _06379_, _06373_);
  nor (_06382_, _06381_, _06380_);
  and (_06383_, _06382_, _06329_);
  nor (_06384_, _06382_, _06329_);
  nor (_06385_, _06384_, _06383_);
  and (_06386_, _06385_, _06372_);
  nor (_06387_, _06385_, _06372_);
  nor (_06388_, _06387_, _06386_);
  and (_06389_, _06388_, _06366_);
  nor (_06390_, _06388_, _06366_);
  nor (_06391_, _06390_, _06389_);
  and (_06392_, _06391_, _06364_);
  nor (_06393_, _06391_, _06364_);
  nor (_06394_, _06393_, _06392_);
  not (_06395_, _06394_);
  nor (_06396_, _06395_, _06362_);
  nor (_06397_, _06392_, _06389_);
  nor (_06398_, _06383_, _06380_);
  not (_06399_, _06398_);
  and (_06400_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_06401_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_06402_, _06401_, _06400_);
  nor (_06403_, _06401_, _06400_);
  nor (_06404_, _06403_, _06402_);
  and (_06405_, _06404_, _06368_);
  nor (_06406_, _06404_, _06368_);
  nor (_06407_, _06406_, _06405_);
  and (_06408_, _06407_, _06376_);
  nor (_06409_, _06407_, _06376_);
  nor (_06410_, _06409_, _06408_);
  and (_06411_, _06410_, _06367_);
  nor (_06412_, _06410_, _06367_);
  nor (_06413_, _06412_, _06411_);
  and (_06414_, _06413_, _06386_);
  nor (_06415_, _06413_, _06386_);
  nor (_06416_, _06415_, _06414_);
  and (_06417_, _06416_, _06399_);
  nor (_06418_, _06416_, _06399_);
  nor (_06419_, _06418_, _06417_);
  not (_06420_, _06419_);
  nor (_06421_, _06420_, _06397_);
  and (_06422_, _06420_, _06397_);
  nor (_06423_, _06422_, _06421_);
  and (_06424_, _06423_, _06396_);
  nor (_06425_, _06417_, _06414_);
  nor (_06426_, _06408_, _06405_);
  not (_06427_, _06426_);
  and (_06428_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_06429_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_06430_, _06429_, _06428_);
  nor (_06431_, _06429_, _06428_);
  nor (_06432_, _06431_, _06430_);
  and (_06433_, _06432_, _06402_);
  nor (_06434_, _06432_, _06402_);
  nor (_06435_, _06434_, _06433_);
  and (_06436_, _06435_, _06411_);
  nor (_06437_, _06435_, _06411_);
  nor (_06438_, _06437_, _06436_);
  and (_06439_, _06438_, _06427_);
  nor (_06440_, _06438_, _06427_);
  nor (_06441_, _06440_, _06439_);
  not (_06442_, _06441_);
  nor (_06443_, _06442_, _06425_);
  and (_06444_, _06442_, _06425_);
  nor (_06445_, _06444_, _06443_);
  and (_06446_, _06445_, _06421_);
  nor (_06447_, _06445_, _06421_);
  nor (_06448_, _06447_, _06446_);
  and (_06449_, _06448_, _06424_);
  nor (_06450_, _06448_, _06424_);
  and (_06451_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_06452_, _06451_, _06264_);
  and (_06453_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_06454_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_06455_, _06454_, _06260_);
  nor (_06456_, _06455_, _06452_);
  and (_06457_, _06456_, _06453_);
  nor (_06458_, _06457_, _06452_);
  not (_06459_, _06458_);
  nor (_06460_, _06266_, _06262_);
  nor (_06461_, _06460_, _06267_);
  and (_06462_, _06461_, _06459_);
  and (_06463_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_06464_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_06465_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_06466_, _06465_, _06464_);
  nor (_06467_, _06465_, _06464_);
  nor (_06468_, _06467_, _06466_);
  and (_06469_, _06468_, _06463_);
  nor (_06470_, _06468_, _06463_);
  nor (_06471_, _06470_, _06469_);
  nor (_06472_, _06461_, _06459_);
  nor (_06473_, _06472_, _06462_);
  and (_06474_, _06473_, _06471_);
  nor (_06475_, _06474_, _06462_);
  nor (_06476_, _06286_, _06284_);
  nor (_06477_, _06476_, _06287_);
  not (_06478_, _06477_);
  nor (_06479_, _06478_, _06475_);
  and (_06480_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_06481_, _06480_, _06307_);
  nor (_06482_, _06469_, _06466_);
  nor (_06483_, _06307_, _06306_);
  nor (_06484_, _06483_, _06308_);
  not (_06485_, _06484_);
  nor (_06486_, _06485_, _06482_);
  and (_06487_, _06485_, _06482_);
  nor (_06488_, _06487_, _06486_);
  and (_06489_, _06488_, _06481_);
  nor (_06490_, _06488_, _06481_);
  nor (_06491_, _06490_, _06489_);
  and (_06492_, _06478_, _06475_);
  nor (_06493_, _06492_, _06479_);
  and (_06494_, _06493_, _06491_);
  nor (_06495_, _06494_, _06479_);
  nor (_06496_, _06323_, _06321_);
  nor (_06497_, _06496_, _06324_);
  not (_06498_, _06497_);
  nor (_06499_, _06498_, _06495_);
  nor (_06500_, _06489_, _06486_);
  not (_06501_, _06500_);
  and (_06502_, _06498_, _06495_);
  nor (_06503_, _06502_, _06499_);
  and (_06504_, _06503_, _06501_);
  nor (_06505_, _06504_, _06499_);
  nor (_06506_, _06360_, _06358_);
  nor (_06507_, _06506_, _06361_);
  not (_06508_, _06507_);
  nor (_06509_, _06508_, _06505_);
  and (_06510_, _06395_, _06362_);
  nor (_06511_, _06510_, _06396_);
  and (_06512_, _06511_, _06509_);
  nor (_06513_, _06423_, _06396_);
  nor (_06514_, _06513_, _06424_);
  and (_06515_, _06514_, _06512_);
  and (_06516_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_06517_, _06516_, _06451_);
  and (_06518_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_06519_, _06516_, _06451_);
  nor (_06520_, _06519_, _06517_);
  and (_06521_, _06520_, _06518_);
  nor (_06522_, _06521_, _06517_);
  not (_06523_, _06522_);
  nor (_06524_, _06456_, _06453_);
  nor (_06525_, _06524_, _06457_);
  and (_06526_, _06525_, _06523_);
  and (_06527_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_06528_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_06529_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_06530_, _06529_, _06528_);
  nor (_06531_, _06529_, _06528_);
  nor (_06532_, _06531_, _06530_);
  and (_06533_, _06532_, _06527_);
  nor (_06534_, _06532_, _06527_);
  nor (_06535_, _06534_, _06533_);
  nor (_06536_, _06525_, _06523_);
  nor (_06537_, _06536_, _06526_);
  and (_06538_, _06537_, _06535_);
  nor (_06539_, _06538_, _06526_);
  not (_06540_, _06539_);
  nor (_06541_, _06473_, _06471_);
  nor (_06542_, _06541_, _06474_);
  and (_06543_, _06542_, _06540_);
  nor (_06544_, _06533_, _06530_);
  and (_06545_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_06546_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_06547_, _06546_, _06545_);
  nor (_06548_, _06547_, _06481_);
  not (_06549_, _06548_);
  nor (_06550_, _06549_, _06544_);
  and (_06551_, _06549_, _06544_);
  nor (_06552_, _06551_, _06550_);
  nor (_06553_, _06542_, _06540_);
  nor (_06554_, _06553_, _06543_);
  and (_06555_, _06554_, _06552_);
  nor (_06556_, _06555_, _06543_);
  nor (_06557_, _06493_, _06491_);
  nor (_06558_, _06557_, _06494_);
  not (_06559_, _06558_);
  nor (_06560_, _06559_, _06556_);
  and (_06561_, _06559_, _06556_);
  nor (_06562_, _06561_, _06560_);
  and (_06563_, _06562_, _06550_);
  nor (_06564_, _06563_, _06560_);
  nor (_06565_, _06503_, _06501_);
  nor (_06566_, _06565_, _06504_);
  not (_06567_, _06566_);
  nor (_06568_, _06567_, _06564_);
  and (_06569_, _06508_, _06505_);
  nor (_06570_, _06569_, _06509_);
  and (_06571_, _06570_, _06568_);
  nor (_06572_, _06511_, _06509_);
  nor (_06573_, _06572_, _06512_);
  and (_06575_, _06573_, _06571_);
  nor (_06576_, _06573_, _06571_);
  nor (_06577_, _06576_, _06575_);
  and (_06578_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_06579_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_06580_, _06579_, _06578_);
  and (_06581_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06582_, _06579_, _06578_);
  nor (_06583_, _06582_, _06580_);
  and (_06584_, _06583_, _06581_);
  nor (_06585_, _06584_, _06580_);
  not (_06586_, _06585_);
  nor (_06587_, _06520_, _06518_);
  nor (_06588_, _06587_, _06521_);
  and (_06589_, _06588_, _06586_);
  and (_06590_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_06591_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_06592_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_06593_, _06592_, _06591_);
  nor (_06594_, _06592_, _06591_);
  nor (_06595_, _06594_, _06593_);
  and (_06596_, _06595_, _06590_);
  nor (_06597_, _06595_, _06590_);
  nor (_06598_, _06597_, _06596_);
  nor (_06599_, _06588_, _06586_);
  nor (_06600_, _06599_, _06589_);
  and (_06601_, _06600_, _06598_);
  nor (_06602_, _06601_, _06589_);
  not (_06603_, _06602_);
  nor (_06604_, _06537_, _06535_);
  nor (_06605_, _06604_, _06538_);
  and (_06606_, _06605_, _06603_);
  not (_06607_, _06480_);
  nor (_06608_, _06596_, _06593_);
  nor (_06609_, _06608_, _06607_);
  and (_06610_, _06608_, _06607_);
  nor (_06611_, _06610_, _06609_);
  nor (_06612_, _06605_, _06603_);
  nor (_06613_, _06612_, _06606_);
  and (_06614_, _06613_, _06611_);
  nor (_06615_, _06614_, _06606_);
  not (_06616_, _06615_);
  nor (_06617_, _06554_, _06552_);
  nor (_06618_, _06617_, _06555_);
  and (_06619_, _06618_, _06616_);
  nor (_06620_, _06618_, _06616_);
  nor (_06621_, _06620_, _06619_);
  and (_06622_, _06621_, _06609_);
  nor (_06623_, _06622_, _06619_);
  nor (_06624_, _06562_, _06550_);
  nor (_06625_, _06624_, _06563_);
  not (_06626_, _06625_);
  nor (_06627_, _06626_, _06623_);
  and (_06628_, _06567_, _06564_);
  nor (_06629_, _06628_, _06568_);
  and (_06630_, _06629_, _06627_);
  nor (_06631_, _06570_, _06568_);
  nor (_06632_, _06631_, _06571_);
  and (_06633_, _06632_, _06630_);
  nor (_06634_, _06632_, _06630_);
  nor (_06635_, _06634_, _06633_);
  and (_06636_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_06637_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_06638_, _06637_, _06636_);
  and (_06639_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_06640_, _06637_, _06636_);
  nor (_06641_, _06640_, _06638_);
  and (_06642_, _06641_, _06639_);
  nor (_06643_, _06642_, _06638_);
  not (_06644_, _06643_);
  nor (_06645_, _06583_, _06581_);
  nor (_06646_, _06645_, _06584_);
  and (_06647_, _06646_, _06644_);
  and (_06648_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_06649_, _06648_, _06592_);
  and (_06650_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_06651_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_06652_, _06651_, _06650_);
  nor (_06653_, _06652_, _06649_);
  nor (_06654_, _06646_, _06644_);
  nor (_06655_, _06654_, _06647_);
  and (_06656_, _06655_, _06653_);
  nor (_06657_, _06656_, _06647_);
  not (_06658_, _06657_);
  nor (_06659_, _06600_, _06598_);
  nor (_06660_, _06659_, _06601_);
  and (_06661_, _06660_, _06658_);
  nor (_06662_, _06660_, _06658_);
  nor (_06663_, _06662_, _06661_);
  and (_06664_, _06663_, _06649_);
  nor (_06665_, _06664_, _06661_);
  not (_06666_, _06665_);
  nor (_06667_, _06613_, _06611_);
  nor (_06668_, _06667_, _06614_);
  and (_06669_, _06668_, _06666_);
  nor (_06670_, _06621_, _06609_);
  nor (_06671_, _06670_, _06622_);
  and (_06672_, _06671_, _06669_);
  and (_06673_, _06626_, _06623_);
  nor (_06674_, _06673_, _06627_);
  and (_06675_, _06674_, _06672_);
  nor (_06676_, _06629_, _06627_);
  nor (_06677_, _06676_, _06630_);
  and (_06678_, _06677_, _06675_);
  nor (_06679_, _06677_, _06675_);
  nor (_06680_, _06679_, _06678_);
  and (_06681_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_06682_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_06683_, _06682_, _06681_);
  and (_06684_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_06685_, _06682_, _06681_);
  nor (_06686_, _06685_, _06683_);
  and (_06687_, _06686_, _06684_);
  nor (_06688_, _06687_, _06683_);
  not (_06689_, _06688_);
  nor (_06690_, _06641_, _06639_);
  nor (_06691_, _06690_, _06642_);
  and (_06692_, _06691_, _06689_);
  nor (_06693_, _06691_, _06689_);
  nor (_06694_, _06693_, _06692_);
  and (_06695_, _06694_, _06648_);
  nor (_06696_, _06695_, _06692_);
  not (_06697_, _06696_);
  nor (_06698_, _06655_, _06653_);
  nor (_06699_, _06698_, _06656_);
  and (_06700_, _06699_, _06697_);
  nor (_06701_, _06663_, _06649_);
  nor (_06702_, _06701_, _06664_);
  and (_06703_, _06702_, _06700_);
  nor (_06704_, _06668_, _06666_);
  nor (_06705_, _06704_, _06669_);
  and (_06706_, _06705_, _06703_);
  nor (_06707_, _06671_, _06669_);
  nor (_06708_, _06707_, _06672_);
  and (_06709_, _06708_, _06706_);
  nor (_06710_, _06674_, _06672_);
  nor (_06711_, _06710_, _06675_);
  and (_06712_, _06711_, _06709_);
  and (_06713_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_06714_, _06713_, _06682_);
  nor (_06715_, _06686_, _06684_);
  nor (_06716_, _06715_, _06687_);
  and (_06717_, _06716_, _06714_);
  nor (_06718_, _06694_, _06648_);
  nor (_06719_, _06718_, _06695_);
  and (_06720_, _06719_, _06717_);
  nor (_06721_, _06699_, _06697_);
  nor (_06722_, _06721_, _06700_);
  and (_06723_, _06722_, _06720_);
  nor (_06724_, _06702_, _06700_);
  nor (_06725_, _06724_, _06703_);
  and (_06726_, _06725_, _06723_);
  nor (_06727_, _06705_, _06703_);
  nor (_06728_, _06727_, _06706_);
  and (_06729_, _06728_, _06726_);
  nor (_06730_, _06708_, _06706_);
  nor (_06731_, _06730_, _06709_);
  and (_06732_, _06731_, _06729_);
  nor (_06733_, _06711_, _06709_);
  nor (_06734_, _06733_, _06712_);
  and (_06735_, _06734_, _06732_);
  nor (_06736_, _06735_, _06712_);
  not (_06737_, _06736_);
  and (_06738_, _06737_, _06680_);
  nor (_06739_, _06738_, _06678_);
  not (_06740_, _06739_);
  and (_06741_, _06740_, _06635_);
  nor (_06742_, _06741_, _06633_);
  not (_06743_, _06742_);
  and (_06744_, _06743_, _06577_);
  nor (_06745_, _06744_, _06575_);
  not (_06746_, _06745_);
  nor (_06747_, _06514_, _06512_);
  nor (_06748_, _06747_, _06515_);
  and (_06749_, _06748_, _06746_);
  nor (_06750_, _06749_, _06515_);
  nor (_06751_, _06750_, _06450_);
  or (_06752_, _06751_, _06449_);
  and (_06753_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_06754_, _06753_);
  nor (_06755_, _06754_, _06401_);
  nor (_06756_, _06755_, _06433_);
  nor (_06757_, _06439_, _06436_);
  nor (_06758_, _06757_, _06756_);
  and (_06759_, _06757_, _06756_);
  nor (_06760_, _06759_, _06758_);
  not (_06761_, _06760_);
  nor (_06762_, _06446_, _06443_);
  and (_06763_, _06762_, _06761_);
  nor (_06764_, _06762_, _06761_);
  nor (_06765_, _06764_, _06763_);
  and (_06766_, _06765_, _06752_);
  or (_06767_, _06758_, _06430_);
  or (_06768_, _06767_, _06764_);
  or (_06769_, _06768_, _06766_);
  or (_06770_, _06769_, _06258_);
  and (_06771_, _06770_, _02986_);
  and (_06772_, _06771_, _06257_);
  not (_06773_, _05321_);
  nor (_06774_, _05531_, _06773_);
  or (_06775_, _06774_, _06236_);
  and (_06776_, _06775_, _02866_);
  or (_06777_, _06776_, _05535_);
  or (_06778_, _06777_, _06772_);
  and (_06779_, _06778_, _06223_);
  or (_06780_, _06779_, _02841_);
  and (_06781_, _05461_, _04721_);
  or (_06782_, _06214_, _02842_);
  or (_06783_, _06782_, _06781_);
  and (_06784_, _06783_, _02839_);
  and (_06785_, _06784_, _06780_);
  and (_06786_, _03028_, _02515_);
  nor (_06787_, _05740_, _06220_);
  or (_06788_, _06787_, _06214_);
  and (_06789_, _06788_, _02567_);
  or (_06790_, _06789_, _06786_);
  or (_06791_, _06790_, _06785_);
  not (_06792_, _06786_);
  not (_06793_, \oc8051_golden_model_1.B [1]);
  nor (_06794_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_06795_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_06796_, _06795_, _06794_);
  and (_06797_, _06796_, _06793_);
  not (_06798_, \oc8051_golden_model_1.B [0]);
  and (_06799_, _06798_, \oc8051_golden_model_1.ACC [7]);
  nor (_06800_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_06801_, _06800_, _06799_);
  and (_06802_, _06801_, _06797_);
  or (_06803_, _06798_, \oc8051_golden_model_1.ACC [7]);
  and (_06804_, _06800_, _06797_);
  and (_06805_, _06804_, _06803_);
  or (_06806_, _06805_, _05364_);
  not (_06807_, \oc8051_golden_model_1.ACC [6]);
  and (_06808_, \oc8051_golden_model_1.B [0], _06807_);
  nor (_06809_, _06808_, _05364_);
  nor (_06810_, _06809_, _06793_);
  and (_06811_, _06800_, _06796_);
  not (_06812_, _06811_);
  nor (_06813_, _06812_, _06810_);
  nor (_06814_, _06813_, _06806_);
  nor (_06815_, _06814_, _06802_);
  and (_06816_, _06813_, \oc8051_golden_model_1.B [0]);
  nor (_06817_, _06816_, _06807_);
  and (_06818_, _06817_, _06793_);
  nor (_06819_, _06817_, _06793_);
  nor (_06820_, _06819_, _06818_);
  nor (_06821_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_06822_, _06821_, _06451_);
  nor (_06823_, _06822_, \oc8051_golden_model_1.ACC [4]);
  nor (_06824_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_06825_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_06826_, _06825_, _06798_);
  nor (_06827_, _06826_, _06824_);
  nor (_06828_, _06827_, _06823_);
  not (_06829_, _06828_);
  and (_06830_, _06829_, _06820_);
  not (_06831_, _06830_);
  nor (_06832_, _06815_, \oc8051_golden_model_1.B [2]);
  nor (_06833_, _06832_, _06818_);
  and (_06834_, _06833_, _06831_);
  not (_06835_, _06834_);
  and (_06836_, _06796_, _06211_);
  and (_06837_, \oc8051_golden_model_1.B [2], _05364_);
  not (_06838_, _06837_);
  and (_06839_, _06838_, _06836_);
  and (_06840_, _06839_, _06835_);
  nor (_06841_, _06840_, _06815_);
  nor (_06842_, _06841_, _06802_);
  nor (_06843_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_06844_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_06845_, _06844_, \oc8051_golden_model_1.ACC [7]);
  and (_06846_, _06845_, _06843_);
  nor (_06847_, _06846_, _06836_);
  nor (_06848_, _06842_, \oc8051_golden_model_1.B [3]);
  nor (_06849_, _06829_, _06820_);
  nor (_06850_, _06849_, _06830_);
  and (_06851_, _06850_, _06840_);
  not (_06852_, _06817_);
  nor (_06853_, _06840_, _06852_);
  nor (_06854_, _06853_, _06851_);
  nor (_06855_, _06854_, \oc8051_golden_model_1.B [2]);
  and (_06856_, _06854_, \oc8051_golden_model_1.B [2]);
  nor (_06857_, _06856_, _06855_);
  not (_06858_, \oc8051_golden_model_1.ACC [5]);
  nor (_06859_, _06840_, _06858_);
  and (_06860_, _06840_, _06822_);
  or (_06861_, _06860_, _06859_);
  and (_06862_, _06861_, _06793_);
  nor (_06863_, _06861_, _06793_);
  not (_06864_, \oc8051_golden_model_1.ACC [4]);
  and (_06865_, \oc8051_golden_model_1.B [0], _06864_);
  nor (_06866_, _06865_, _06863_);
  nor (_06867_, _06866_, _06862_);
  not (_06868_, _06867_);
  and (_06869_, _06868_, _06857_);
  or (_06870_, _06869_, _06855_);
  nor (_06871_, _06870_, _06848_);
  nor (_06872_, _06871_, _06847_);
  nor (_06873_, _06872_, _06842_);
  nor (_06874_, _06873_, _06802_);
  nor (_06875_, _06874_, \oc8051_golden_model_1.B [4]);
  not (_06876_, \oc8051_golden_model_1.B [3]);
  nor (_06877_, _06872_, _06854_);
  nor (_06878_, _06868_, _06857_);
  nor (_06879_, _06878_, _06869_);
  and (_06880_, _06879_, _06872_);
  or (_06881_, _06880_, _06877_);
  and (_06882_, _06881_, _06876_);
  nor (_06883_, _06881_, _06876_);
  nor (_06884_, _06883_, _06882_);
  not (_06885_, _06884_);
  nor (_06886_, _06872_, _06861_);
  nor (_06887_, _06863_, _06862_);
  and (_06888_, _06887_, _06865_);
  nor (_06889_, _06887_, _06865_);
  nor (_06890_, _06889_, _06888_);
  and (_06891_, _06890_, _06872_);
  or (_06892_, _06891_, _06886_);
  nor (_06893_, _06892_, \oc8051_golden_model_1.B [2]);
  and (_06894_, _06892_, \oc8051_golden_model_1.B [2]);
  nor (_06895_, _06872_, _06864_);
  nor (_06896_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_06897_, _06896_, _06578_);
  and (_06898_, _06872_, _06897_);
  or (_06899_, _06898_, _06895_);
  and (_06900_, _06899_, _06793_);
  nor (_06901_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_06902_, _06901_, _06636_);
  nor (_06903_, _06902_, \oc8051_golden_model_1.ACC [2]);
  nor (_06904_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_06905_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_06906_, _06905_, _06798_);
  nor (_06907_, _06906_, _06904_);
  nor (_06908_, _06907_, _06903_);
  not (_06909_, _06908_);
  nor (_06910_, _06899_, _06793_);
  nor (_06911_, _06910_, _06900_);
  and (_06912_, _06911_, _06909_);
  nor (_06913_, _06912_, _06900_);
  nor (_06914_, _06913_, _06894_);
  nor (_06915_, _06914_, _06893_);
  nor (_06916_, _06915_, _06885_);
  or (_06917_, _06916_, _06882_);
  nor (_06918_, _06917_, _06875_);
  not (_06919_, \oc8051_golden_model_1.B [5]);
  and (_06920_, _06844_, _06919_);
  not (_06921_, _06920_);
  and (_06922_, \oc8051_golden_model_1.B [4], _05364_);
  nor (_06923_, _06922_, _06921_);
  not (_06924_, _06923_);
  nor (_06925_, _06924_, _06918_);
  nor (_06926_, _06925_, _06874_);
  nor (_06927_, _06926_, _06802_);
  nor (_06928_, _06845_, _06920_);
  nor (_06929_, _06927_, \oc8051_golden_model_1.B [5]);
  not (_06930_, \oc8051_golden_model_1.B [4]);
  and (_06931_, _06915_, _06885_);
  nor (_06932_, _06931_, _06916_);
  not (_06933_, _06932_);
  and (_06934_, _06933_, _06925_);
  nor (_06935_, _06925_, _06881_);
  nor (_06936_, _06935_, _06934_);
  and (_06937_, _06936_, _06930_);
  nor (_06938_, _06936_, _06930_);
  nor (_06939_, _06938_, _06937_);
  not (_06940_, _06939_);
  nor (_06941_, _06925_, _06892_);
  nor (_06942_, _06894_, _06893_);
  and (_06943_, _06942_, _06913_);
  nor (_06944_, _06942_, _06913_);
  nor (_06945_, _06944_, _06943_);
  not (_06946_, _06945_);
  and (_06947_, _06946_, _06925_);
  nor (_06948_, _06947_, _06941_);
  nor (_06949_, _06948_, \oc8051_golden_model_1.B [3]);
  and (_06950_, _06948_, \oc8051_golden_model_1.B [3]);
  not (_06951_, \oc8051_golden_model_1.B [2]);
  nor (_06952_, _06911_, _06909_);
  nor (_06953_, _06952_, _06912_);
  not (_06954_, _06953_);
  and (_06955_, _06954_, _06925_);
  nor (_06956_, _06925_, _06899_);
  nor (_06957_, _06956_, _06955_);
  and (_06958_, _06957_, _06951_);
  nor (_06959_, _06925_, _02625_);
  and (_06960_, _06925_, _06902_);
  or (_06961_, _06960_, _06959_);
  and (_06962_, _06961_, _06793_);
  nor (_06963_, _06961_, _06793_);
  not (_06964_, \oc8051_golden_model_1.ACC [2]);
  and (_06965_, \oc8051_golden_model_1.B [0], _06964_);
  nor (_06966_, _06965_, _06963_);
  nor (_06967_, _06966_, _06962_);
  nor (_06968_, _06957_, _06951_);
  nor (_06969_, _06968_, _06958_);
  not (_06970_, _06969_);
  nor (_06971_, _06970_, _06967_);
  nor (_06972_, _06971_, _06958_);
  nor (_06973_, _06972_, _06950_);
  nor (_06974_, _06973_, _06949_);
  nor (_06975_, _06974_, _06940_);
  or (_06976_, _06975_, _06937_);
  nor (_06977_, _06976_, _06929_);
  nor (_06978_, _06977_, _06928_);
  nor (_06979_, _06978_, _06927_);
  nor (_06980_, _06979_, _06802_);
  nor (_06981_, _06980_, \oc8051_golden_model_1.B [6]);
  and (_06982_, \oc8051_golden_model_1.B [6], _05364_);
  not (_06983_, _06978_);
  and (_06984_, _06974_, _06940_);
  nor (_06985_, _06984_, _06975_);
  nor (_06986_, _06985_, _06983_);
  nor (_06987_, _06978_, _06936_);
  nor (_06988_, _06987_, _06986_);
  and (_06989_, _06988_, _06919_);
  nor (_06990_, _06988_, _06919_);
  nor (_06991_, _06990_, _06989_);
  nor (_06992_, _06978_, _06948_);
  nor (_06993_, _06950_, _06949_);
  nor (_06994_, _06993_, _06972_);
  and (_06995_, _06993_, _06972_);
  or (_06996_, _06995_, _06994_);
  and (_06997_, _06996_, _06978_);
  or (_06998_, _06997_, _06992_);
  and (_06999_, _06998_, _06930_);
  nor (_07000_, _06998_, _06930_);
  and (_07001_, _06970_, _06967_);
  nor (_07002_, _07001_, _06971_);
  nor (_07003_, _07002_, _06983_);
  nor (_07004_, _06978_, _06957_);
  nor (_07005_, _07004_, _07003_);
  and (_07006_, _07005_, _06876_);
  nor (_07007_, _06963_, _06962_);
  nor (_07008_, _07007_, _06965_);
  and (_07009_, _07007_, _06965_);
  or (_07010_, _07009_, _07008_);
  nor (_07011_, _07010_, _06983_);
  nor (_07012_, _06978_, _06961_);
  nor (_07013_, _07012_, _07011_);
  and (_07014_, _07013_, _06951_);
  nor (_07015_, _07013_, _06951_);
  nor (_07016_, _06978_, _06964_);
  nor (_07017_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07018_, _07017_, _06681_);
  and (_07019_, _06978_, _07018_);
  or (_07020_, _07019_, _07016_);
  and (_07021_, _07020_, _06793_);
  and (_07022_, \oc8051_golden_model_1.B [0], _02543_);
  not (_07023_, _07022_);
  nor (_07024_, _07020_, _06793_);
  nor (_07025_, _07024_, _07021_);
  and (_07026_, _07025_, _07023_);
  nor (_07027_, _07026_, _07021_);
  nor (_07028_, _07027_, _07015_);
  nor (_07029_, _07028_, _07014_);
  not (_07030_, _07029_);
  nor (_07031_, _07005_, _06876_);
  nor (_07032_, _07031_, _07006_);
  and (_07033_, _07032_, _07030_);
  nor (_07034_, _07033_, _07006_);
  nor (_07035_, _07034_, _07000_);
  nor (_07036_, _07035_, _06999_);
  not (_07037_, _07036_);
  and (_07038_, _07037_, _06991_);
  nor (_07039_, _07038_, _06989_);
  nor (_07040_, _07039_, _06982_);
  nor (_07041_, _07040_, _06981_);
  nor (_07042_, _07041_, \oc8051_golden_model_1.B [7]);
  nor (_07043_, _07042_, _06980_);
  or (_07044_, _07043_, _06802_);
  nor (_07045_, _07044_, \oc8051_golden_model_1.B [7]);
  nor (_07046_, _07045_, _06753_);
  nor (_07047_, _07037_, _06991_);
  nor (_07048_, _07047_, _07038_);
  and (_07049_, _07048_, _07042_);
  not (_07050_, _07042_);
  and (_07051_, _07050_, _06988_);
  nor (_07052_, _07051_, _07049_);
  and (_07053_, _07052_, \oc8051_golden_model_1.B [6]);
  not (_07054_, _07053_);
  nor (_07055_, _07054_, _07046_);
  nor (_07056_, _07015_, _07014_);
  nor (_07057_, _07056_, _07027_);
  and (_07058_, _07056_, _07027_);
  or (_07059_, _07058_, _07057_);
  nor (_07060_, _07059_, _07050_);
  nor (_07061_, _07042_, _07013_);
  nor (_07062_, _07061_, _07060_);
  nor (_07063_, _07062_, _06876_);
  and (_07064_, _07062_, _06876_);
  nor (_07065_, _07064_, _07063_);
  nor (_07066_, _07025_, _07023_);
  or (_07067_, _07066_, _07026_);
  and (_07068_, _07067_, _07042_);
  nor (_07069_, _07042_, _07020_);
  nor (_07070_, _07069_, _07068_);
  nor (_07071_, _07070_, _06951_);
  and (_07072_, _07070_, _06951_);
  nor (_07073_, _07072_, _07071_);
  and (_07074_, _07073_, _07065_);
  nor (_07075_, _07042_, \oc8051_golden_model_1.ACC [1]);
  and (_07076_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07077_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  or (_07078_, _07077_, _07076_);
  and (_07079_, _07042_, _07078_);
  nor (_07080_, _07079_, _07075_);
  and (_07081_, _07080_, _06793_);
  nor (_07082_, _07080_, _06793_);
  and (_07083_, _06798_, \oc8051_golden_model_1.ACC [0]);
  not (_07084_, _07083_);
  nor (_07085_, _07084_, _07082_);
  nor (_07086_, _07085_, _07081_);
  and (_07087_, _07086_, _07074_);
  not (_07088_, _07087_);
  and (_07089_, _07071_, _07065_);
  nor (_07090_, _07089_, _07063_);
  and (_07091_, _07090_, _07088_);
  nor (_07092_, _07052_, \oc8051_golden_model_1.B [6]);
  nor (_07093_, _07092_, _07053_);
  not (_07094_, _07093_);
  nor (_07095_, _07094_, _07046_);
  nor (_07096_, _07032_, _07030_);
  nor (_07097_, _07096_, _07033_);
  and (_07098_, _07097_, _07042_);
  and (_07099_, _07050_, _07005_);
  nor (_07100_, _07099_, _07098_);
  and (_07101_, _07100_, \oc8051_golden_model_1.B [4]);
  nor (_07102_, _07100_, \oc8051_golden_model_1.B [4]);
  nor (_07103_, _07102_, _07101_);
  nor (_07104_, _07000_, _06999_);
  nor (_07105_, _07104_, _07034_);
  and (_07106_, _07104_, _07034_);
  or (_07107_, _07106_, _07105_);
  nor (_07108_, _07107_, _07050_);
  nor (_07109_, _07042_, _06998_);
  nor (_07110_, _07109_, _07108_);
  nor (_07111_, _07110_, _06919_);
  and (_07112_, _07110_, _06919_);
  nor (_07113_, _07112_, _07111_);
  and (_07114_, _07113_, _07103_);
  and (_07115_, _07114_, _07095_);
  not (_07116_, _07115_);
  nor (_07117_, _07116_, _07091_);
  and (_07118_, _06980_, \oc8051_golden_model_1.B [7]);
  and (_07119_, _07113_, _07101_);
  nor (_07120_, _07119_, _07111_);
  not (_07121_, _07120_);
  and (_07122_, _07121_, _07095_);
  or (_07123_, _07122_, _07118_);
  or (_07124_, _07123_, _07117_);
  nor (_07125_, _07124_, _07055_);
  and (_07126_, \oc8051_golden_model_1.B [0], _02696_);
  not (_07127_, _07126_);
  nor (_07128_, _07082_, _07081_);
  and (_07129_, _07128_, _07127_);
  and (_07130_, _07129_, _07084_);
  and (_07131_, _07130_, _07074_);
  and (_07132_, _07131_, _07115_);
  nor (_07133_, _07132_, _07125_);
  or (_07134_, _07133_, _06802_);
  and (_07135_, _07134_, _07044_);
  or (_07136_, _07135_, _06792_);
  and (_07137_, _07136_, _06791_);
  or (_07138_, _07137_, _02834_);
  not (_07139_, _03051_);
  not (_07140_, _02834_);
  or (_07141_, _06217_, _07140_);
  and (_07142_, _07141_, _07139_);
  and (_07143_, _07142_, _07138_);
  and (_07144_, _05764_, _04721_);
  or (_07145_, _06214_, _03148_);
  nor (_07146_, _07145_, _07144_);
  nor (_07147_, _07146_, _03149_);
  or (_07148_, _07147_, _07143_);
  and (_07149_, _05772_, _04721_);
  not (_07150_, _03148_);
  or (_07151_, _06214_, _07150_);
  or (_07152_, _07151_, _07149_);
  and (_07153_, _07152_, _03023_);
  and (_07154_, _07153_, _07148_);
  or (_07155_, _07154_, _06219_);
  and (_07156_, _07155_, _06213_);
  and (_07157_, _06228_, _03137_);
  and (_07158_, _07157_, _06215_);
  or (_07159_, _07158_, _03042_);
  or (_07160_, _07159_, _07156_);
  not (_07161_, _03143_);
  nor (_07162_, _05763_, _06220_);
  or (_07163_, _06214_, _03043_);
  or (_07164_, _07163_, _07162_);
  and (_07165_, _07164_, _07161_);
  and (_07166_, _07165_, _07160_);
  nor (_07167_, _05771_, _06220_);
  or (_07168_, _07167_, _06214_);
  and (_07169_, _07168_, _03143_);
  or (_07170_, _07169_, _03174_);
  or (_07171_, _07170_, _07166_);
  or (_07172_, _06225_, _03179_);
  and (_07173_, _07172_, _03183_);
  and (_07174_, _07173_, _07171_);
  and (_07175_, _06248_, _02799_);
  or (_07176_, _07175_, _02887_);
  or (_07177_, _07176_, _07174_);
  and (_07178_, _05246_, _04721_);
  or (_07179_, _06214_, _02888_);
  or (_07180_, _07179_, _07178_);
  and (_07181_, _07180_, _34655_);
  and (_07182_, _07181_, _07177_);
  or (_07183_, _07182_, _06212_);
  and (_35828_[7], _07183_, _35796_);
  nor (_07184_, _34655_, _05364_);
  and (_07185_, _02840_, _02509_);
  nor (_07186_, _03728_, _03272_);
  and (_07187_, _02845_, _02509_);
  nor (_07188_, _07187_, _03570_);
  and (_07189_, _07188_, _07186_);
  and (_07190_, _04630_, _05364_);
  nor (_07191_, _04630_, _05364_);
  nor (_07192_, _07191_, _07190_);
  nor (_07193_, _04790_, _06807_);
  and (_07194_, _04790_, _06807_);
  nor (_07195_, _07194_, _07193_);
  nor (_07196_, _04894_, _06858_);
  and (_07197_, _04894_, _06858_);
  nor (_07198_, _07197_, _07196_);
  not (_07199_, _07198_);
  nor (_07200_, _05192_, _06864_);
  and (_07201_, _05192_, _06864_);
  nor (_07202_, _07201_, _07200_);
  nor (_07203_, _04275_, _02625_);
  and (_07204_, _04275_, _02625_);
  nor (_07205_, _04449_, _06964_);
  and (_07206_, _04449_, _06964_);
  nor (_07207_, _07206_, _07205_);
  not (_07208_, _07207_);
  nor (_07209_, _04020_, _02543_);
  and (_07210_, _04020_, _02543_);
  nor (_07211_, _07210_, _07209_);
  and (_07212_, _03838_, \oc8051_golden_model_1.ACC [0]);
  and (_07213_, _07212_, _07211_);
  nor (_07214_, _07213_, _07209_);
  nor (_07215_, _07214_, _07208_);
  nor (_07216_, _07215_, _07205_);
  nor (_07217_, _07216_, _07204_);
  or (_07218_, _07217_, _07203_);
  and (_07219_, _07218_, _07202_);
  nor (_07220_, _07219_, _07200_);
  nor (_07221_, _07220_, _07199_);
  or (_07222_, _07221_, _07196_);
  and (_07223_, _07222_, _07195_);
  nor (_07224_, _07223_, _07193_);
  nor (_07225_, _07224_, _07192_);
  and (_07226_, _07224_, _07192_);
  or (_07227_, _07226_, _07225_);
  or (_07228_, _07227_, _07189_);
  and (_07229_, _02840_, _02527_);
  nor (_07230_, _02856_, _03551_);
  and (_07231_, _02849_, _02539_);
  nand (_07232_, _07231_, _02527_);
  not (_07233_, _07232_);
  nor (_07234_, _07233_, _07230_);
  not (_07235_, _04790_);
  and (_07236_, _05254_, _07235_);
  and (_07237_, _07236_, \oc8051_golden_model_1.PSW [7]);
  nor (_07238_, _07237_, _04630_);
  and (_07239_, _07237_, _04630_);
  nor (_07240_, _07239_, _07238_);
  and (_07241_, _07240_, \oc8051_golden_model_1.ACC [7]);
  nor (_07242_, _07240_, \oc8051_golden_model_1.ACC [7]);
  nor (_07243_, _07242_, _07241_);
  and (_07244_, _05254_, \oc8051_golden_model_1.PSW [7]);
  nor (_07245_, _07244_, _07235_);
  nor (_07246_, _07245_, _07237_);
  and (_07247_, _07246_, \oc8051_golden_model_1.ACC [6]);
  and (_07248_, _07246_, _06807_);
  nor (_07249_, _07246_, _06807_);
  nor (_07250_, _07249_, _07248_);
  and (_07251_, _05253_, \oc8051_golden_model_1.PSW [7]);
  nor (_07252_, _07251_, _05248_);
  nor (_07253_, _07252_, _07244_);
  and (_07254_, _07253_, \oc8051_golden_model_1.ACC [5]);
  and (_07255_, _07253_, _06858_);
  nor (_07256_, _07253_, _06858_);
  nor (_07257_, _07256_, _07255_);
  and (_07258_, _05250_, \oc8051_golden_model_1.PSW [7]);
  and (_07259_, _07258_, _05251_);
  nor (_07260_, _07259_, _05249_);
  nor (_07261_, _07260_, _07251_);
  and (_07262_, _07261_, \oc8051_golden_model_1.ACC [4]);
  nor (_07263_, _07261_, _06864_);
  and (_07264_, _07261_, _06864_);
  nor (_07265_, _07264_, _07263_);
  not (_07266_, _04275_);
  and (_07267_, _05250_, _04450_);
  and (_07268_, _07267_, \oc8051_golden_model_1.PSW [7]);
  nor (_07269_, _07268_, _07266_);
  nor (_07270_, _07269_, _07259_);
  and (_07271_, _07270_, \oc8051_golden_model_1.ACC [3]);
  nor (_07272_, _07270_, _02625_);
  and (_07273_, _07270_, _02625_);
  nor (_07274_, _07273_, _07272_);
  nor (_07275_, _07258_, _04450_);
  nor (_07276_, _07275_, _07268_);
  and (_07277_, _07276_, \oc8051_golden_model_1.ACC [2]);
  nor (_07278_, _07276_, _06964_);
  and (_07279_, _07276_, _06964_);
  nor (_07280_, _07279_, _07278_);
  and (_07281_, _03838_, \oc8051_golden_model_1.PSW [7]);
  nor (_07282_, _07281_, _04021_);
  nor (_07283_, _07282_, _07258_);
  and (_07284_, _07283_, \oc8051_golden_model_1.ACC [1]);
  nor (_07285_, _07283_, _02543_);
  and (_07286_, _07283_, _02543_);
  nor (_07287_, _07286_, _07285_);
  not (_07288_, \oc8051_golden_model_1.PSW [7]);
  and (_07289_, _03872_, _07288_);
  nor (_07290_, _07289_, _07281_);
  and (_07291_, _07290_, \oc8051_golden_model_1.ACC [0]);
  not (_07292_, _07291_);
  nor (_07293_, _07292_, _07287_);
  nor (_07294_, _07293_, _07284_);
  nor (_07295_, _07294_, _07280_);
  nor (_07296_, _07295_, _07277_);
  nor (_07297_, _07296_, _07274_);
  nor (_07298_, _07297_, _07271_);
  nor (_07299_, _07298_, _07265_);
  nor (_07300_, _07299_, _07262_);
  nor (_07301_, _07300_, _07257_);
  nor (_07302_, _07301_, _07254_);
  nor (_07303_, _07302_, _07250_);
  nor (_07304_, _07303_, _07247_);
  nor (_07305_, _07304_, _07243_);
  and (_07306_, _07304_, _07243_);
  nor (_07307_, _07306_, _07305_);
  or (_07308_, _07307_, _07234_);
  nor (_07309_, _02856_, _03543_);
  nand (_07310_, _07309_, _07190_);
  and (_07311_, _03028_, _02529_);
  not (_07312_, _07311_);
  or (_07313_, _05770_, _03136_);
  and (_07314_, _07313_, _07312_);
  nor (_07315_, _04731_, _05364_);
  and (_07316_, _05764_, _04731_);
  nor (_07317_, _07316_, _07315_);
  nand (_07318_, _07317_, _03051_);
  not (_07319_, _04731_);
  nor (_07320_, _07319_, _04630_);
  nor (_07321_, _07320_, _07315_);
  nand (_07322_, _07321_, _05535_);
  and (_07323_, _06174_, \oc8051_golden_model_1.PSW [7]);
  nor (_07324_, _07323_, _05461_);
  and (_07325_, _06173_, \oc8051_golden_model_1.PSW [7]);
  and (_07326_, _07325_, _06162_);
  and (_07327_, _07326_, _05461_);
  nor (_07328_, _07327_, _07324_);
  nor (_07329_, _07328_, _05364_);
  and (_07330_, _07328_, _05364_);
  nor (_07331_, _07330_, _07329_);
  not (_07332_, _07331_);
  nor (_07333_, _07325_, _06162_);
  nor (_07334_, _07333_, _07323_);
  nor (_07335_, _07334_, _06807_);
  and (_07336_, _07334_, _06807_);
  and (_07337_, _06169_, _06171_);
  and (_07338_, _07337_, \oc8051_golden_model_1.PSW [7]);
  nor (_07339_, _07338_, _06170_);
  nor (_07340_, _07339_, _07325_);
  and (_07341_, _07340_, _06858_);
  nor (_07342_, _07340_, _06858_);
  and (_07343_, _06165_, \oc8051_golden_model_1.PSW [7]);
  and (_07344_, _07343_, _06168_);
  nor (_07345_, _07344_, _06171_);
  nor (_07346_, _07345_, _07338_);
  nor (_07347_, _07346_, _06864_);
  nor (_07348_, _07347_, _07342_);
  nor (_07349_, _07348_, _07341_);
  nor (_07350_, _07342_, _07341_);
  and (_07351_, _07346_, _06864_);
  nor (_07352_, _07351_, _07347_);
  and (_07353_, _07352_, _07350_);
  not (_07354_, _07353_);
  and (_07355_, _06165_, _06167_);
  and (_07356_, _07355_, \oc8051_golden_model_1.PSW [7]);
  nor (_07357_, _07356_, _06166_);
  nor (_07358_, _07357_, _07344_);
  nor (_07359_, _07358_, _02625_);
  and (_07360_, _07358_, _02625_);
  nor (_07361_, _07360_, _07359_);
  nor (_07362_, _07343_, _06167_);
  nor (_07363_, _07362_, _07356_);
  nor (_07364_, _07363_, _06964_);
  and (_07365_, _07363_, _06964_);
  nor (_07366_, _07365_, _07364_);
  and (_07367_, _07366_, _07361_);
  and (_07368_, _06164_, \oc8051_golden_model_1.PSW [7]);
  nor (_07369_, _07368_, _06163_);
  nor (_07370_, _07369_, _07343_);
  and (_07371_, _07370_, _02543_);
  nor (_07372_, _07370_, _02543_);
  and (_07373_, _05945_, _07288_);
  nor (_07374_, _07373_, _07368_);
  nor (_07375_, _07374_, _02696_);
  nor (_07376_, _07375_, _07372_);
  nor (_07377_, _07376_, _07371_);
  not (_07378_, _07377_);
  and (_07379_, _07378_, _07367_);
  not (_07380_, _07379_);
  and (_07381_, _07365_, _07361_);
  nor (_07382_, _07381_, _07360_);
  and (_07383_, _07382_, _07380_);
  nor (_07384_, _07372_, _07371_);
  and (_07385_, _07374_, _02696_);
  nor (_07386_, _07375_, _07385_);
  and (_07387_, _07386_, _07384_);
  and (_07388_, _07387_, _07367_);
  nor (_07389_, _07388_, _07383_);
  nor (_07390_, _07389_, _07354_);
  nor (_07391_, _07390_, _07349_);
  nor (_07392_, _07391_, _07336_);
  or (_07393_, _07392_, _07335_);
  and (_07394_, _07393_, _07332_);
  nor (_07395_, _07393_, _07332_);
  or (_07396_, _07395_, _07394_);
  and (_07397_, _02840_, _02864_);
  and (_07398_, _07397_, _07396_);
  or (_07399_, _02568_, _02564_);
  not (_07400_, _07399_);
  nor (_07401_, _03765_, _03413_);
  and (_07402_, _07401_, _04046_);
  not (_07403_, _07402_);
  nand (_07404_, _07403_, _04630_);
  and (_07405_, _03028_, _02883_);
  and (_07406_, _05474_, _04731_);
  nor (_07407_, _07406_, _07315_);
  nand (_07408_, _07407_, _02948_);
  nor (_07409_, _05497_, _03401_);
  and (_07410_, _02840_, _02949_);
  not (_07411_, _07410_);
  or (_07412_, _07411_, _05461_);
  not (_07413_, _03724_);
  and (_07414_, _02962_, _02949_);
  not (_07415_, _07414_);
  nor (_07416_, _02966_, _02854_);
  nor (_07417_, _07416_, _02600_);
  nor (_07418_, _03019_, _02600_);
  nor (_07419_, _07418_, _07417_);
  and (_07420_, _07419_, _07415_);
  and (_07421_, _07420_, _07413_);
  nor (_07422_, _07421_, _04630_);
  and (_07423_, _03028_, _03382_);
  or (_07424_, _07423_, \oc8051_golden_model_1.ACC [7]);
  nand (_07425_, _07423_, \oc8051_golden_model_1.ACC [7]);
  and (_07426_, _07425_, _07424_);
  and (_07427_, _07426_, _07421_);
  or (_07428_, _07427_, _07410_);
  or (_07429_, _07428_, _07422_);
  and (_07430_, _07429_, _03401_);
  and (_07431_, _07430_, _07412_);
  or (_07432_, _07431_, _07409_);
  and (_07433_, _02798_, _02949_);
  nor (_07434_, _03028_, _02541_);
  nor (_07435_, _07434_, _02600_);
  or (_07436_, _07435_, _03394_);
  nor (_07437_, _07436_, _07433_);
  and (_07438_, _07437_, _07432_);
  nor (_07439_, _02538_, _02305_);
  and (_07440_, _07439_, _02949_);
  or (_07441_, _07440_, _07433_);
  and (_07442_, _07441_, xram_data_in_reg[7]);
  or (_07443_, _07442_, _02948_);
  or (_07444_, _07443_, _07438_);
  and (_07445_, _07444_, _07408_);
  or (_07446_, _07445_, _07405_);
  nor (_07447_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07448_, _07447_, _02625_);
  and (_07449_, _07448_, _06825_);
  and (_07450_, _07449_, \oc8051_golden_model_1.ACC [6]);
  and (_07451_, _07450_, \oc8051_golden_model_1.ACC [7]);
  nor (_07452_, _07450_, \oc8051_golden_model_1.ACC [7]);
  nor (_07453_, _07452_, _07451_);
  and (_07454_, _07448_, \oc8051_golden_model_1.ACC [4]);
  nor (_07455_, _07454_, \oc8051_golden_model_1.ACC [5]);
  nor (_07456_, _07455_, _07449_);
  nor (_07457_, _07449_, \oc8051_golden_model_1.ACC [6]);
  nor (_07458_, _07457_, _07450_);
  nor (_07459_, _07458_, _07456_);
  not (_07460_, _07459_);
  and (_07461_, _07460_, _07453_);
  nor (_07462_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_07463_, _07462_, _07459_);
  nor (_07464_, _07463_, _07453_);
  nor (_07465_, _07464_, _07461_);
  not (_07466_, _07465_);
  nand (_07467_, _07466_, _07405_);
  and (_07468_, _07467_, _02976_);
  and (_07469_, _07468_, _07446_);
  nor (_07470_, _05313_, _05364_);
  and (_07471_, _05348_, _05313_);
  nor (_07472_, _07471_, _07470_);
  nor (_07473_, _07472_, _02934_);
  not (_07474_, _02946_);
  nor (_07475_, _07321_, _07474_);
  or (_07476_, _07475_, _07403_);
  or (_07477_, _07476_, _07473_);
  or (_07478_, _07477_, _07469_);
  and (_07479_, _07478_, _07404_);
  or (_07480_, _07479_, _03873_);
  not (_07481_, _03873_);
  or (_07482_, _05461_, _07481_);
  and (_07483_, _07482_, _02992_);
  and (_07484_, _07483_, _07480_);
  and (_07485_, _03028_, _02875_);
  nor (_07486_, _05497_, _02992_);
  or (_07487_, _07486_, _07485_);
  or (_07488_, _07487_, _07484_);
  nand (_07489_, _07485_, _02625_);
  and (_07490_, _07489_, _07488_);
  or (_07491_, _07490_, _02877_);
  and (_07492_, _05344_, _05313_);
  nor (_07493_, _07492_, _07470_);
  nand (_07494_, _07493_, _02877_);
  and (_07495_, _07494_, _06246_);
  and (_07496_, _07495_, _07491_);
  and (_07497_, _07471_, _05502_);
  nor (_07498_, _07497_, _07470_);
  nor (_07499_, _07498_, _06246_);
  or (_07500_, _07499_, _06252_);
  or (_07501_, _07500_, _07496_);
  nor (_07502_, _06731_, _06729_);
  nor (_07503_, _07502_, _06732_);
  or (_07504_, _07503_, _06258_);
  and (_07505_, _07504_, _07501_);
  or (_07506_, _07505_, _07400_);
  not (_07507_, _07397_);
  not (_07508_, _07243_);
  and (_07509_, _07265_, _07257_);
  not (_07510_, _07509_);
  and (_07511_, _07280_, _07274_);
  nor (_07512_, _07290_, _02696_);
  nor (_07513_, _07512_, _07285_);
  or (_07514_, _07513_, _07286_);
  and (_07515_, _07514_, _07511_);
  not (_07516_, _07515_);
  and (_07517_, _07279_, _07274_);
  nor (_07518_, _07517_, _07273_);
  and (_07519_, _07518_, _07516_);
  and (_07520_, _07290_, _02696_);
  nor (_07521_, _07512_, _07520_);
  and (_07522_, _07521_, _07287_);
  and (_07523_, _07522_, _07511_);
  nor (_07524_, _07523_, _07519_);
  nor (_07525_, _07524_, _07510_);
  not (_07526_, _07525_);
  and (_07527_, _07263_, _07257_);
  nor (_07528_, _07527_, _07256_);
  and (_07529_, _07528_, _07526_);
  nor (_07530_, _07529_, _07248_);
  or (_07531_, _07530_, _07249_);
  and (_07532_, _07531_, _07508_);
  nor (_07533_, _07531_, _07508_);
  or (_07534_, _07533_, _07532_);
  or (_07535_, _07534_, _07399_);
  and (_07536_, _07535_, _07507_);
  and (_07537_, _07536_, _07506_);
  or (_07538_, _07537_, _02979_);
  or (_07539_, _07538_, _07398_);
  and (_07540_, _03028_, _02864_);
  not (_07541_, _07540_);
  and (_07542_, _04666_, \oc8051_golden_model_1.P2INREG [6]);
  and (_07543_, _04670_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_07544_, _07543_, _07542_);
  and (_07545_, _04654_, \oc8051_golden_model_1.P0INREG [6]);
  and (_07546_, _04660_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_07547_, _07546_, _07545_);
  and (_07548_, _07547_, _07544_);
  and (_07549_, _07548_, _04826_);
  and (_07550_, _07549_, _04817_);
  and (_07551_, _07550_, _04811_);
  and (_07552_, _07551_, _04791_);
  not (_07553_, _07552_);
  and (_07554_, _04654_, \oc8051_golden_model_1.P0INREG [3]);
  not (_07555_, _07554_);
  and (_07556_, _04660_, \oc8051_golden_model_1.P1INREG [3]);
  not (_07557_, _07556_);
  and (_07558_, _04666_, \oc8051_golden_model_1.P2INREG [3]);
  and (_07559_, _04670_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_07560_, _07559_, _07558_);
  and (_07561_, _07560_, _07557_);
  and (_07562_, _07561_, _04981_);
  and (_07563_, _07562_, _07555_);
  and (_07564_, _07563_, _04972_);
  and (_07565_, _07564_, _04966_);
  and (_07566_, _07565_, _04946_);
  not (_07567_, _07566_);
  and (_07568_, _04666_, \oc8051_golden_model_1.P2INREG [2]);
  and (_07569_, _04670_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_07570_, _07569_, _07568_);
  and (_07571_, _04654_, \oc8051_golden_model_1.P0INREG [2]);
  and (_07572_, _04660_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_07573_, _07572_, _07571_);
  and (_07574_, _07573_, _07570_);
  and (_07575_, _07574_, _05122_);
  and (_07576_, _07575_, _05112_);
  and (_07577_, _07576_, _05087_);
  not (_07578_, _07577_);
  not (_07579_, _05011_);
  nor (_07580_, _05015_, _05012_);
  and (_07581_, _07580_, _05023_);
  and (_07582_, _07581_, _07579_);
  and (_07583_, _07582_, _05034_);
  and (_07584_, _05020_, _04999_);
  and (_07585_, _04666_, \oc8051_golden_model_1.P2INREG [1]);
  and (_07586_, _04670_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_07587_, _07586_, _07585_);
  and (_07588_, _04660_, \oc8051_golden_model_1.P1INREG [1]);
  and (_07589_, _04654_, \oc8051_golden_model_1.P0INREG [1]);
  nor (_07590_, _07589_, _07588_);
  and (_07591_, _07590_, _07587_);
  and (_07592_, _07591_, _05010_);
  and (_07593_, _07592_, _07584_);
  and (_07594_, _07593_, _07583_);
  and (_07595_, _07594_, _04994_);
  not (_07596_, _07595_);
  and (_07597_, _04666_, \oc8051_golden_model_1.P2INREG [0]);
  and (_07598_, _04670_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_07599_, _07598_, _07597_);
  and (_07600_, _04654_, \oc8051_golden_model_1.P0INREG [0]);
  and (_07601_, _04660_, \oc8051_golden_model_1.P1INREG [0]);
  nor (_07602_, _07601_, _07600_);
  and (_07603_, _07602_, _07599_);
  and (_07604_, _07603_, _05074_);
  and (_07605_, _07604_, _05065_);
  and (_07606_, _07605_, _05059_);
  and (_07607_, _07606_, _05039_);
  nor (_07608_, _07607_, _07288_);
  and (_07609_, _07608_, _07596_);
  and (_07610_, _07609_, _07578_);
  and (_07611_, _07610_, _07567_);
  and (_07612_, _04666_, \oc8051_golden_model_1.P2INREG [5]);
  and (_07613_, _04670_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_07614_, _07613_, _07612_);
  and (_07615_, _04654_, \oc8051_golden_model_1.P0INREG [5]);
  and (_07616_, _04660_, \oc8051_golden_model_1.P1INREG [5]);
  nor (_07617_, _07616_, _07615_);
  and (_07618_, _07617_, _07614_);
  and (_07619_, _07618_, _04901_);
  and (_07620_, _07619_, _04942_);
  and (_07621_, _07620_, _04895_);
  not (_07622_, _05213_);
  nor (_07623_, _05217_, _05214_);
  and (_07624_, _07623_, _05225_);
  and (_07625_, _07624_, _07622_);
  and (_07626_, _07625_, _05236_);
  and (_07627_, _05222_, _05204_);
  and (_07628_, _04666_, \oc8051_golden_model_1.P2INREG [4]);
  and (_07629_, _04670_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_07630_, _07629_, _07628_);
  and (_07631_, _04660_, \oc8051_golden_model_1.P1INREG [4]);
  and (_07632_, _04654_, \oc8051_golden_model_1.P0INREG [4]);
  nor (_07633_, _07632_, _07631_);
  and (_07634_, _07633_, _07630_);
  and (_07635_, _07634_, _05212_);
  and (_07636_, _07635_, _07627_);
  and (_07637_, _07636_, _07626_);
  and (_07638_, _07637_, _05193_);
  nor (_07639_, _07638_, _07621_);
  and (_07640_, _07639_, _07611_);
  and (_07641_, _07640_, _07553_);
  nor (_07642_, _07641_, _05497_);
  and (_07643_, _07641_, _05497_);
  nor (_07644_, _07643_, _07642_);
  and (_07645_, _07644_, \oc8051_golden_model_1.ACC [7]);
  nor (_07646_, _07644_, \oc8051_golden_model_1.ACC [7]);
  nor (_07647_, _07646_, _07645_);
  not (_07648_, _07647_);
  nor (_07649_, _07640_, _07553_);
  nor (_07650_, _07649_, _07641_);
  nor (_07651_, _07650_, _06807_);
  and (_07652_, _07650_, _06807_);
  not (_07653_, _07621_);
  not (_07654_, _07638_);
  and (_07655_, _07611_, _07654_);
  nor (_07656_, _07655_, _07653_);
  nor (_07657_, _07656_, _07640_);
  and (_07658_, _07657_, _06858_);
  nor (_07659_, _07657_, _06858_);
  nor (_07660_, _07611_, _07654_);
  nor (_07661_, _07660_, _07655_);
  nor (_07662_, _07661_, _06864_);
  nor (_07663_, _07662_, _07659_);
  nor (_07664_, _07663_, _07658_);
  nor (_07665_, _07659_, _07658_);
  and (_07666_, _07661_, _06864_);
  nor (_07667_, _07666_, _07662_);
  and (_07668_, _07667_, _07665_);
  not (_07669_, _07668_);
  nor (_07670_, _07610_, _07567_);
  nor (_07671_, _07670_, _07611_);
  nor (_07672_, _07671_, _02625_);
  and (_07673_, _07671_, _02625_);
  nor (_07674_, _07673_, _07672_);
  nor (_07675_, _07609_, _07578_);
  nor (_07676_, _07675_, _07610_);
  nor (_07677_, _07676_, _06964_);
  and (_07678_, _07676_, _06964_);
  nor (_07679_, _07678_, _07677_);
  and (_07680_, _07679_, _07674_);
  not (_07681_, _07680_);
  nor (_07682_, _07608_, _07596_);
  nor (_07683_, _07682_, _07609_);
  and (_07684_, _07683_, _02543_);
  nor (_07685_, _07683_, _02543_);
  and (_07686_, _07607_, _07288_);
  nor (_07687_, _07686_, _07608_);
  nor (_07688_, _07687_, _02696_);
  nor (_07689_, _07688_, _07685_);
  nor (_07690_, _07689_, _07684_);
  nor (_07691_, _07690_, _07681_);
  nor (_07692_, _07678_, _07673_);
  or (_07693_, _07692_, _07672_);
  not (_07694_, _07693_);
  nor (_07695_, _07694_, _07691_);
  and (_07696_, _07687_, _02696_);
  nor (_07697_, _07688_, _07696_);
  nor (_07698_, _07595_, \oc8051_golden_model_1.ACC [1]);
  and (_07699_, _07595_, \oc8051_golden_model_1.ACC [1]);
  nor (_07700_, _07699_, _07698_);
  and (_07701_, \oc8051_golden_model_1.PSW [7], _02696_);
  and (_07702_, _07288_, \oc8051_golden_model_1.ACC [0]);
  nor (_07703_, _07607_, _07702_);
  nor (_07704_, _07703_, _07701_);
  and (_07705_, _07704_, _07700_);
  nor (_07706_, _07704_, _07700_);
  or (_07707_, _07706_, _07705_);
  nand (_07708_, _07707_, _07697_);
  nor (_07709_, _07708_, _07681_);
  nor (_07710_, _07709_, _07695_);
  nor (_07711_, _07710_, _07669_);
  nor (_07712_, _07711_, _07664_);
  nor (_07713_, _07712_, _07652_);
  or (_07714_, _07713_, _07651_);
  nand (_07715_, _07714_, _07648_);
  or (_07716_, _07714_, _07648_);
  and (_07717_, _07716_, _07715_);
  nand (_07718_, _07717_, _02979_);
  and (_07719_, _07718_, _07541_);
  and (_07720_, _07719_, _07539_);
  not (_07721_, _02571_);
  and (_07722_, _04677_, \oc8051_golden_model_1.PSW [7]);
  and (_07723_, _07722_, _04683_);
  and (_07724_, _07723_, _04668_);
  and (_07725_, _07724_, _04374_);
  nor (_07726_, _07725_, _02763_);
  and (_07727_, _07724_, _02925_);
  nor (_07728_, _07727_, _07726_);
  and (_07729_, _07728_, \oc8051_golden_model_1.ACC [7]);
  nor (_07730_, _07728_, \oc8051_golden_model_1.ACC [7]);
  nor (_07731_, _07730_, _07729_);
  not (_07732_, _07731_);
  nor (_07733_, _07724_, _04374_);
  nor (_07734_, _07733_, _07725_);
  nor (_07735_, _07734_, _06807_);
  and (_07736_, _07734_, _06807_);
  and (_07737_, _07723_, _04657_);
  nor (_07738_, _07737_, _04663_);
  nor (_07739_, _07738_, _07724_);
  and (_07740_, _07739_, _06858_);
  nor (_07741_, _07739_, _06858_);
  nor (_07742_, _07723_, _04657_);
  nor (_07743_, _07742_, _07737_);
  nor (_07744_, _07743_, _06864_);
  nor (_07745_, _07744_, _07741_);
  nor (_07746_, _07745_, _07740_);
  nor (_07747_, _07741_, _07740_);
  and (_07748_, _07743_, _06864_);
  nor (_07749_, _07748_, _07744_);
  and (_07750_, _07749_, _07747_);
  not (_07751_, _07750_);
  nor (_07752_, _05530_, _02794_);
  nor (_07753_, _07752_, _07723_);
  nor (_07754_, _07753_, _02625_);
  and (_07755_, _07753_, _02625_);
  nor (_07756_, _07755_, _07754_);
  nor (_07757_, _07722_, _04385_);
  nor (_07758_, _07757_, _05530_);
  nor (_07759_, _07758_, _06964_);
  and (_07760_, _07758_, _06964_);
  nor (_07761_, _07760_, _07759_);
  and (_07762_, _07761_, _07756_);
  and (_07763_, _02833_, \oc8051_golden_model_1.PSW [7]);
  nor (_07764_, _07763_, _03951_);
  nor (_07765_, _07764_, _07722_);
  and (_07766_, _07765_, _02543_);
  nor (_07767_, _07765_, _02543_);
  and (_07768_, _02837_, _07288_);
  nor (_07769_, _07768_, _07763_);
  nor (_07770_, _07769_, _02696_);
  nor (_07771_, _07770_, _07767_);
  or (_07772_, _07771_, _07766_);
  and (_07773_, _07772_, _07762_);
  not (_07774_, _07773_);
  and (_07775_, _07760_, _07756_);
  nor (_07776_, _07775_, _07755_);
  and (_07777_, _07776_, _07774_);
  not (_07778_, _07762_);
  and (_07779_, _07769_, _02696_);
  nor (_07780_, _07770_, _07779_);
  nor (_07781_, _03687_, _02543_);
  and (_07782_, _03687_, _02543_);
  or (_07783_, _07782_, _07781_);
  not (_07784_, _07702_);
  and (_07785_, _07784_, _02833_);
  nor (_07786_, _07785_, _07701_);
  and (_07787_, _07786_, _07783_);
  nor (_07788_, _07786_, _07783_);
  or (_07789_, _07788_, _07787_);
  nand (_07790_, _07789_, _07780_);
  nor (_07791_, _07790_, _07778_);
  nor (_07792_, _07791_, _07777_);
  nor (_07793_, _07792_, _07751_);
  nor (_07794_, _07793_, _07746_);
  nor (_07795_, _07794_, _07736_);
  or (_07796_, _07795_, _07735_);
  and (_07797_, _07796_, _07732_);
  nor (_07798_, _07796_, _07732_);
  or (_07799_, _07798_, _07797_);
  and (_07800_, _07799_, _07540_);
  or (_07801_, _07800_, _07721_);
  or (_07802_, _07801_, _07720_);
  nand (_07803_, _02763_, _07721_);
  and (_07804_, _07803_, _02986_);
  and (_07805_, _07804_, _07802_);
  not (_07806_, _05313_);
  nor (_07807_, _05531_, _07806_);
  nor (_07808_, _07807_, _07470_);
  nor (_07809_, _07808_, _02986_);
  or (_07810_, _07809_, _05535_);
  or (_07811_, _07810_, _07805_);
  and (_07812_, _07811_, _07322_);
  or (_07813_, _07812_, _02841_);
  and (_07814_, _05461_, _04731_);
  or (_07815_, _07814_, _07315_);
  or (_07816_, _07815_, _02842_);
  and (_07817_, _07816_, _02839_);
  and (_07818_, _07817_, _07813_);
  nor (_07819_, _05740_, _07319_);
  nor (_07820_, _07819_, _07315_);
  nor (_07821_, _07820_, _02839_);
  or (_07822_, _07821_, _06786_);
  or (_07823_, _07822_, _07818_);
  or (_07824_, _06805_, _06792_);
  and (_07825_, _07824_, _07823_);
  and (_07826_, _07825_, _02609_);
  nor (_07827_, _02763_, _02609_);
  or (_07828_, _07827_, _02834_);
  or (_07829_, _07828_, _07826_);
  and (_07830_, _03028_, _02521_);
  not (_07831_, _07830_);
  and (_07832_, _05549_, _04731_);
  nor (_07833_, _07832_, _07315_);
  nand (_07834_, _07833_, _02834_);
  and (_07835_, _07834_, _07831_);
  and (_07836_, _07835_, _07829_);
  nor (_07837_, _07831_, _02763_);
  nand (_07838_, _07231_, _02523_);
  and (_07839_, _02854_, _02523_);
  or (_07840_, _07839_, _03517_);
  and (_07841_, _03009_, _02523_);
  nor (_07842_, _07841_, _03281_);
  not (_07843_, _07842_);
  nor (_07844_, _07843_, _07840_);
  and (_07845_, _07844_, _07838_);
  not (_07846_, _07845_);
  or (_07847_, _07846_, _07837_);
  or (_07848_, _07847_, _07836_);
  and (_07849_, _02840_, _02523_);
  not (_07850_, _07849_);
  or (_07851_, _07845_, _07192_);
  and (_07852_, _07851_, _07850_);
  and (_07853_, _07852_, _07848_);
  and (_07854_, _05810_, _05364_);
  and (_07855_, _05461_, \oc8051_golden_model_1.ACC [7]);
  nor (_07856_, _07855_, _07854_);
  and (_07857_, _07849_, _07856_);
  or (_07858_, _07857_, _03146_);
  or (_07859_, _07858_, _07853_);
  and (_07860_, _03028_, _02523_);
  not (_07861_, _07860_);
  or (_07862_, _05772_, _03147_);
  and (_07863_, _07862_, _07861_);
  and (_07864_, _07863_, _07859_);
  nor (_07865_, _02763_, _05364_);
  and (_07866_, _02763_, _05364_);
  nor (_07867_, _07866_, _07865_);
  and (_07868_, _07860_, _07867_);
  or (_07869_, _07868_, _03051_);
  or (_07870_, _07869_, _07864_);
  and (_07871_, _07870_, _07318_);
  or (_07872_, _07871_, _03148_);
  or (_07873_, _07315_, _07150_);
  and (_07874_, _02966_, _02529_);
  nor (_07875_, _07874_, _03764_);
  not (_07876_, _07875_);
  nor (_07877_, _07876_, _03758_);
  and (_07878_, _07877_, _07873_);
  and (_07879_, _07878_, _07872_);
  and (_07880_, _02849_, _02529_);
  not (_07881_, _07880_);
  and (_07882_, _07881_, _07875_);
  not (_07883_, _07882_);
  and (_07884_, _02845_, _02529_);
  or (_07885_, _07884_, _07191_);
  and (_07886_, _07885_, _07883_);
  or (_07887_, _07886_, _07879_);
  not (_07888_, _07884_);
  or (_07889_, _07888_, _07191_);
  and (_07890_, _02840_, _02529_);
  not (_07891_, _07890_);
  and (_07892_, _07891_, _07889_);
  and (_07893_, _07892_, _07887_);
  and (_07894_, _07890_, _07855_);
  or (_07895_, _07894_, _03135_);
  or (_07896_, _07895_, _07893_);
  and (_07897_, _07896_, _07314_);
  and (_07898_, _07865_, _07311_);
  or (_07899_, _07898_, _07897_);
  and (_07900_, _07899_, _03023_);
  or (_07901_, _07833_, _05771_);
  nor (_07902_, _07901_, _03023_);
  or (_07903_, _07902_, _07309_);
  or (_07904_, _07903_, _07900_);
  and (_07905_, _07904_, _07310_);
  nor (_07906_, _03019_, _03543_);
  or (_07907_, _07906_, _07905_);
  and (_07908_, _07231_, _02532_);
  and (_07909_, _02962_, _02532_);
  or (_07910_, _07190_, _07909_);
  nand (_07911_, _07910_, _07908_);
  and (_07912_, _07911_, _07907_);
  not (_07913_, _07909_);
  nor (_07914_, _07190_, _07913_);
  and (_07915_, _02840_, _02532_);
  or (_07916_, _07915_, _07914_);
  or (_07917_, _07916_, _07912_);
  nand (_07918_, _07915_, _07854_);
  and (_07919_, _07918_, _03142_);
  and (_07920_, _07919_, _07917_);
  and (_07921_, _03028_, _02532_);
  nor (_07922_, _05771_, _03142_);
  or (_07923_, _07922_, _07921_);
  or (_07924_, _07923_, _07920_);
  nand (_07925_, _07921_, _07866_);
  and (_07926_, _07925_, _03043_);
  and (_07927_, _07926_, _07924_);
  nor (_07928_, _05763_, _07319_);
  nor (_07929_, _07928_, _07315_);
  nor (_07930_, _07929_, _03043_);
  not (_07931_, _07234_);
  or (_07932_, _07931_, _07930_);
  or (_07933_, _07932_, _07927_);
  and (_07934_, _07933_, _07308_);
  or (_07935_, _07934_, _07229_);
  not (_07936_, _07229_);
  and (_07937_, _07334_, \oc8051_golden_model_1.ACC [6]);
  nor (_07938_, _07335_, _07336_);
  and (_07939_, _07340_, \oc8051_golden_model_1.ACC [5]);
  and (_07940_, _07346_, \oc8051_golden_model_1.ACC [4]);
  and (_07941_, _07358_, \oc8051_golden_model_1.ACC [3]);
  and (_07942_, _07363_, \oc8051_golden_model_1.ACC [2]);
  and (_07943_, _07370_, \oc8051_golden_model_1.ACC [1]);
  and (_07944_, _07374_, \oc8051_golden_model_1.ACC [0]);
  not (_07945_, _07944_);
  nor (_07946_, _07945_, _07384_);
  nor (_07947_, _07946_, _07943_);
  nor (_07948_, _07947_, _07366_);
  nor (_07949_, _07948_, _07942_);
  nor (_07950_, _07949_, _07361_);
  nor (_07951_, _07950_, _07941_);
  nor (_07952_, _07951_, _07352_);
  nor (_07953_, _07952_, _07940_);
  nor (_07954_, _07953_, _07350_);
  nor (_07955_, _07954_, _07939_);
  nor (_07956_, _07955_, _07938_);
  nor (_07957_, _07956_, _07937_);
  nor (_07958_, _07957_, _07331_);
  and (_07959_, _07957_, _07331_);
  nor (_07960_, _07959_, _07958_);
  or (_07961_, _07960_, _07936_);
  and (_07962_, _07961_, _03134_);
  and (_07963_, _07962_, _07935_);
  and (_07964_, _03028_, _02527_);
  nor (_07965_, _07964_, _03133_);
  not (_07966_, _07965_);
  and (_07967_, _07650_, \oc8051_golden_model_1.ACC [6]);
  nor (_07968_, _07651_, _07652_);
  and (_07969_, _07657_, \oc8051_golden_model_1.ACC [5]);
  and (_07970_, _07661_, \oc8051_golden_model_1.ACC [4]);
  and (_07971_, _07671_, \oc8051_golden_model_1.ACC [3]);
  and (_07972_, _07676_, \oc8051_golden_model_1.ACC [2]);
  and (_07973_, _07683_, \oc8051_golden_model_1.ACC [1]);
  nor (_07974_, _07685_, _07684_);
  and (_07975_, _07687_, \oc8051_golden_model_1.ACC [0]);
  not (_07976_, _07975_);
  nor (_07977_, _07976_, _07974_);
  nor (_07978_, _07977_, _07973_);
  nor (_07979_, _07978_, _07679_);
  nor (_07980_, _07979_, _07972_);
  nor (_07981_, _07980_, _07674_);
  nor (_07982_, _07981_, _07971_);
  nor (_07983_, _07982_, _07667_);
  nor (_07984_, _07983_, _07970_);
  nor (_07985_, _07984_, _07665_);
  nor (_07986_, _07985_, _07969_);
  nor (_07987_, _07986_, _07968_);
  nor (_07988_, _07987_, _07967_);
  nor (_07989_, _07988_, _07647_);
  and (_07990_, _07988_, _07647_);
  nor (_07991_, _07990_, _07989_);
  or (_07992_, _07991_, _07964_);
  and (_07993_, _07992_, _07966_);
  or (_07994_, _07993_, _07963_);
  and (_07995_, _02541_, _02527_);
  not (_07996_, _07995_);
  not (_07997_, _07964_);
  and (_07998_, _07734_, \oc8051_golden_model_1.ACC [6]);
  nor (_07999_, _07735_, _07736_);
  and (_08000_, _07739_, \oc8051_golden_model_1.ACC [5]);
  and (_08001_, _07743_, \oc8051_golden_model_1.ACC [4]);
  and (_08002_, _07753_, \oc8051_golden_model_1.ACC [3]);
  and (_08003_, _07758_, \oc8051_golden_model_1.ACC [2]);
  and (_08004_, _07765_, \oc8051_golden_model_1.ACC [1]);
  nor (_08005_, _07766_, _07767_);
  and (_08006_, _07769_, \oc8051_golden_model_1.ACC [0]);
  not (_08007_, _08006_);
  nor (_08008_, _08007_, _08005_);
  nor (_08009_, _08008_, _08004_);
  nor (_08010_, _08009_, _07761_);
  nor (_08011_, _08010_, _08003_);
  nor (_08012_, _08011_, _07756_);
  nor (_08013_, _08012_, _08002_);
  nor (_08014_, _08013_, _07749_);
  nor (_08015_, _08014_, _08001_);
  nor (_08016_, _08015_, _07747_);
  nor (_08017_, _08016_, _08000_);
  nor (_08018_, _08017_, _07999_);
  nor (_08019_, _08018_, _07998_);
  nor (_08020_, _08019_, _07731_);
  and (_08021_, _08019_, _07731_);
  nor (_08022_, _08021_, _08020_);
  or (_08023_, _08022_, _07997_);
  and (_08024_, _08023_, _07996_);
  and (_08025_, _08024_, _07994_);
  nand (_08026_, _07995_, \oc8051_golden_model_1.ACC [6]);
  nand (_08027_, _07189_, _08026_);
  or (_08028_, _08027_, _08025_);
  and (_08029_, _08028_, _07228_);
  or (_08030_, _08029_, _07185_);
  not (_08031_, _07185_);
  and (_08032_, _06162_, \oc8051_golden_model_1.ACC [6]);
  and (_08033_, _05855_, _06807_);
  nor (_08034_, _08032_, _08033_);
  and (_08035_, _06170_, \oc8051_golden_model_1.ACC [5]);
  and (_08036_, _06083_, _06858_);
  nor (_08037_, _08036_, _08035_);
  not (_08038_, _08037_);
  and (_08039_, _06171_, \oc8051_golden_model_1.ACC [4]);
  and (_08040_, _06128_, _06864_);
  nor (_08041_, _08039_, _08040_);
  and (_08042_, _06166_, \oc8051_golden_model_1.ACC [3]);
  and (_08043_, _05991_, _02625_);
  and (_08044_, _06167_, \oc8051_golden_model_1.ACC [2]);
  and (_08045_, _06036_, _06964_);
  nor (_08046_, _08044_, _08045_);
  not (_08047_, _08046_);
  and (_08048_, _06163_, \oc8051_golden_model_1.ACC [1]);
  and (_08049_, _05900_, _02543_);
  nor (_08050_, _08048_, _08049_);
  and (_08051_, _06164_, \oc8051_golden_model_1.ACC [0]);
  and (_08052_, _08051_, _08050_);
  nor (_08053_, _08052_, _08048_);
  nor (_08054_, _08053_, _08047_);
  nor (_08055_, _08054_, _08044_);
  nor (_08056_, _08055_, _08043_);
  or (_08057_, _08056_, _08042_);
  and (_08058_, _08057_, _08041_);
  nor (_08059_, _08058_, _08039_);
  nor (_08060_, _08059_, _08038_);
  or (_08061_, _08060_, _08035_);
  and (_08062_, _08061_, _08034_);
  nor (_08063_, _08062_, _08032_);
  nor (_08064_, _08063_, _07856_);
  and (_08065_, _08063_, _07856_);
  or (_08066_, _08065_, _08064_);
  or (_08067_, _08066_, _08031_);
  and (_08068_, _08067_, _03166_);
  and (_08069_, _08068_, _08030_);
  and (_08070_, _03028_, _02509_);
  and (_08071_, _05497_, _05364_);
  nor (_08072_, _05497_, _05364_);
  nor (_08073_, _08072_, _08071_);
  nor (_08074_, _07552_, _06807_);
  and (_08075_, _07552_, \oc8051_golden_model_1.ACC [6]);
  nor (_08076_, _07552_, \oc8051_golden_model_1.ACC [6]);
  nor (_08077_, _08076_, _08075_);
  nor (_08078_, _07621_, _06858_);
  nor (_08079_, _07621_, \oc8051_golden_model_1.ACC [5]);
  and (_08080_, _07621_, \oc8051_golden_model_1.ACC [5]);
  nor (_08081_, _08080_, _08079_);
  nor (_08082_, _07638_, _06864_);
  and (_08083_, _07638_, \oc8051_golden_model_1.ACC [4]);
  nor (_08084_, _07638_, \oc8051_golden_model_1.ACC [4]);
  nor (_08085_, _08084_, _08083_);
  not (_08086_, _08085_);
  nor (_08087_, _07577_, _06964_);
  and (_08088_, _07577_, \oc8051_golden_model_1.ACC [2]);
  nor (_08089_, _07577_, \oc8051_golden_model_1.ACC [2]);
  nor (_08090_, _08089_, _08088_);
  nor (_08091_, _07595_, _02543_);
  nor (_08092_, _07607_, _02696_);
  not (_08093_, _08092_);
  nor (_08094_, _08093_, _07700_);
  nor (_08095_, _08094_, _08091_);
  nor (_08096_, _08095_, _08090_);
  nor (_08097_, _08096_, _08087_);
  nor (_08098_, _08097_, _07566_);
  or (_08099_, _08098_, \oc8051_golden_model_1.ACC [3]);
  nand (_08100_, _08097_, _07566_);
  and (_08101_, _08100_, _08099_);
  and (_08102_, _08101_, _08086_);
  nor (_08103_, _08102_, _08082_);
  nor (_08104_, _08103_, _08081_);
  nor (_08105_, _08104_, _08078_);
  nor (_08106_, _08105_, _08077_);
  nor (_08107_, _08106_, _08074_);
  nor (_08108_, _08107_, _08073_);
  and (_08109_, _08107_, _08073_);
  or (_08110_, _08109_, _08108_);
  or (_08111_, _08110_, _08070_);
  or (_08112_, _08070_, _02892_);
  and (_08113_, _08112_, _08111_);
  or (_08114_, _08113_, _08069_);
  and (_08115_, _02541_, _02509_);
  not (_08116_, _08115_);
  not (_08117_, _08070_);
  nor (_08118_, _02924_, _06807_);
  and (_08119_, _02924_, _06807_);
  nor (_08120_, _08119_, _08118_);
  nor (_08121_, _03220_, _06858_);
  and (_08122_, _03220_, _06858_);
  nor (_08123_, _03647_, _06864_);
  and (_08124_, _03647_, _06864_);
  nor (_08125_, _08124_, _08123_);
  and (_08126_, _02794_, \oc8051_golden_model_1.ACC [3]);
  nor (_08127_, _02794_, \oc8051_golden_model_1.ACC [3]);
  nor (_08128_, _03356_, _06964_);
  and (_08129_, _03356_, _06964_);
  nor (_08130_, _08129_, _08128_);
  not (_08131_, _08130_);
  and (_08132_, _02833_, \oc8051_golden_model_1.ACC [0]);
  not (_08133_, _08132_);
  nor (_08134_, _07783_, _08133_);
  nor (_08135_, _08134_, _07781_);
  nor (_08136_, _08135_, _08131_);
  nor (_08137_, _08136_, _08128_);
  nor (_08138_, _08137_, _08127_);
  or (_08139_, _08138_, _08126_);
  and (_08140_, _08139_, _08125_);
  nor (_08141_, _08140_, _08123_);
  nor (_08142_, _08141_, _08122_);
  or (_08143_, _08142_, _08121_);
  and (_08144_, _08143_, _08120_);
  nor (_08145_, _08144_, _08118_);
  nor (_08146_, _08145_, _07867_);
  and (_08147_, _08145_, _07867_);
  or (_08148_, _08147_, _08146_);
  or (_08149_, _08148_, _08117_);
  and (_08150_, _08149_, _08116_);
  and (_08151_, _08150_, _08114_);
  and (_08152_, _08115_, \oc8051_golden_model_1.ACC [6]);
  or (_08153_, _08152_, _03174_);
  or (_08154_, _08153_, _08151_);
  and (_08155_, _03028_, _02504_);
  not (_08156_, _08155_);
  nand (_08157_, _07407_, _03174_);
  and (_08158_, _08157_, _08156_);
  and (_08159_, _08158_, _08154_);
  and (_08160_, _02541_, _02504_);
  nor (_08161_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08162_, _08161_, _06904_);
  and (_08163_, _08162_, _06824_);
  and (_08164_, _08163_, _06807_);
  nor (_08165_, _08164_, _05364_);
  and (_08166_, _08164_, _05364_);
  nor (_08167_, _08166_, _08165_);
  nor (_08168_, _08167_, _08156_);
  or (_08169_, _08168_, _08160_);
  or (_08170_, _08169_, _08159_);
  nand (_08171_, _08160_, _07288_);
  and (_08172_, _08171_, _03183_);
  and (_08173_, _08172_, _08170_);
  nor (_08174_, _07493_, _03183_);
  or (_08175_, _08174_, _02887_);
  or (_08176_, _08175_, _08173_);
  and (_08177_, _03028_, _02498_);
  not (_08178_, _08177_);
  and (_08179_, _05246_, _04731_);
  nor (_08180_, _08179_, _07315_);
  nand (_08181_, _08180_, _02887_);
  and (_08182_, _08181_, _08178_);
  and (_08183_, _08182_, _08176_);
  and (_08184_, _02541_, _02498_);
  and (_08185_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08186_, _08185_, _06905_);
  nor (_08187_, _08186_, _06864_);
  and (_08188_, _08187_, \oc8051_golden_model_1.ACC [5]);
  and (_08189_, _08188_, \oc8051_golden_model_1.ACC [6]);
  nor (_08190_, _08189_, \oc8051_golden_model_1.ACC [7]);
  and (_08191_, _08189_, \oc8051_golden_model_1.ACC [7]);
  nor (_08192_, _08191_, _08190_);
  and (_08193_, _08192_, _08177_);
  or (_08194_, _08193_, _08184_);
  or (_08195_, _08194_, _08183_);
  nand (_08196_, _08184_, _02696_);
  and (_08197_, _08196_, _34655_);
  and (_08198_, _08197_, _08195_);
  or (_08199_, _08198_, _07184_);
  and (_35827_[7], _08199_, _35796_);
  not (_08200_, \oc8051_golden_model_1.DPL [7]);
  nor (_08201_, _34655_, _08200_);
  nor (_08202_, _04643_, _08200_);
  not (_08203_, _04643_);
  nor (_08204_, _05771_, _08203_);
  or (_08205_, _08204_, _08202_);
  and (_08206_, _08205_, _03143_);
  not (_08207_, _03052_);
  nor (_08208_, _08203_, _04630_);
  or (_08209_, _08208_, _08202_);
  or (_08210_, _08209_, _02859_);
  not (_08211_, _03046_);
  and (_08212_, _05474_, _04643_);
  or (_08213_, _08212_, _08202_);
  or (_08214_, _08213_, _03006_);
  and (_08215_, _04643_, \oc8051_golden_model_1.ACC [7]);
  or (_08216_, _08215_, _08202_);
  and (_08217_, _08216_, _03845_);
  nor (_08218_, _03845_, _08200_);
  or (_08219_, _08218_, _02948_);
  or (_08220_, _08219_, _08217_);
  and (_08221_, _08220_, _07474_);
  and (_08222_, _08221_, _08214_);
  and (_08223_, _08209_, _02946_);
  or (_08224_, _08223_, _02880_);
  or (_08225_, _08224_, _08222_);
  nor (_08226_, _02588_, _02540_);
  not (_08227_, _08226_);
  or (_08228_, _08216_, _02992_);
  and (_08229_, _08228_, _08227_);
  and (_08230_, _08229_, _08225_);
  and (_08231_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_08232_, _08231_, \oc8051_golden_model_1.DPL [2]);
  and (_08233_, _08232_, \oc8051_golden_model_1.DPL [3]);
  and (_08234_, _08233_, \oc8051_golden_model_1.DPL [4]);
  and (_08235_, _08234_, \oc8051_golden_model_1.DPL [5]);
  and (_08236_, _08235_, \oc8051_golden_model_1.DPL [6]);
  nor (_08237_, _08236_, \oc8051_golden_model_1.DPL [7]);
  and (_08238_, _08236_, \oc8051_golden_model_1.DPL [7]);
  nor (_08239_, _08238_, _08237_);
  and (_08240_, _08239_, _08226_);
  or (_08241_, _08240_, _08230_);
  and (_08242_, _08241_, _08211_);
  nor (_08243_, _05302_, _08211_);
  or (_08244_, _08243_, _05535_);
  or (_08245_, _08244_, _08242_);
  and (_08246_, _08245_, _08210_);
  or (_08247_, _08246_, _02841_);
  and (_08248_, _05461_, _04643_);
  or (_08249_, _08202_, _02842_);
  or (_08250_, _08249_, _08248_);
  and (_08251_, _08250_, _02839_);
  and (_08252_, _08251_, _08247_);
  nor (_08253_, _05740_, _08203_);
  or (_08254_, _08253_, _08202_);
  and (_08255_, _08254_, _02567_);
  or (_08256_, _08255_, _08252_);
  or (_08257_, _08256_, _08207_);
  and (_08258_, _05764_, _04643_);
  or (_08259_, _08202_, _07139_);
  or (_08260_, _08259_, _08258_);
  and (_08261_, _05549_, _04643_);
  or (_08262_, _08261_, _08202_);
  or (_08263_, _08262_, _07140_);
  and (_08264_, _08263_, _07150_);
  and (_08265_, _08264_, _08260_);
  and (_08266_, _08265_, _08257_);
  and (_08267_, _05772_, _04643_);
  or (_08268_, _08267_, _08202_);
  and (_08269_, _08268_, _03148_);
  or (_08270_, _08269_, _08266_);
  and (_08271_, _08270_, _03138_);
  or (_08272_, _08202_, _04740_);
  and (_08273_, _08216_, _03137_);
  and (_08274_, _08262_, _03022_);
  or (_08275_, _08274_, _08273_);
  and (_08276_, _08275_, _08272_);
  or (_08277_, _08276_, _03042_);
  or (_08278_, _08277_, _08271_);
  nor (_08279_, _05763_, _08203_);
  or (_08280_, _08202_, _03043_);
  or (_08281_, _08280_, _08279_);
  and (_08282_, _08281_, _07161_);
  and (_08283_, _08282_, _08278_);
  or (_08284_, _08283_, _08206_);
  and (_08285_, _08284_, _03179_);
  and (_08286_, _08213_, _03174_);
  or (_08287_, _08286_, _02887_);
  or (_08288_, _08287_, _08285_);
  and (_08289_, _05246_, _04643_);
  or (_08290_, _08202_, _02888_);
  or (_08291_, _08290_, _08289_);
  and (_08292_, _08291_, _34655_);
  and (_08293_, _08292_, _08288_);
  or (_08294_, _08293_, _08201_);
  and (_35830_[7], _08294_, _35796_);
  not (_08295_, \oc8051_golden_model_1.DPH [7]);
  nor (_08296_, _34655_, _08295_);
  and (_08297_, _04677_, _04652_);
  and (_08298_, _08297_, _04634_);
  nor (_08299_, _08298_, _08295_);
  not (_08300_, _04696_);
  nor (_08301_, _05771_, _08300_);
  or (_08302_, _08301_, _08299_);
  and (_08303_, _08302_, _03143_);
  nor (_08304_, _08300_, _04630_);
  or (_08305_, _08304_, _08299_);
  or (_08306_, _08305_, _02859_);
  and (_08307_, _05474_, _04696_);
  or (_08308_, _08307_, _08299_);
  or (_08309_, _08308_, _03006_);
  and (_08310_, _08298_, \oc8051_golden_model_1.ACC [7]);
  or (_08311_, _08310_, _08299_);
  and (_08312_, _08311_, _03845_);
  nor (_08313_, _03845_, _08295_);
  or (_08314_, _08313_, _02948_);
  or (_08315_, _08314_, _08312_);
  and (_08316_, _08315_, _07474_);
  and (_08317_, _08316_, _08309_);
  and (_08318_, _08305_, _02946_);
  or (_08319_, _08318_, _02880_);
  or (_08320_, _08319_, _08317_);
  or (_08321_, _08311_, _02992_);
  and (_08322_, _08321_, _08227_);
  and (_08323_, _08322_, _08320_);
  and (_08324_, _08238_, \oc8051_golden_model_1.DPH [0]);
  and (_08325_, _08324_, \oc8051_golden_model_1.DPH [1]);
  and (_08326_, _08325_, \oc8051_golden_model_1.DPH [2]);
  and (_08327_, _08326_, \oc8051_golden_model_1.DPH [3]);
  and (_08328_, _08327_, \oc8051_golden_model_1.DPH [4]);
  and (_08329_, _08328_, \oc8051_golden_model_1.DPH [5]);
  and (_08330_, _08329_, \oc8051_golden_model_1.DPH [6]);
  nor (_08331_, _08330_, _08295_);
  and (_08332_, _08330_, _08295_);
  or (_08333_, _08332_, _08331_);
  and (_08334_, _08333_, _08226_);
  or (_08335_, _08334_, _08323_);
  and (_08336_, _08335_, _08211_);
  nor (_08337_, _08211_, _02763_);
  or (_08338_, _08337_, _05535_);
  or (_08339_, _08338_, _08336_);
  and (_08340_, _08339_, _08306_);
  or (_08341_, _08340_, _02841_);
  or (_08342_, _08299_, _02842_);
  and (_08343_, _05461_, _08298_);
  or (_08344_, _08343_, _08342_);
  and (_08345_, _08344_, _08341_);
  or (_08346_, _08345_, _02567_);
  nor (_08347_, _05740_, _08300_);
  or (_08348_, _08299_, _02839_);
  or (_08349_, _08348_, _08347_);
  and (_08350_, _08349_, _08346_);
  or (_08351_, _08350_, _08207_);
  and (_08352_, _05764_, _04696_);
  or (_08353_, _08299_, _07139_);
  or (_08354_, _08353_, _08352_);
  and (_08355_, _05549_, _08298_);
  or (_08356_, _08355_, _08299_);
  or (_08357_, _08356_, _07140_);
  and (_08358_, _08357_, _07150_);
  and (_08359_, _08358_, _08354_);
  and (_08360_, _08359_, _08351_);
  and (_08361_, _05772_, _04696_);
  or (_08362_, _08361_, _08299_);
  and (_08363_, _08362_, _03148_);
  or (_08364_, _08363_, _08360_);
  and (_08365_, _08364_, _03138_);
  or (_08366_, _08299_, _04740_);
  and (_08367_, _08311_, _03137_);
  and (_08368_, _08356_, _03022_);
  or (_08369_, _08368_, _08367_);
  and (_08370_, _08369_, _08366_);
  or (_08371_, _08370_, _03042_);
  or (_08372_, _08371_, _08365_);
  nor (_08373_, _05763_, _08300_);
  or (_08374_, _08299_, _03043_);
  or (_08375_, _08374_, _08373_);
  and (_08376_, _08375_, _07161_);
  and (_08377_, _08376_, _08372_);
  or (_08378_, _08377_, _08303_);
  and (_08379_, _08378_, _03179_);
  and (_08380_, _08308_, _03174_);
  or (_08381_, _08380_, _02887_);
  or (_08382_, _08381_, _08379_);
  and (_08383_, _05246_, _04696_);
  or (_08384_, _08299_, _02888_);
  or (_08385_, _08384_, _08383_);
  and (_08386_, _08385_, _34655_);
  and (_08387_, _08386_, _08382_);
  or (_08388_, _08387_, _08296_);
  and (_35829_[7], _08388_, _35796_);
  and (_35831_[7], \oc8051_golden_model_1.IE [7], _35796_);
  and (_35832_[7], \oc8051_golden_model_1.IP [7], _35796_);
  not (_08389_, \oc8051_golden_model_1.P0 [7]);
  nor (_08390_, _34655_, _08389_);
  or (_08391_, _08390_, rst);
  nor (_08392_, _04654_, _08389_);
  not (_08393_, _04654_);
  nor (_08394_, _08393_, _04630_);
  or (_08395_, _08394_, _08392_);
  or (_08396_, _08395_, _02859_);
  nor (_08397_, _04635_, _08389_);
  and (_08398_, _05348_, _04635_);
  or (_08399_, _08398_, _08397_);
  or (_08400_, _08397_, _05502_);
  and (_08401_, _08400_, _02871_);
  and (_08402_, _08401_, _08399_);
  and (_08403_, _05474_, _04654_);
  or (_08404_, _08403_, _08392_);
  or (_08405_, _08404_, _03006_);
  and (_08406_, _04654_, \oc8051_golden_model_1.ACC [7]);
  or (_08407_, _08406_, _08392_);
  and (_08408_, _08407_, _03845_);
  nor (_08409_, _03845_, _08389_);
  or (_08410_, _08409_, _02948_);
  or (_08411_, _08410_, _08408_);
  and (_08412_, _08411_, _02976_);
  and (_08413_, _08412_, _08405_);
  and (_08414_, _08395_, _02946_);
  and (_08415_, _08399_, _02884_);
  or (_08416_, _08415_, _08414_);
  or (_08417_, _08416_, _02880_);
  or (_08418_, _08417_, _08413_);
  or (_08419_, _08407_, _02992_);
  and (_08420_, _08419_, _08418_);
  or (_08421_, _08420_, _02877_);
  and (_08422_, _05344_, _04635_);
  or (_08423_, _08422_, _08397_);
  or (_08424_, _08423_, _02987_);
  and (_08425_, _08424_, _06246_);
  and (_08426_, _08425_, _08421_);
  or (_08427_, _08426_, _08402_);
  and (_08428_, _08427_, _02986_);
  or (_08429_, _05530_, _05344_);
  and (_08430_, _08429_, _04635_);
  or (_08431_, _08430_, _08397_);
  and (_08432_, _08431_, _02866_);
  or (_08433_, _08432_, _05535_);
  or (_08434_, _08433_, _08428_);
  and (_08435_, _08434_, _08396_);
  or (_08436_, _08435_, _02841_);
  and (_08437_, _05461_, _04654_);
  or (_08438_, _08392_, _02842_);
  or (_08439_, _08438_, _08437_);
  and (_08440_, _08439_, _02839_);
  and (_08441_, _08440_, _08436_);
  nor (_08442_, _05740_, _08393_);
  or (_08443_, _08442_, _08392_);
  and (_08444_, _08443_, _02567_);
  or (_08445_, _08444_, _08207_);
  or (_08446_, _08445_, _08441_);
  and (_08447_, _05764_, _04654_);
  or (_08448_, _08392_, _07139_);
  or (_08449_, _08448_, _08447_);
  and (_08450_, _05549_, _04654_);
  or (_08451_, _08450_, _08392_);
  or (_08452_, _08451_, _07140_);
  and (_08453_, _08452_, _07150_);
  and (_08454_, _08453_, _08449_);
  and (_08455_, _08454_, _08446_);
  and (_08456_, _05772_, _04654_);
  or (_08457_, _08456_, _08392_);
  and (_08458_, _08457_, _03148_);
  or (_08459_, _08458_, _08455_);
  and (_08460_, _08459_, _03138_);
  or (_08461_, _08392_, _04740_);
  and (_08462_, _08407_, _03137_);
  and (_08463_, _08451_, _03022_);
  or (_08464_, _08463_, _08462_);
  and (_08465_, _08464_, _08461_);
  or (_08466_, _08465_, _03042_);
  or (_08467_, _08466_, _08460_);
  nor (_08468_, _05763_, _08393_);
  or (_08469_, _08392_, _03043_);
  or (_08470_, _08469_, _08468_);
  and (_08471_, _08470_, _07161_);
  and (_08472_, _08471_, _08467_);
  nor (_08473_, _05771_, _08393_);
  or (_08474_, _08473_, _08392_);
  and (_08475_, _08474_, _03143_);
  or (_08476_, _08475_, _03174_);
  or (_08477_, _08476_, _08472_);
  or (_08478_, _08404_, _03179_);
  and (_08479_, _08478_, _03183_);
  and (_08480_, _08479_, _08477_);
  and (_08481_, _08423_, _02799_);
  or (_08482_, _08481_, _02887_);
  or (_08483_, _08482_, _08480_);
  and (_08484_, _05246_, _04654_);
  or (_08485_, _08392_, _02888_);
  or (_08486_, _08485_, _08484_);
  and (_08487_, _08486_, _34655_);
  and (_08488_, _08487_, _08483_);
  or (_35834_[7], _08488_, _08391_);
  not (_08489_, \oc8051_golden_model_1.P1 [7]);
  nor (_08490_, _34655_, _08489_);
  or (_08491_, _08490_, rst);
  nor (_08492_, _04660_, _08489_);
  not (_08493_, _04660_);
  nor (_08494_, _08493_, _04630_);
  or (_08495_, _08494_, _08492_);
  or (_08496_, _08495_, _02859_);
  nor (_08497_, _05332_, _08489_);
  and (_08498_, _05348_, _05332_);
  or (_08499_, _08498_, _08497_);
  or (_08500_, _08497_, _05502_);
  and (_08501_, _08500_, _02871_);
  and (_08502_, _08501_, _08499_);
  and (_08503_, _05474_, _04660_);
  or (_08504_, _08503_, _08492_);
  or (_08505_, _08504_, _03006_);
  and (_08506_, _04660_, \oc8051_golden_model_1.ACC [7]);
  or (_08507_, _08506_, _08492_);
  and (_08508_, _08507_, _03845_);
  nor (_08509_, _03845_, _08489_);
  or (_08510_, _08509_, _02948_);
  or (_08511_, _08510_, _08508_);
  and (_08512_, _08511_, _02976_);
  and (_08513_, _08512_, _08505_);
  and (_08514_, _08495_, _02946_);
  and (_08515_, _08499_, _02884_);
  or (_08516_, _08515_, _08514_);
  or (_08517_, _08516_, _02880_);
  or (_08518_, _08517_, _08513_);
  or (_08519_, _08507_, _02992_);
  and (_08520_, _08519_, _08518_);
  or (_08521_, _08520_, _02877_);
  and (_08522_, _05344_, _05332_);
  or (_08523_, _08522_, _08497_);
  or (_08524_, _08523_, _02987_);
  and (_08525_, _08524_, _06246_);
  and (_08526_, _08525_, _08521_);
  or (_08527_, _08526_, _08502_);
  and (_08528_, _08527_, _02986_);
  and (_08529_, _08429_, _05332_);
  or (_08530_, _08529_, _08497_);
  and (_08531_, _08530_, _02866_);
  or (_08532_, _08531_, _05535_);
  or (_08533_, _08532_, _08528_);
  and (_08534_, _08533_, _08496_);
  or (_08535_, _08534_, _02841_);
  and (_08536_, _05461_, _04660_);
  or (_08537_, _08492_, _02842_);
  or (_08538_, _08537_, _08536_);
  and (_08539_, _08538_, _02839_);
  and (_08540_, _08539_, _08535_);
  nor (_08541_, _05740_, _08493_);
  or (_08542_, _08541_, _08492_);
  and (_08543_, _08542_, _02567_);
  or (_08544_, _08543_, _08207_);
  or (_08545_, _08544_, _08540_);
  and (_08546_, _05764_, _04660_);
  or (_08547_, _08492_, _07139_);
  or (_08548_, _08547_, _08546_);
  and (_08549_, _05549_, _04660_);
  or (_08550_, _08549_, _08492_);
  or (_08551_, _08550_, _07140_);
  and (_08552_, _08551_, _07150_);
  and (_08553_, _08552_, _08548_);
  and (_08554_, _08553_, _08545_);
  and (_08555_, _05772_, _04660_);
  or (_08556_, _08555_, _08492_);
  and (_08557_, _08556_, _03148_);
  or (_08558_, _08557_, _08554_);
  and (_08559_, _08558_, _03138_);
  or (_08560_, _08492_, _04740_);
  and (_08561_, _08507_, _03137_);
  and (_08562_, _08550_, _03022_);
  or (_08563_, _08562_, _08561_);
  and (_08564_, _08563_, _08560_);
  or (_08565_, _08564_, _03042_);
  or (_08566_, _08565_, _08559_);
  nor (_08567_, _05763_, _08493_);
  or (_08568_, _08492_, _03043_);
  or (_08569_, _08568_, _08567_);
  and (_08570_, _08569_, _07161_);
  and (_08571_, _08570_, _08566_);
  nor (_08572_, _05771_, _08493_);
  or (_08573_, _08572_, _08492_);
  and (_08574_, _08573_, _03143_);
  or (_08575_, _08574_, _03174_);
  or (_08576_, _08575_, _08571_);
  or (_08577_, _08504_, _03179_);
  and (_08578_, _08577_, _03183_);
  and (_08579_, _08578_, _08576_);
  and (_08580_, _08523_, _02799_);
  or (_08581_, _08580_, _02887_);
  or (_08582_, _08581_, _08579_);
  and (_08583_, _05246_, _04660_);
  or (_08584_, _08492_, _02888_);
  or (_08585_, _08584_, _08583_);
  and (_08586_, _08585_, _34655_);
  and (_08587_, _08586_, _08582_);
  or (_35836_[7], _08587_, _08491_);
  not (_08588_, \oc8051_golden_model_1.P2 [7]);
  nor (_08589_, _34655_, _08588_);
  or (_08590_, _08589_, rst);
  nor (_08591_, _04666_, _08588_);
  not (_08592_, _04666_);
  nor (_08593_, _08592_, _04630_);
  or (_08594_, _08593_, _08591_);
  or (_08595_, _08594_, _02859_);
  nor (_08596_, _05335_, _08588_);
  and (_08597_, _05348_, _05335_);
  or (_08598_, _08597_, _08596_);
  or (_08599_, _08596_, _05502_);
  and (_08600_, _08599_, _02871_);
  and (_08601_, _08600_, _08598_);
  and (_08602_, _05474_, _04666_);
  or (_08603_, _08602_, _08591_);
  or (_08604_, _08603_, _03006_);
  and (_08605_, _04666_, \oc8051_golden_model_1.ACC [7]);
  or (_08606_, _08605_, _08591_);
  and (_08607_, _08606_, _03845_);
  nor (_08608_, _03845_, _08588_);
  or (_08609_, _08608_, _02948_);
  or (_08610_, _08609_, _08607_);
  and (_08611_, _08610_, _02976_);
  and (_08612_, _08611_, _08604_);
  and (_08613_, _08594_, _02946_);
  and (_08614_, _08598_, _02884_);
  or (_08615_, _08614_, _08613_);
  or (_08616_, _08615_, _02880_);
  or (_08617_, _08616_, _08612_);
  or (_08618_, _08606_, _02992_);
  and (_08619_, _08618_, _08617_);
  or (_08620_, _08619_, _02877_);
  and (_08621_, _05344_, _05335_);
  or (_08622_, _08621_, _08596_);
  or (_08623_, _08622_, _02987_);
  and (_08624_, _08623_, _06246_);
  and (_08625_, _08624_, _08620_);
  or (_08626_, _08625_, _08601_);
  and (_08627_, _08626_, _02986_);
  and (_08628_, _08429_, _05335_);
  or (_08629_, _08628_, _08596_);
  and (_08630_, _08629_, _02866_);
  or (_08631_, _08630_, _05535_);
  or (_08632_, _08631_, _08627_);
  and (_08633_, _08632_, _08595_);
  or (_08634_, _08633_, _02841_);
  and (_08635_, _05461_, _04666_);
  or (_08636_, _08591_, _02842_);
  or (_08637_, _08636_, _08635_);
  and (_08638_, _08637_, _02839_);
  and (_08639_, _08638_, _08634_);
  nor (_08640_, _05740_, _08592_);
  or (_08641_, _08640_, _08591_);
  and (_08642_, _08641_, _02567_);
  or (_08643_, _08642_, _08207_);
  or (_08644_, _08643_, _08639_);
  and (_08645_, _05764_, _04666_);
  or (_08646_, _08591_, _07139_);
  or (_08647_, _08646_, _08645_);
  and (_08648_, _05549_, _04666_);
  or (_08649_, _08648_, _08591_);
  or (_08650_, _08649_, _07140_);
  and (_08651_, _08650_, _07150_);
  and (_08652_, _08651_, _08647_);
  and (_08653_, _08652_, _08644_);
  and (_08654_, _05772_, _04666_);
  or (_08655_, _08654_, _08591_);
  and (_08656_, _08655_, _03148_);
  or (_08657_, _08656_, _08653_);
  and (_08658_, _08657_, _03138_);
  or (_08659_, _08591_, _04740_);
  and (_08660_, _08606_, _03137_);
  and (_08661_, _08649_, _03022_);
  or (_08662_, _08661_, _08660_);
  and (_08663_, _08662_, _08659_);
  or (_08664_, _08663_, _03042_);
  or (_08665_, _08664_, _08658_);
  nor (_08666_, _05763_, _08592_);
  or (_08667_, _08591_, _03043_);
  or (_08668_, _08667_, _08666_);
  and (_08669_, _08668_, _07161_);
  and (_08670_, _08669_, _08665_);
  nor (_08671_, _05771_, _08592_);
  or (_08672_, _08671_, _08591_);
  and (_08673_, _08672_, _03143_);
  or (_08674_, _08673_, _03174_);
  or (_08675_, _08674_, _08670_);
  or (_08676_, _08603_, _03179_);
  and (_08677_, _08676_, _03183_);
  and (_08678_, _08677_, _08675_);
  and (_08679_, _08622_, _02799_);
  or (_08680_, _08679_, _02887_);
  or (_08681_, _08680_, _08678_);
  and (_08682_, _05246_, _04666_);
  or (_08683_, _08591_, _02888_);
  or (_08684_, _08683_, _08682_);
  and (_08685_, _08684_, _34655_);
  and (_08686_, _08685_, _08681_);
  or (_35838_[7], _08686_, _08590_);
  not (_08687_, \oc8051_golden_model_1.P3 [7]);
  nor (_08688_, _34655_, _08687_);
  or (_08689_, _08688_, rst);
  nor (_08690_, _04670_, _08687_);
  not (_08691_, _04670_);
  nor (_08692_, _08691_, _04630_);
  or (_08693_, _08692_, _08690_);
  or (_08694_, _08693_, _02859_);
  and (_08695_, _05474_, _04670_);
  or (_08696_, _08695_, _08690_);
  or (_08697_, _08696_, _03006_);
  and (_08698_, _04670_, \oc8051_golden_model_1.ACC [7]);
  or (_08699_, _08698_, _08690_);
  and (_08700_, _08699_, _03845_);
  nor (_08701_, _03845_, _08687_);
  or (_08702_, _08701_, _02948_);
  or (_08703_, _08702_, _08700_);
  and (_08704_, _08703_, _02976_);
  and (_08705_, _08704_, _08697_);
  and (_08706_, _08693_, _02946_);
  nor (_08707_, _05337_, _08687_);
  and (_08708_, _05348_, _05337_);
  or (_08709_, _08708_, _08707_);
  and (_08710_, _08709_, _02884_);
  or (_08711_, _08710_, _08706_);
  or (_08712_, _08711_, _02880_);
  or (_08713_, _08712_, _08705_);
  or (_08714_, _08699_, _02992_);
  and (_08715_, _08714_, _08713_);
  or (_08716_, _08715_, _02877_);
  and (_08717_, _05344_, _05337_);
  or (_08718_, _08717_, _08707_);
  or (_08719_, _08718_, _02987_);
  and (_08720_, _08719_, _06246_);
  and (_08721_, _08720_, _08716_);
  and (_08722_, _05503_, _05337_);
  or (_08723_, _08722_, _08707_);
  and (_08724_, _08723_, _02871_);
  or (_08725_, _08724_, _08721_);
  and (_08726_, _08725_, _02986_);
  and (_08727_, _08429_, _05337_);
  or (_08728_, _08727_, _08707_);
  and (_08729_, _08728_, _02866_);
  or (_08730_, _08729_, _05535_);
  or (_08731_, _08730_, _08726_);
  and (_08732_, _08731_, _08694_);
  or (_08733_, _08732_, _02841_);
  and (_08734_, _05461_, _04670_);
  or (_08735_, _08690_, _02842_);
  or (_08736_, _08735_, _08734_);
  and (_08737_, _08736_, _02839_);
  and (_08738_, _08737_, _08733_);
  nor (_08739_, _05740_, _08691_);
  or (_08740_, _08739_, _08690_);
  and (_08741_, _08740_, _02567_);
  or (_08742_, _08741_, _08207_);
  or (_08743_, _08742_, _08738_);
  and (_08744_, _05764_, _04670_);
  or (_08745_, _08690_, _07139_);
  or (_08746_, _08745_, _08744_);
  and (_08747_, _05549_, _04670_);
  or (_08748_, _08747_, _08690_);
  or (_08749_, _08748_, _07140_);
  and (_08750_, _08749_, _07150_);
  and (_08751_, _08750_, _08746_);
  and (_08752_, _08751_, _08743_);
  and (_08753_, _05772_, _04670_);
  or (_08754_, _08753_, _08690_);
  and (_08755_, _08754_, _03148_);
  or (_08756_, _08755_, _08752_);
  and (_08757_, _08756_, _03138_);
  or (_08758_, _08690_, _04740_);
  and (_08759_, _08699_, _03137_);
  and (_08760_, _08748_, _03022_);
  or (_08761_, _08760_, _08759_);
  and (_08762_, _08761_, _08758_);
  or (_08763_, _08762_, _03042_);
  or (_08764_, _08763_, _08757_);
  nor (_08765_, _05763_, _08691_);
  or (_08766_, _08690_, _03043_);
  or (_08767_, _08766_, _08765_);
  and (_08768_, _08767_, _07161_);
  and (_08769_, _08768_, _08764_);
  nor (_08770_, _05771_, _08691_);
  or (_08771_, _08770_, _08690_);
  and (_08772_, _08771_, _03143_);
  or (_08773_, _08772_, _03174_);
  or (_08774_, _08773_, _08769_);
  or (_08775_, _08696_, _03179_);
  and (_08776_, _08775_, _03183_);
  and (_08777_, _08776_, _08774_);
  and (_08778_, _08718_, _02799_);
  or (_08779_, _08778_, _02887_);
  or (_08780_, _08779_, _08777_);
  and (_08781_, _05246_, _04670_);
  or (_08782_, _08690_, _02888_);
  or (_08783_, _08782_, _08781_);
  and (_08784_, _08783_, _34655_);
  and (_08785_, _08784_, _08780_);
  or (_35840_[7], _08785_, _08689_);
  and (_08786_, _02798_, _02498_);
  not (_08787_, _08786_);
  not (_08788_, _02510_);
  not (_08789_, _08112_);
  not (_08790_, _02234_);
  and (_08791_, _05265_, _08790_);
  and (_08792_, _08791_, \oc8051_golden_model_1.PC [7]);
  and (_08793_, _08792_, \oc8051_golden_model_1.PC [8]);
  and (_08794_, _08793_, \oc8051_golden_model_1.PC [9]);
  and (_08795_, _08794_, \oc8051_golden_model_1.PC [10]);
  and (_08796_, _08795_, \oc8051_golden_model_1.PC [11]);
  and (_08797_, _08796_, \oc8051_golden_model_1.PC [12]);
  and (_08798_, _08797_, \oc8051_golden_model_1.PC [13]);
  and (_08799_, _08798_, \oc8051_golden_model_1.PC [14]);
  nor (_08800_, _08799_, \oc8051_golden_model_1.PC [15]);
  and (_08801_, _08799_, \oc8051_golden_model_1.PC [15]);
  nor (_08802_, _08801_, _08800_);
  and (_08803_, _08031_, _07189_);
  nor (_08804_, _08803_, _08802_);
  and (_08806_, _07936_, _07234_);
  nor (_08807_, _08806_, _08802_);
  and (_08808_, _02798_, _02532_);
  nor (_08809_, _03143_, _02533_);
  nor (_08810_, _08809_, _06206_);
  or (_08811_, _08810_, _08808_);
  nor (_08812_, _07921_, _03141_);
  not (_08813_, _07915_);
  nor (_08814_, _07908_, _07309_);
  and (_08815_, _08814_, _08813_);
  nor (_08817_, _08815_, _08802_);
  and (_08818_, _02798_, _02529_);
  nor (_08819_, _03137_, _02530_);
  nor (_08820_, _08819_, _06206_);
  or (_08821_, _08820_, _08818_);
  nor (_08822_, _07860_, _03146_);
  and (_08823_, _07850_, _07845_);
  nor (_08824_, _08823_, _08802_);
  nor (_08825_, _06191_, \oc8051_golden_model_1.PC [14]);
  nor (_08826_, _08825_, _06192_);
  not (_08828_, _08826_);
  nor (_08829_, _08828_, _05302_);
  and (_08830_, _08828_, _05302_);
  nor (_08831_, _08830_, _08829_);
  not (_08832_, _08831_);
  nor (_08833_, _06190_, \oc8051_golden_model_1.PC [13]);
  nor (_08834_, _08833_, _06191_);
  not (_08835_, _08834_);
  nor (_08836_, _08835_, _05302_);
  and (_08837_, _08835_, _05302_);
  nor (_08839_, _06189_, \oc8051_golden_model_1.PC [12]);
  nor (_08840_, _08839_, _06190_);
  not (_08841_, _08840_);
  nor (_08842_, _08841_, _05302_);
  nor (_08843_, _06188_, \oc8051_golden_model_1.PC [11]);
  nor (_08844_, _08843_, _06189_);
  not (_08845_, _08844_);
  nor (_08846_, _08845_, _05302_);
  and (_08847_, _08845_, _05302_);
  nor (_08848_, _08847_, _08846_);
  nor (_08850_, _06187_, \oc8051_golden_model_1.PC [10]);
  nor (_08851_, _08850_, _06188_);
  not (_08852_, _08851_);
  nor (_08853_, _08852_, _05302_);
  and (_08854_, _08852_, _05302_);
  nor (_08855_, _08854_, _08853_);
  and (_08856_, _08855_, _08848_);
  nor (_08857_, _06186_, \oc8051_golden_model_1.PC [9]);
  nor (_08858_, _08857_, _06187_);
  not (_08859_, _08858_);
  nor (_08861_, _08859_, _05302_);
  and (_08862_, _08859_, _05302_);
  nor (_08863_, _08862_, _08861_);
  nor (_08864_, _06147_, _05302_);
  and (_08865_, _06147_, _05302_);
  and (_08866_, _06142_, _05264_);
  nor (_08867_, _08866_, \oc8051_golden_model_1.PC [6]);
  nor (_08868_, _08867_, _06143_);
  not (_08869_, _08868_);
  nor (_08870_, _08869_, _05585_);
  and (_08872_, _08869_, _05585_);
  nor (_08873_, _08872_, _08870_);
  not (_08874_, _08873_);
  and (_08875_, _06142_, \oc8051_golden_model_1.PC [4]);
  nor (_08876_, _08875_, \oc8051_golden_model_1.PC [5]);
  nor (_08877_, _08876_, _08866_);
  not (_08878_, _08877_);
  nor (_08879_, _08878_, _05649_);
  and (_08880_, _08878_, _05649_);
  nor (_08881_, _06142_, \oc8051_golden_model_1.PC [4]);
  nor (_08882_, _08881_, _08875_);
  not (_08883_, _08882_);
  nor (_08884_, _08883_, _05617_);
  nor (_08885_, _06141_, \oc8051_golden_model_1.PC [3]);
  nor (_08886_, _08885_, _06142_);
  not (_08887_, _08886_);
  nor (_08888_, _08887_, _03128_);
  and (_08889_, _08887_, _03128_);
  nor (_08890_, _02251_, \oc8051_golden_model_1.PC [2]);
  nor (_08891_, _08890_, _06141_);
  not (_08892_, _08891_);
  nor (_08893_, _08892_, _03262_);
  not (_08894_, _02544_);
  nor (_08895_, _03720_, _08894_);
  nor (_08896_, _03505_, \oc8051_golden_model_1.PC [0]);
  and (_08897_, _03720_, _08894_);
  nor (_08898_, _08897_, _08895_);
  and (_08899_, _08898_, _08896_);
  nor (_08900_, _08899_, _08895_);
  and (_08901_, _08892_, _03262_);
  nor (_08902_, _08901_, _08893_);
  not (_08903_, _08902_);
  nor (_08904_, _08903_, _08900_);
  nor (_08905_, _08904_, _08893_);
  nor (_08906_, _08905_, _08889_);
  nor (_08907_, _08906_, _08888_);
  and (_08908_, _08883_, _05617_);
  nor (_08909_, _08908_, _08884_);
  not (_08910_, _08909_);
  nor (_08911_, _08910_, _08907_);
  nor (_08912_, _08911_, _08884_);
  nor (_08913_, _08912_, _08880_);
  nor (_08914_, _08913_, _08879_);
  nor (_08915_, _08914_, _08874_);
  nor (_08916_, _08915_, _08870_);
  nor (_08917_, _08916_, _08865_);
  or (_08918_, _08917_, _08864_);
  nor (_08919_, _06144_, \oc8051_golden_model_1.PC [8]);
  nor (_08920_, _08919_, _06186_);
  not (_08921_, _08920_);
  nor (_08922_, _08921_, _05302_);
  and (_08923_, _08921_, _05302_);
  nor (_08924_, _08923_, _08922_);
  and (_08925_, _08924_, _08918_);
  and (_08926_, _08925_, _08863_);
  and (_08927_, _08926_, _08856_);
  nor (_08928_, _08922_, _08861_);
  not (_08929_, _08928_);
  and (_08930_, _08929_, _08856_);
  or (_08931_, _08930_, _08853_);
  or (_08932_, _08931_, _08927_);
  nor (_08933_, _08932_, _08846_);
  not (_08934_, _08933_);
  and (_08935_, _08841_, _05302_);
  nor (_08936_, _08935_, _08842_);
  and (_08937_, _08936_, _08934_);
  nor (_08938_, _08937_, _08842_);
  nor (_08939_, _08938_, _08837_);
  nor (_08940_, _08939_, _08836_);
  nor (_08941_, _08940_, _08832_);
  nor (_08942_, _08941_, _08829_);
  not (_08943_, _06195_);
  and (_08944_, _08943_, _05302_);
  nor (_08945_, _08943_, _05302_);
  nor (_08946_, _08945_, _08944_);
  and (_08947_, _08946_, _08942_);
  nor (_08948_, _08946_, _08942_);
  nor (_08949_, _08948_, _08947_);
  not (_08950_, _05514_);
  or (_08951_, _05461_, _02763_);
  and (_08952_, _08951_, _08950_);
  or (_08953_, _06162_, _02924_);
  or (_08954_, _05855_, _04374_);
  and (_08955_, _08954_, _08953_);
  and (_08956_, _08955_, _08952_);
  or (_08957_, _06083_, _04663_);
  or (_08958_, _06170_, _03220_);
  and (_08959_, _08958_, _08957_);
  or (_08960_, _06128_, _04657_);
  or (_08961_, _06171_, _03647_);
  and (_08962_, _08961_, _08960_);
  and (_08963_, _08962_, _08959_);
  and (_08964_, _08963_, _08956_);
  or (_08965_, _06166_, _04353_);
  and (_08966_, _06166_, _04353_);
  not (_08967_, _08966_);
  and (_08968_, _08967_, _08965_);
  or (_08969_, _06167_, _03356_);
  or (_08970_, _06036_, _04385_);
  and (_08971_, _08970_, _08969_);
  and (_08972_, _08971_, _08968_);
  or (_08973_, _05945_, _02833_);
  or (_08974_, _06163_, _03687_);
  or (_08975_, _05900_, _03951_);
  and (_08976_, _08975_, _08974_);
  and (_08977_, _08976_, _08973_);
  nand (_08978_, _08977_, _08972_);
  and (_08979_, _05945_, _02833_);
  nor (_08980_, _08979_, _08978_);
  nand (_08981_, _08980_, _08964_);
  and (_08982_, _08981_, _08949_);
  nor (_08983_, _08981_, _06195_);
  nor (_08984_, _08983_, _08982_);
  and (_08985_, _02840_, _02870_);
  not (_08986_, _08985_);
  nor (_08987_, _08986_, _08984_);
  not (_08988_, _06206_);
  not (_08989_, _02595_);
  nor (_08990_, _02877_, _08989_);
  and (_08991_, _08990_, _03962_);
  nor (_08992_, _08991_, _08988_);
  nor (_08993_, _02884_, _04225_);
  and (_08994_, _08993_, _07474_);
  nor (_08995_, _08994_, _06206_);
  nor (_08996_, _02596_, _02540_);
  nor (_08997_, _08996_, _07405_);
  not (_08998_, _08997_);
  and (_08999_, _05085_, _05037_);
  and (_09000_, _05468_, _08999_);
  and (_09001_, _04837_, _04739_);
  and (_09002_, _09001_, _05465_);
  and (_09003_, _09002_, _09000_);
  and (_09004_, _09003_, _08943_);
  not (_09005_, _08949_);
  nor (_09006_, _09003_, _09005_);
  or (_09007_, _09006_, _03006_);
  or (_09008_, _09007_, _09004_);
  and (_09009_, _05353_, _05351_);
  and (_09010_, _04020_, _03838_);
  and (_09011_, _09010_, _05259_);
  and (_09012_, _09011_, _09009_);
  and (_09013_, _09012_, _06206_);
  nor (_09014_, _06202_, \oc8051_golden_model_1.PC [14]);
  nor (_09015_, _09014_, _06203_);
  not (_09016_, _09015_);
  nor (_09017_, _09016_, _02763_);
  and (_09018_, _09016_, _02763_);
  nor (_09019_, _09018_, _09017_);
  nor (_09020_, _06201_, \oc8051_golden_model_1.PC [13]);
  nor (_09021_, _09020_, _06202_);
  not (_09022_, _09021_);
  nor (_09023_, _09022_, _02763_);
  and (_09024_, _09022_, _02763_);
  nor (_09025_, _06200_, \oc8051_golden_model_1.PC [12]);
  nor (_09026_, _09025_, _06201_);
  not (_09027_, _09026_);
  nor (_09028_, _09027_, _02763_);
  nor (_09029_, _06199_, \oc8051_golden_model_1.PC [11]);
  nor (_09030_, _09029_, _06200_);
  not (_09031_, _09030_);
  nor (_09032_, _09031_, _02763_);
  and (_09033_, _09031_, _02763_);
  nor (_09034_, _09033_, _09032_);
  nor (_09035_, _06198_, \oc8051_golden_model_1.PC [10]);
  nor (_09036_, _09035_, _06199_);
  not (_09037_, _09036_);
  nor (_09038_, _09037_, _02763_);
  and (_09039_, _09037_, _02763_);
  nor (_09040_, _09039_, _09038_);
  and (_09041_, _09040_, _09034_);
  nor (_09042_, _06197_, \oc8051_golden_model_1.PC [9]);
  nor (_09043_, _09042_, _06198_);
  not (_09044_, _09043_);
  nor (_09045_, _09044_, _02763_);
  and (_09046_, _09044_, _02763_);
  nor (_09047_, _09046_, _09045_);
  nor (_09048_, _05507_, _02763_);
  and (_09049_, _05507_, _02763_);
  nor (_09050_, _09049_, _09048_);
  not (_09051_, _09050_);
  and (_09052_, _05264_, _02638_);
  nor (_09053_, _09052_, \oc8051_golden_model_1.PC [6]);
  nor (_09054_, _09053_, _05266_);
  not (_09055_, _09054_);
  nor (_09056_, _09055_, _02924_);
  and (_09057_, _09055_, _02924_);
  nor (_09058_, _09057_, _09056_);
  and (_09059_, _02638_, \oc8051_golden_model_1.PC [4]);
  nor (_09060_, _09059_, \oc8051_golden_model_1.PC [5]);
  nor (_09061_, _09060_, _09052_);
  not (_09062_, _09061_);
  nor (_09063_, _09062_, _03220_);
  and (_09064_, _09062_, _03220_);
  nor (_09065_, _02638_, \oc8051_golden_model_1.PC [4]);
  nor (_09066_, _09065_, _09059_);
  not (_09067_, _09066_);
  nor (_09068_, _09067_, _03647_);
  and (_09069_, _02794_, _02640_);
  nor (_09070_, _02794_, _02640_);
  nor (_09071_, _03356_, _02620_);
  nor (_09072_, _03687_, \oc8051_golden_model_1.PC [1]);
  and (_09073_, _02833_, \oc8051_golden_model_1.PC [0]);
  and (_09074_, _03687_, \oc8051_golden_model_1.PC [1]);
  nor (_09075_, _09074_, _09072_);
  and (_09076_, _09075_, _09073_);
  nor (_09077_, _09076_, _09072_);
  and (_09078_, _03356_, _02620_);
  nor (_09079_, _09078_, _09071_);
  not (_09080_, _09079_);
  nor (_09081_, _09080_, _09077_);
  nor (_09082_, _09081_, _09071_);
  nor (_09083_, _09082_, _09070_);
  nor (_09084_, _09083_, _09069_);
  not (_09085_, _09084_);
  and (_09086_, _09067_, _03647_);
  nor (_09087_, _09086_, _09068_);
  and (_09088_, _09087_, _09085_);
  nor (_09089_, _09088_, _09068_);
  nor (_09090_, _09089_, _09064_);
  or (_09091_, _09090_, _09063_);
  and (_09092_, _09091_, _09058_);
  nor (_09093_, _09092_, _09056_);
  nor (_09094_, _09093_, _09051_);
  nor (_09095_, _09094_, _09048_);
  nor (_09096_, _05267_, \oc8051_golden_model_1.PC [8]);
  nor (_09097_, _09096_, _06197_);
  not (_09098_, _09097_);
  nor (_09099_, _09098_, _02763_);
  and (_09100_, _09098_, _02763_);
  nor (_09101_, _09100_, _09099_);
  not (_09102_, _09101_);
  nor (_09103_, _09102_, _09095_);
  and (_09104_, _09103_, _09047_);
  and (_09105_, _09104_, _09041_);
  nor (_09106_, _09099_, _09045_);
  not (_09107_, _09106_);
  and (_09108_, _09107_, _09041_);
  or (_09109_, _09108_, _09038_);
  or (_09110_, _09109_, _09105_);
  nor (_09111_, _09110_, _09032_);
  not (_09112_, _09111_);
  and (_09113_, _09027_, _02763_);
  nor (_09114_, _09113_, _09028_);
  and (_09115_, _09114_, _09112_);
  nor (_09116_, _09115_, _09028_);
  nor (_09117_, _09116_, _09024_);
  nor (_09118_, _09117_, _09023_);
  not (_09119_, _09118_);
  and (_09120_, _09119_, _09019_);
  nor (_09121_, _09120_, _09017_);
  and (_09122_, _08988_, _02763_);
  nor (_09123_, _08988_, _02763_);
  nor (_09124_, _09123_, _09122_);
  and (_09125_, _09124_, _09121_);
  nor (_09126_, _09124_, _09121_);
  nor (_09127_, _09126_, _09125_);
  nor (_09128_, _09012_, _09127_);
  or (_09129_, _09128_, _05361_);
  nor (_09130_, _09129_, _09013_);
  and (_09131_, _08802_, _07433_);
  not (_09132_, _05361_);
  not (_09133_, _07433_);
  and (_09134_, _07439_, _03382_);
  nor (_09135_, _09134_, _07423_);
  and (_09136_, _06206_, _03845_);
  nor (_09137_, _02840_, _02304_);
  nor (_09138_, _09137_, _02602_);
  nand (_09139_, _04194_, \oc8051_golden_model_1.PC [15]);
  nor (_09140_, _09139_, _09138_);
  or (_09141_, _09140_, _09136_);
  and (_09142_, _09141_, _09135_);
  not (_09143_, _08802_);
  not (_09144_, _09138_);
  and (_09145_, _09144_, _09135_);
  nor (_09146_, _09145_, _09143_);
  or (_09147_, _09146_, _09142_);
  and (_09148_, _09147_, _02603_);
  nor (_09149_, _07410_, _07414_);
  and (_09150_, _02798_, _03382_);
  nor (_09151_, _09150_, _03724_);
  and (_09152_, _09151_, _09149_);
  and (_09153_, _09152_, _07419_);
  not (_09154_, _09153_);
  and (_09155_, _06206_, _03849_);
  or (_09156_, _09155_, _09154_);
  nor (_09157_, _09156_, _09148_);
  nor (_09158_, _09153_, _08802_);
  nor (_09159_, _09158_, _02951_);
  not (_09160_, _09159_);
  nor (_09161_, _09160_, _09157_);
  and (_09162_, _06206_, _02951_);
  nor (_09163_, _09162_, _07436_);
  not (_09164_, _09163_);
  nor (_09165_, _09164_, _09161_);
  and (_09166_, _09143_, _07436_);
  nor (_09167_, _09166_, _09165_);
  and (_09168_, _09167_, _02601_);
  not (_09169_, _02601_);
  and (_09170_, _06206_, _09169_);
  or (_09171_, _09170_, _09168_);
  and (_09172_, _09171_, _09133_);
  or (_09173_, _09172_, _09132_);
  nor (_09174_, _09173_, _09131_);
  not (_09175_, _09174_);
  nor (_09176_, _03840_, _02948_);
  nand (_09177_, _09176_, _09175_);
  or (_09178_, _09177_, _09130_);
  and (_09179_, _09178_, _09008_);
  or (_09180_, _09179_, _08998_);
  nand (_09181_, _08997_, _05371_);
  nand (_09182_, _09181_, _08802_);
  and (_09183_, _09182_, _08994_);
  and (_09184_, _09183_, _09180_);
  nor (_09185_, _09184_, _08995_);
  and (_09186_, _07402_, _07481_);
  not (_09187_, _09186_);
  nor (_09188_, _09187_, _09185_);
  nor (_09189_, _09186_, _08802_);
  nor (_09190_, _09189_, _02880_);
  not (_09191_, _09190_);
  nor (_09192_, _09191_, _09188_);
  nor (_09193_, _07434_, _02594_);
  or (_09194_, _09193_, _02880_);
  not (_09195_, _09194_);
  nor (_09196_, _09193_, _06206_);
  nor (_09197_, _09196_, _09195_);
  nor (_09198_, _09197_, _09192_);
  not (_09199_, _08991_);
  not (_09200_, _09193_);
  nor (_09201_, _09200_, _08802_);
  nor (_09202_, _09201_, _09199_);
  not (_09203_, _09202_);
  nor (_09204_, _09203_, _09198_);
  nor (_09205_, _09204_, _08992_);
  nor (_09206_, _07231_, _03298_);
  nor (_09207_, _09206_, _02590_);
  not (_09208_, _09207_);
  and (_09209_, _09208_, _03005_);
  not (_09210_, _09209_);
  or (_09211_, _09210_, _09205_);
  not (_09212_, _04631_);
  and (_09213_, _04630_, _02838_);
  nor (_09214_, _09213_, _09212_);
  nor (_09215_, _04790_, _04374_);
  and (_09216_, _04790_, _04374_);
  nor (_09217_, _09216_, _09215_);
  and (_09218_, _09217_, _09214_);
  nor (_09219_, _04894_, _04663_);
  and (_09220_, _04894_, _04663_);
  nor (_09221_, _09220_, _09219_);
  and (_09222_, _05192_, _04657_);
  nor (_09223_, _05192_, _04657_);
  nor (_09224_, _09223_, _09222_);
  and (_09225_, _09224_, _09221_);
  and (_09226_, _09225_, _09218_);
  and (_09227_, _04275_, _02794_);
  and (_09228_, _04449_, _04385_);
  nor (_09229_, _09228_, _09227_);
  nor (_09230_, _04275_, _02794_);
  nor (_09231_, _04449_, _04385_);
  nor (_09232_, _09231_, _09230_);
  and (_09233_, _09232_, _09229_);
  nor (_09234_, _04020_, _03951_);
  and (_09235_, _04020_, _03951_);
  nor (_09236_, _09235_, _09234_);
  and (_09237_, _03838_, _02837_);
  and (_09238_, _03872_, _02833_);
  nor (_09239_, _09238_, _09237_);
  and (_09240_, _09239_, _09236_);
  and (_09241_, _09240_, _09233_);
  and (_09242_, _09241_, _09226_);
  and (_09243_, _09242_, _08943_);
  nor (_09244_, _09242_, _09005_);
  or (_09245_, _09244_, _09209_);
  or (_09246_, _09245_, _09243_);
  and (_09247_, _09246_, _08986_);
  and (_09248_, _09247_, _09211_);
  nor (_09249_, _02590_, _02540_);
  not (_09250_, _09249_);
  and (_09251_, _09250_, _03030_);
  not (_09252_, _09251_);
  or (_09253_, _09252_, _09248_);
  nor (_09254_, _09253_, _08987_);
  and (_09255_, _09249_, _08802_);
  not (_09256_, _09255_);
  not (_09257_, _02591_);
  nor (_09258_, _02871_, _09257_);
  and (_09259_, _05379_, _02965_);
  nor (_09260_, _02969_, _02937_);
  and (_09261_, _09260_, _04063_);
  and (_09262_, _09261_, _09259_);
  and (_09263_, _09262_, _09258_);
  and (_09264_, _09263_, _09256_);
  nor (_09265_, _08122_, _08121_);
  nor (_09266_, _09265_, _08125_);
  nor (_09267_, _08120_, _07867_);
  and (_09268_, _09267_, _09266_);
  nor (_09269_, _08126_, _08127_);
  nor (_09270_, _09269_, _08130_);
  and (_09271_, _02837_, _02696_);
  nor (_09272_, _09271_, _08132_);
  not (_09273_, _07783_);
  nor (_09274_, _09273_, _09272_);
  and (_09275_, _09274_, _09270_);
  and (_09276_, _09275_, _09268_);
  not (_09277_, _09276_);
  and (_09278_, _09277_, _08949_);
  not (_09279_, _03029_);
  and (_09280_, _09276_, _08943_);
  nor (_09281_, _09280_, _09279_);
  not (_09282_, _09281_);
  nor (_09283_, _09282_, _09278_);
  nor (_09284_, _07566_, \oc8051_golden_model_1.ACC [3]);
  and (_09285_, _07566_, \oc8051_golden_model_1.ACC [3]);
  nor (_09286_, _09285_, _09284_);
  and (_09287_, _09286_, _08090_);
  nor (_09288_, _07607_, \oc8051_golden_model_1.ACC [0]);
  and (_09289_, _07607_, \oc8051_golden_model_1.ACC [0]);
  nor (_09290_, _09289_, _09288_);
  and (_09291_, _09290_, _07700_);
  and (_09292_, _09291_, _09287_);
  and (_09293_, _08081_, _08085_);
  not (_09294_, _08073_);
  and (_09295_, _08077_, _09294_);
  and (_09296_, _09295_, _09293_);
  and (_09297_, _09296_, _09292_);
  and (_09298_, _09297_, _08943_);
  not (_09299_, _02954_);
  nor (_09300_, _09297_, _09005_);
  or (_09301_, _09300_, _09299_);
  nor (_09302_, _09301_, _09298_);
  nor (_09303_, _09302_, _09283_);
  and (_09304_, _09303_, _09264_);
  not (_09305_, _09304_);
  nor (_09306_, _09305_, _09254_);
  and (_09307_, _02939_, _02566_);
  nor (_09308_, _09307_, _06252_);
  and (_09309_, _09308_, _08227_);
  not (_09310_, _09309_);
  nor (_09311_, _09263_, _06206_);
  nor (_09312_, _09311_, _09310_);
  not (_09313_, _09312_);
  nor (_09314_, _09313_, _09306_);
  and (_09315_, _09310_, _08802_);
  and (_09316_, _02942_, _02589_);
  not (_09317_, _09316_);
  or (_09318_, _09317_, _09315_);
  or (_09319_, _09318_, _09314_);
  nor (_09320_, _07400_, _07397_);
  or (_09321_, _09316_, _06206_);
  and (_09322_, _09321_, _09320_);
  and (_09323_, _09322_, _09319_);
  nor (_09324_, _07540_, _02979_);
  not (_09325_, _09324_);
  not (_09326_, _09320_);
  and (_09327_, _09326_, _08802_);
  nor (_09328_, _09327_, _09325_);
  not (_09329_, _09328_);
  nor (_09330_, _09329_, _09323_);
  nor (_09331_, _09324_, _06206_);
  nor (_09332_, _09331_, _07721_);
  not (_09333_, _09332_);
  nor (_09334_, _09333_, _09330_);
  nor (_09335_, _02866_, _02569_);
  and (_09336_, _09335_, _02571_);
  not (_09337_, _09335_);
  nor (_09338_, _09337_, _08802_);
  nor (_09339_, _09338_, _09336_);
  nor (_09340_, _09339_, _09334_);
  nor (_09341_, _09335_, _06206_);
  nor (_09342_, _09341_, _03046_);
  not (_09343_, _09342_);
  or (_09344_, _09343_, _09340_);
  and (_09345_, _02860_, _08211_);
  and (_09346_, _08943_, _02860_);
  or (_09347_, _09346_, _09345_);
  nand (_09348_, _09347_, _09344_);
  nor (_09349_, _06206_, _02860_);
  nor (_09350_, _09349_, _02567_);
  and (_09351_, _09350_, _09348_);
  or (_09352_, _06786_, _02542_);
  nor (_09353_, _09352_, _02567_);
  nor (_09354_, _09352_, _06195_);
  nor (_09355_, _09354_, _09353_);
  nor (_09356_, _09355_, _09351_);
  not (_09357_, _09352_);
  nor (_09358_, _09357_, _08802_);
  or (_09359_, _09358_, _09356_);
  nor (_09360_, _02930_, _02516_);
  and (_09361_, _09360_, _09359_);
  and (_09362_, _02798_, _02515_);
  nor (_09363_, _09360_, _06206_);
  or (_09364_, _09363_, _09362_);
  or (_09365_, _09364_, _09361_);
  not (_09366_, _09362_);
  nor (_09367_, _09366_, _09127_);
  nor (_09368_, _09367_, _05749_);
  nand (_09369_, _09368_, _09365_);
  nor (_09370_, _06206_, _05748_);
  nor (_09371_, _09370_, _02834_);
  nand (_09372_, _09371_, _09369_);
  and (_09373_, _06195_, _02834_);
  nor (_09374_, _09373_, _07830_);
  nand (_09375_, _09374_, _09372_);
  and (_09376_, _02541_, _02521_);
  nor (_09377_, _07831_, _06206_);
  nor (_09378_, _09377_, _09376_);
  nand (_09379_, _09378_, _09375_);
  not (_09380_, \oc8051_golden_model_1.DPH [0]);
  and (_09381_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_09382_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_09383_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09384_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09385_, _09384_, _09383_);
  not (_09386_, _09385_);
  and (_09387_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_09388_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_09389_, _09388_, _09387_);
  not (_09390_, _09389_);
  and (_09391_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09392_, _02649_, _02645_);
  nor (_09393_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09394_, _09393_, _09391_);
  not (_09395_, _09394_);
  nor (_09396_, _09395_, _09392_);
  nor (_09397_, _09396_, _09391_);
  nor (_09398_, _09397_, _09390_);
  nor (_09399_, _09398_, _09387_);
  nor (_09400_, _09399_, _09386_);
  nor (_09401_, _09400_, _09383_);
  nor (_09402_, _09401_, _09382_);
  nor (_09403_, _09402_, _09381_);
  nor (_09404_, _09403_, _09380_);
  and (_09405_, _09404_, \oc8051_golden_model_1.DPH [1]);
  and (_09406_, _09405_, \oc8051_golden_model_1.DPH [2]);
  and (_09407_, _09406_, \oc8051_golden_model_1.DPH [3]);
  and (_09408_, _09407_, \oc8051_golden_model_1.DPH [4]);
  and (_09409_, _09408_, \oc8051_golden_model_1.DPH [5]);
  and (_09410_, _09409_, \oc8051_golden_model_1.DPH [6]);
  nor (_09411_, _09410_, \oc8051_golden_model_1.DPH [7]);
  and (_09412_, _09410_, \oc8051_golden_model_1.DPH [7]);
  nor (_09413_, _09412_, _09411_);
  and (_09414_, _09413_, _09376_);
  nor (_09415_, _02928_, _02522_);
  not (_09416_, _09415_);
  nor (_09417_, _09416_, _09414_);
  nand (_09418_, _09417_, _09379_);
  and (_09419_, _02798_, _02521_);
  nor (_09420_, _09415_, _06206_);
  nor (_09421_, _09420_, _09419_);
  nand (_09423_, _09421_, _09418_);
  and (_09424_, _08166_, _06206_);
  nor (_09425_, _09127_, _08166_);
  or (_09426_, _09425_, _09424_);
  and (_09427_, _09426_, _09419_);
  not (_09428_, _08823_);
  nor (_09429_, _09428_, _09427_);
  and (_09430_, _09429_, _09423_);
  or (_09431_, _09430_, _08824_);
  nand (_09432_, _09431_, _08822_);
  nor (_09433_, _08822_, _06206_);
  nor (_09434_, _09433_, _03051_);
  nand (_09435_, _09434_, _09432_);
  and (_09436_, _06195_, _03051_);
  nor (_09437_, _03148_, _02524_);
  not (_09438_, _09437_);
  nor (_09439_, _09438_, _09436_);
  nand (_09440_, _09439_, _09435_);
  and (_09441_, _02798_, _02523_);
  nor (_09442_, _09437_, _06206_);
  nor (_09444_, _09442_, _09441_);
  nand (_09445_, _09444_, _09440_);
  not (_09446_, _09441_);
  not (_09447_, _08166_);
  nand (_09448_, _09447_, _06206_);
  or (_09449_, _09127_, _09447_);
  and (_09450_, _09449_, _09448_);
  or (_09451_, _09450_, _09446_);
  nand (_09452_, _09451_, _09445_);
  and (_09453_, _07891_, _07882_);
  nand (_09454_, _09453_, _09452_);
  nor (_09455_, _07311_, _03135_);
  not (_09456_, _09455_);
  nor (_09457_, _09453_, _09143_);
  nor (_09458_, _09457_, _09456_);
  nand (_09459_, _09458_, _09454_);
  nor (_09460_, _09455_, _06206_);
  nor (_09461_, _09460_, _03022_);
  nand (_09462_, _09461_, _09459_);
  not (_09463_, _08819_);
  and (_09464_, _06195_, _03022_);
  nor (_09465_, _09464_, _09463_);
  and (_09466_, _09465_, _09462_);
  or (_09467_, _09466_, _08821_);
  not (_09468_, _08815_);
  and (_09469_, _09127_, _07288_);
  not (_09470_, _08818_);
  nor (_09471_, _06206_, _07288_);
  nor (_09472_, _09471_, _09470_);
  not (_09473_, _09472_);
  nor (_09474_, _09473_, _09469_);
  nor (_09475_, _09474_, _09468_);
  and (_09476_, _09475_, _09467_);
  or (_09477_, _09476_, _08817_);
  nand (_09478_, _09477_, _08812_);
  nor (_09479_, _08812_, _06206_);
  nor (_09480_, _09479_, _03042_);
  nand (_09481_, _09480_, _09478_);
  not (_09482_, _08809_);
  and (_09483_, _06195_, _03042_);
  nor (_09484_, _09483_, _09482_);
  and (_09485_, _09484_, _09481_);
  or (_09486_, _09485_, _08811_);
  not (_09487_, _08806_);
  nand (_09488_, _09127_, \oc8051_golden_model_1.PSW [7]);
  or (_09489_, _06206_, \oc8051_golden_model_1.PSW [7]);
  and (_09490_, _09489_, _08808_);
  and (_09491_, _09490_, _09488_);
  nor (_09492_, _09491_, _09487_);
  and (_09493_, _09492_, _09486_);
  or (_09494_, _09493_, _08807_);
  nand (_09495_, _09494_, _07965_);
  nor (_09496_, _07965_, _06206_);
  nor (_09497_, _09496_, _07995_);
  and (_09498_, _09497_, _09495_);
  and (_09499_, _08802_, _07995_);
  or (_09500_, _09499_, _03155_);
  nor (_09501_, _09500_, _09498_);
  and (_09502_, _04630_, _03155_);
  or (_09503_, _09502_, _09501_);
  nand (_09504_, _09503_, _05790_);
  nor (_09505_, _06206_, _05790_);
  nor (_09506_, _09505_, _03040_);
  nand (_09507_, _09506_, _09504_);
  not (_09508_, _04642_);
  and (_09509_, _05316_, \oc8051_golden_model_1.PSW [2]);
  and (_09510_, _05313_, \oc8051_golden_model_1.ACC [2]);
  nor (_09511_, _09510_, _09509_);
  and (_09512_, _05319_, \oc8051_golden_model_1.IP [2]);
  and (_09513_, _05321_, \oc8051_golden_model_1.B [2]);
  nor (_09514_, _09513_, _09512_);
  and (_09515_, _09514_, _09511_);
  and (_09516_, _05337_, \oc8051_golden_model_1.P3INREG [2]);
  not (_09517_, _09516_);
  and (_09518_, _04635_, \oc8051_golden_model_1.P0INREG [2]);
  and (_09519_, _05335_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_09520_, _09519_, _09518_);
  and (_09521_, _09520_, _09517_);
  and (_09522_, _05326_, \oc8051_golden_model_1.SCON [2]);
  and (_09523_, _05328_, \oc8051_golden_model_1.IE [2]);
  nor (_09524_, _09523_, _09522_);
  and (_09525_, _05310_, \oc8051_golden_model_1.TCON [2]);
  and (_09526_, _05332_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_09527_, _09526_, _09525_);
  and (_09528_, _09527_, _09524_);
  and (_09529_, _09528_, _09521_);
  and (_09530_, _09529_, _09515_);
  and (_09531_, _09530_, _05087_);
  nor (_09532_, _09531_, _09508_);
  not (_09533_, _04637_);
  and (_09534_, _05310_, \oc8051_golden_model_1.TCON [1]);
  and (_09535_, _05321_, \oc8051_golden_model_1.B [1]);
  nor (_09536_, _09535_, _09534_);
  and (_09537_, _05316_, \oc8051_golden_model_1.PSW [1]);
  not (_09538_, _09537_);
  and (_09539_, _05319_, \oc8051_golden_model_1.IP [1]);
  and (_09540_, _05313_, \oc8051_golden_model_1.ACC [1]);
  nor (_09541_, _09540_, _09539_);
  and (_09542_, _09541_, _09538_);
  and (_09543_, _09542_, _09536_);
  and (_09544_, _05326_, \oc8051_golden_model_1.SCON [1]);
  and (_09545_, _05328_, \oc8051_golden_model_1.IE [1]);
  nor (_09546_, _09545_, _09544_);
  and (_09547_, _04635_, \oc8051_golden_model_1.P0INREG [1]);
  and (_09548_, _05335_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_09549_, _09548_, _09547_);
  and (_09550_, _05332_, \oc8051_golden_model_1.P1INREG [1]);
  and (_09551_, _05337_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_09552_, _09551_, _09550_);
  and (_09553_, _09552_, _09549_);
  and (_09554_, _09553_, _09546_);
  and (_09555_, _09554_, _09543_);
  and (_09556_, _09555_, _04994_);
  nor (_09557_, _09556_, _09533_);
  nor (_09558_, _09557_, _09532_);
  and (_09559_, _04645_, _04385_);
  not (_09560_, _09559_);
  and (_09561_, _05316_, \oc8051_golden_model_1.PSW [4]);
  and (_09562_, _05321_, \oc8051_golden_model_1.B [4]);
  nor (_09563_, _09562_, _09561_);
  and (_09564_, _05319_, \oc8051_golden_model_1.IP [4]);
  and (_09565_, _05313_, \oc8051_golden_model_1.ACC [4]);
  nor (_09566_, _09565_, _09564_);
  and (_09567_, _09566_, _09563_);
  and (_09568_, _05326_, \oc8051_golden_model_1.SCON [4]);
  and (_09569_, _05328_, \oc8051_golden_model_1.IE [4]);
  nor (_09570_, _09569_, _09568_);
  and (_09571_, _05310_, \oc8051_golden_model_1.TCON [4]);
  and (_09572_, _05337_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_09573_, _09572_, _09571_);
  and (_09574_, _09573_, _09570_);
  and (_09575_, _05332_, \oc8051_golden_model_1.P1INREG [4]);
  not (_09576_, _09575_);
  and (_09577_, _04635_, \oc8051_golden_model_1.P0INREG [4]);
  and (_09578_, _05335_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_09579_, _09578_, _09577_);
  and (_09580_, _09579_, _09576_);
  and (_09581_, _09580_, _09574_);
  and (_09582_, _09581_, _09567_);
  and (_09583_, _09582_, _05193_);
  nor (_09584_, _09583_, _09560_);
  nor (_09585_, _05528_, _05347_);
  nor (_09586_, _09585_, _09584_);
  and (_09587_, _09586_, _09558_);
  not (_09588_, _04646_);
  and (_09589_, _05319_, \oc8051_golden_model_1.IP [0]);
  and (_09590_, _05321_, \oc8051_golden_model_1.B [0]);
  nor (_09591_, _09590_, _09589_);
  and (_09592_, _05316_, \oc8051_golden_model_1.PSW [0]);
  and (_09593_, _05313_, \oc8051_golden_model_1.ACC [0]);
  nor (_09594_, _09593_, _09592_);
  and (_09595_, _09594_, _09591_);
  and (_09596_, _05326_, \oc8051_golden_model_1.SCON [0]);
  and (_09597_, _05328_, \oc8051_golden_model_1.IE [0]);
  nor (_09598_, _09597_, _09596_);
  and (_09599_, _05310_, \oc8051_golden_model_1.TCON [0]);
  and (_09600_, _05337_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_09601_, _09600_, _09599_);
  and (_09602_, _09601_, _09598_);
  and (_09603_, _05332_, \oc8051_golden_model_1.P1INREG [0]);
  not (_09604_, _09603_);
  and (_09605_, _04635_, \oc8051_golden_model_1.P0INREG [0]);
  and (_09606_, _05335_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_09607_, _09606_, _09605_);
  and (_09608_, _09607_, _09604_);
  and (_09609_, _09608_, _09602_);
  and (_09610_, _09609_, _09595_);
  and (_09611_, _09610_, _05039_);
  nor (_09612_, _09611_, _09588_);
  and (_09613_, _04641_, _04385_);
  not (_09614_, _09613_);
  and (_09615_, _05319_, \oc8051_golden_model_1.IP [6]);
  and (_09616_, _05313_, \oc8051_golden_model_1.ACC [6]);
  nor (_09617_, _09616_, _09615_);
  and (_09618_, _05316_, \oc8051_golden_model_1.PSW [6]);
  and (_09619_, _05321_, \oc8051_golden_model_1.B [6]);
  nor (_09620_, _09619_, _09618_);
  and (_09621_, _09620_, _09617_);
  and (_09622_, _05337_, \oc8051_golden_model_1.P3INREG [6]);
  not (_09623_, _09622_);
  and (_09624_, _05332_, \oc8051_golden_model_1.P1INREG [6]);
  and (_09625_, _05335_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_09626_, _09625_, _09624_);
  and (_09627_, _09626_, _09623_);
  and (_09628_, _05326_, \oc8051_golden_model_1.SCON [6]);
  and (_09629_, _05328_, \oc8051_golden_model_1.IE [6]);
  nor (_09630_, _09629_, _09628_);
  and (_09631_, _05310_, \oc8051_golden_model_1.TCON [6]);
  and (_09632_, _04635_, \oc8051_golden_model_1.P0INREG [6]);
  nor (_09633_, _09632_, _09631_);
  and (_09634_, _09633_, _09630_);
  and (_09635_, _09634_, _09627_);
  and (_09636_, _09635_, _09621_);
  and (_09637_, _09636_, _04791_);
  nor (_09638_, _09637_, _09614_);
  nor (_09639_, _09638_, _09612_);
  not (_09640_, _04695_);
  and (_09641_, _05319_, \oc8051_golden_model_1.IP [3]);
  and (_09642_, _05321_, \oc8051_golden_model_1.B [3]);
  nor (_09643_, _09642_, _09641_);
  and (_09644_, _05316_, \oc8051_golden_model_1.PSW [3]);
  and (_09645_, _05313_, \oc8051_golden_model_1.ACC [3]);
  nor (_09646_, _09645_, _09644_);
  and (_09647_, _09646_, _09643_);
  and (_09648_, _05337_, \oc8051_golden_model_1.P3INREG [3]);
  not (_09649_, _09648_);
  and (_09650_, _05332_, \oc8051_golden_model_1.P1INREG [3]);
  and (_09651_, _05335_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_09652_, _09651_, _09650_);
  and (_09653_, _09652_, _09649_);
  and (_09654_, _05326_, \oc8051_golden_model_1.SCON [3]);
  and (_09655_, _05328_, \oc8051_golden_model_1.IE [3]);
  nor (_09656_, _09655_, _09654_);
  and (_09657_, _05310_, \oc8051_golden_model_1.TCON [3]);
  and (_09658_, _04635_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_09659_, _09658_, _09657_);
  and (_09660_, _09659_, _09656_);
  and (_09661_, _09660_, _09653_);
  and (_09662_, _09661_, _09647_);
  and (_09663_, _09662_, _04946_);
  nor (_09664_, _09663_, _09640_);
  and (_09665_, _04636_, _04385_);
  not (_09666_, _09665_);
  and (_09667_, _05326_, \oc8051_golden_model_1.SCON [5]);
  and (_09668_, _05328_, \oc8051_golden_model_1.IE [5]);
  nor (_09669_, _09668_, _09667_);
  and (_09670_, _05310_, \oc8051_golden_model_1.TCON [5]);
  and (_09671_, _05337_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_09672_, _09671_, _09670_);
  and (_09673_, _09672_, _09669_);
  and (_09674_, _05319_, \oc8051_golden_model_1.IP [5]);
  and (_09675_, _05321_, \oc8051_golden_model_1.B [5]);
  nor (_09676_, _09675_, _09674_);
  and (_09677_, _05316_, \oc8051_golden_model_1.PSW [5]);
  and (_09678_, _05313_, \oc8051_golden_model_1.ACC [5]);
  nor (_09679_, _09678_, _09677_);
  and (_09680_, _09679_, _09676_);
  and (_09681_, _05332_, \oc8051_golden_model_1.P1INREG [5]);
  and (_09682_, _05335_, \oc8051_golden_model_1.P2INREG [5]);
  and (_09683_, _04635_, \oc8051_golden_model_1.P0INREG [5]);
  or (_09684_, _09683_, _09682_);
  nor (_09685_, _09684_, _09681_);
  and (_09686_, _09685_, _09680_);
  and (_09687_, _09686_, _09673_);
  and (_09688_, _09687_, _04895_);
  nor (_09689_, _09688_, _09666_);
  nor (_09690_, _09689_, _09664_);
  and (_09691_, _09690_, _09639_);
  and (_09692_, _09691_, _09587_);
  and (_09693_, _09692_, _08949_);
  nor (_09694_, _09692_, _06195_);
  or (_09695_, _09694_, _03223_);
  or (_09696_, _09695_, _09693_);
  and (_09697_, _09696_, _08803_);
  and (_09698_, _09697_, _09507_);
  or (_09699_, _09698_, _08804_);
  nand (_09700_, _09699_, _08789_);
  nor (_09701_, _08789_, _06206_);
  nor (_09702_, _09701_, _08115_);
  nand (_09703_, _09702_, _09700_);
  and (_09704_, _08802_, _08115_);
  nor (_09705_, _09704_, _02890_);
  and (_09706_, _09705_, _09703_);
  and (_09707_, _04630_, _02890_);
  or (_09708_, _09707_, _09706_);
  nand (_09709_, _09708_, _08788_);
  nor (_09710_, _06206_, _08788_);
  nor (_09711_, _09710_, _02889_);
  nand (_09712_, _09711_, _09709_);
  nor (_09713_, _09692_, _09005_);
  and (_09714_, _09692_, _08943_);
  nor (_09715_, _09714_, _09713_);
  and (_09716_, _09715_, _02889_);
  and (_09717_, _03009_, _02504_);
  not (_09718_, _09717_);
  and (_09719_, _03007_, _02504_);
  nor (_09720_, _09719_, _03591_);
  and (_09721_, _09720_, _09718_);
  and (_09722_, _04130_, _09721_);
  and (_09723_, _09722_, _04105_);
  and (_09724_, _09723_, _05809_);
  not (_09725_, _09724_);
  nor (_09726_, _09725_, _09716_);
  nand (_09727_, _09726_, _09712_);
  nor (_09728_, _09724_, _08802_);
  nor (_09729_, _09728_, _03174_);
  nand (_09730_, _09729_, _09727_);
  and (_09731_, _06206_, _03174_);
  nor (_09732_, _08160_, _08155_);
  not (_09733_, _09732_);
  nor (_09734_, _09733_, _09731_);
  nand (_09735_, _09734_, _09730_);
  nor (_09736_, _09732_, _08802_);
  nor (_09737_, _09736_, _03034_);
  and (_09738_, _09737_, _09735_);
  nor (_09739_, _06185_, _02763_);
  or (_09740_, _09739_, _02505_);
  or (_09741_, _09740_, _09738_);
  not (_09742_, _02505_);
  nor (_09743_, _06206_, _09742_);
  nor (_09744_, _09743_, _02799_);
  nand (_09745_, _09744_, _09741_);
  and (_09746_, _09715_, _02799_);
  and (_09747_, _05257_, _06161_);
  not (_09748_, _09747_);
  nor (_09749_, _09748_, _09746_);
  nand (_09750_, _09749_, _09745_);
  nor (_09751_, _09747_, _08802_);
  nor (_09752_, _09751_, _02887_);
  nand (_09753_, _09752_, _09750_);
  and (_09754_, _06206_, _02887_);
  nor (_09755_, _08184_, _08177_);
  not (_09756_, _09755_);
  nor (_09757_, _09756_, _09754_);
  nand (_09758_, _09757_, _09753_);
  nor (_09759_, _09755_, _08802_);
  nor (_09760_, _09759_, _03036_);
  and (_09761_, _09760_, _09758_);
  nor (_09762_, _03038_, _02763_);
  or (_09763_, _09762_, _09761_);
  and (_09764_, _09763_, _02500_);
  and (_09765_, _06206_, _02499_);
  or (_09766_, _09765_, _09764_);
  and (_09767_, _09766_, _08787_);
  and (_09768_, _08802_, _08786_);
  or (_09769_, _09768_, _09767_);
  or (_09770_, _09769_, _34659_);
  or (_09771_, _34655_, \oc8051_golden_model_1.PC [15]);
  and (_09772_, _09771_, _35796_);
  and (_35842_[15], _09772_, _09770_);
  nor (_09773_, _04718_, _07288_);
  not (_09774_, _09773_);
  nand (_09775_, _05772_, _04718_);
  and (_09776_, _09775_, _09774_);
  or (_09777_, _09776_, _07150_);
  not (_09778_, _02928_);
  not (_09779_, _04718_);
  or (_09780_, _05740_, _09779_);
  and (_09781_, _09780_, _09774_);
  or (_09782_, _09781_, _02839_);
  or (_09783_, _09779_, _04630_);
  and (_09784_, _09783_, _09774_);
  and (_09785_, _09784_, _05535_);
  nand (_09786_, _07655_, _07653_);
  or (_09787_, _09786_, _07552_);
  or (_09788_, _09787_, _05497_);
  and (_09789_, _07651_, _07647_);
  nor (_09790_, _09789_, _07645_);
  and (_09791_, _07968_, _07647_);
  not (_09792_, _09791_);
  nor (_09793_, _09792_, _07712_);
  not (_09794_, _09793_);
  and (_09795_, _09794_, _09790_);
  not (_09796_, _09795_);
  and (_09797_, _09796_, _09788_);
  or (_09798_, _09797_, _02991_);
  not (_09799_, _02941_);
  or (_09800_, _09692_, _09799_);
  nand (_09801_, _09249_, _07288_);
  not (_09802_, _07700_);
  nor (_09803_, _09289_, _09802_);
  or (_09804_, _09803_, _07698_);
  nand (_09805_, _09804_, _09287_);
  and (_09806_, _09286_, _08089_);
  nor (_09807_, _09806_, _09284_);
  nand (_09808_, _09807_, _09805_);
  nand (_09809_, _09808_, _09296_);
  and (_09810_, _08081_, _08084_);
  or (_09811_, _09810_, _08079_);
  nand (_09812_, _09811_, _09295_);
  or (_09813_, _05497_, \oc8051_golden_model_1.ACC [7]);
  nand (_09814_, _08076_, _09294_);
  and (_09815_, _09814_, _09813_);
  and (_09816_, _09815_, _09812_);
  and (_09817_, _09816_, _09809_);
  or (_09818_, _09297_, _09299_);
  or (_09819_, _09818_, _09817_);
  or (_09820_, _03687_, \oc8051_golden_model_1.ACC [1]);
  and (_09821_, _03687_, \oc8051_golden_model_1.ACC [1]);
  and (_09822_, _02837_, \oc8051_golden_model_1.ACC [0]);
  or (_09823_, _09822_, _09821_);
  nand (_09824_, _09823_, _09820_);
  nand (_09825_, _09824_, _09270_);
  nor (_09826_, _02794_, _02625_);
  and (_09827_, _02794_, _02625_);
  nor (_09828_, _03356_, \oc8051_golden_model_1.ACC [2]);
  nor (_09829_, _09828_, _09827_);
  or (_09830_, _09829_, _09826_);
  nand (_09831_, _09830_, _09825_);
  nand (_09832_, _09831_, _09268_);
  and (_09833_, _03220_, \oc8051_golden_model_1.ACC [5]);
  nor (_09834_, _03220_, \oc8051_golden_model_1.ACC [5]);
  nor (_09835_, _03647_, \oc8051_golden_model_1.ACC [4]);
  nor (_09836_, _09835_, _09834_);
  nor (_09837_, _09836_, _09833_);
  nand (_09838_, _09837_, _09267_);
  or (_09839_, _02763_, \oc8051_golden_model_1.ACC [7]);
  or (_09840_, _02924_, \oc8051_golden_model_1.ACC [6]);
  or (_09841_, _09840_, _07867_);
  and (_09842_, _09841_, _09839_);
  and (_09843_, _09842_, _09838_);
  and (_09844_, _09843_, _09832_);
  or (_09845_, _09844_, _09279_);
  or (_09846_, _09845_, _09276_);
  and (_09847_, _09846_, _09819_);
  and (_09848_, _09847_, _09801_);
  and (_09849_, _05474_, _04718_);
  nor (_09850_, _09849_, _09773_);
  and (_09851_, _09850_, _02948_);
  and (_09852_, _04718_, \oc8051_golden_model_1.ACC [7]);
  nor (_09853_, _09852_, _09773_);
  or (_09854_, _09853_, _04194_);
  or (_09855_, _03845_, _07288_);
  and (_09856_, _09855_, _03006_);
  and (_09857_, _09856_, _09854_);
  or (_09858_, _09857_, _07405_);
  or (_09859_, _09858_, _09851_);
  nor (_09860_, _07451_, \oc8051_golden_model_1.PSW [7]);
  not (_09861_, _09860_);
  nor (_09862_, _09861_, _07461_);
  not (_09863_, _09862_);
  and (_09864_, _09863_, _03028_);
  nor (_09865_, _09864_, _07439_);
  or (_09866_, _09865_, _02596_);
  and (_09867_, _09866_, _09859_);
  nor (_09868_, _05316_, _07288_);
  not (_09869_, _09868_);
  nand (_09870_, _05348_, _05316_);
  and (_09871_, _09870_, _09869_);
  and (_09872_, _09871_, _02884_);
  or (_09873_, _09872_, _02946_);
  or (_09874_, _09873_, _09867_);
  or (_09875_, _09784_, _07474_);
  and (_09876_, _09875_, _02992_);
  and (_09877_, _09876_, _09874_);
  nand (_09878_, _09853_, _02880_);
  nand (_09879_, _07439_, _02875_);
  nand (_09880_, _09879_, _09878_);
  or (_09881_, _09880_, _09877_);
  and (_09882_, _05344_, _05316_);
  nor (_09883_, _09882_, _09868_);
  or (_09884_, _09883_, _02987_);
  and (_09885_, _09884_, _09209_);
  and (_09886_, _09885_, _09881_);
  nor (_09887_, _09237_, _09234_);
  or (_09888_, _09235_, _09887_);
  nand (_09889_, _09888_, _09233_);
  or (_09890_, _09230_, _09229_);
  nand (_09891_, _09890_, _09889_);
  nand (_09892_, _09891_, _09226_);
  and (_09893_, _09221_, _09222_);
  or (_09894_, _09893_, _09220_);
  nand (_09895_, _09894_, _09218_);
  and (_09896_, _09216_, _04631_);
  nor (_09897_, _09896_, _09213_);
  and (_09898_, _09897_, _09895_);
  and (_09899_, _09898_, _09892_);
  or (_09900_, _09899_, _09242_);
  and (_09901_, _09900_, _09210_);
  or (_09902_, _09901_, _08985_);
  or (_09903_, _09902_, _09886_);
  not (_09904_, _08972_);
  or (_09905_, _08974_, _09904_);
  or (_09906_, _08966_, _08969_);
  and (_09907_, _09906_, _08965_);
  and (_09908_, _09907_, _08978_);
  nand (_09909_, _09908_, _09905_);
  nand (_09910_, _09909_, _08964_);
  nand (_09911_, _08961_, _08958_);
  and (_09912_, _08956_, _09911_);
  nand (_09913_, _09912_, _08957_);
  and (_09914_, _08951_, _08953_);
  or (_09915_, _09914_, _05514_);
  and (_09916_, _09915_, _09913_);
  and (_09917_, _09916_, _09910_);
  and (_09918_, _08980_, _08964_);
  or (_09919_, _08986_, _09918_);
  or (_09920_, _09919_, _09917_);
  and (_09921_, _09920_, _09903_);
  or (_09922_, _09921_, _09252_);
  and (_09923_, _09922_, _09848_);
  or (_09924_, _09923_, _03434_);
  and (_09925_, _09869_, _05501_);
  or (_09926_, _09925_, _06246_);
  or (_09927_, _09926_, _09871_);
  and (_09928_, _04635_, \oc8051_golden_model_1.P0 [2]);
  and (_09929_, _05332_, \oc8051_golden_model_1.P1 [2]);
  nor (_09930_, _09929_, _09928_);
  and (_09931_, _05337_, \oc8051_golden_model_1.P3 [2]);
  and (_09932_, _05335_, \oc8051_golden_model_1.P2 [2]);
  or (_09933_, _09932_, _09931_);
  nor (_09934_, _09933_, _09525_);
  and (_09935_, _09934_, _09515_);
  and (_09936_, _09935_, _09524_);
  and (_09937_, _09936_, _09930_);
  and (_09938_, _09937_, _05087_);
  nor (_09939_, _09938_, _09508_);
  and (_09940_, _05335_, \oc8051_golden_model_1.P2 [1]);
  and (_09941_, _05337_, \oc8051_golden_model_1.P3 [1]);
  nor (_09942_, _09941_, _09940_);
  and (_09943_, _04635_, \oc8051_golden_model_1.P0 [1]);
  and (_09944_, _05332_, \oc8051_golden_model_1.P1 [1]);
  nor (_09945_, _09944_, _09943_);
  and (_09946_, _09945_, _09942_);
  and (_09947_, _09946_, _09546_);
  and (_09948_, _09947_, _09543_);
  and (_09949_, _09948_, _04994_);
  nor (_09950_, _09949_, _09533_);
  nor (_09951_, _09950_, _09939_);
  and (_09952_, _05337_, \oc8051_golden_model_1.P3 [4]);
  not (_09953_, _09952_);
  and (_09954_, _05335_, \oc8051_golden_model_1.P2 [4]);
  nor (_09955_, _09954_, _09571_);
  and (_09956_, _09955_, _09953_);
  and (_09957_, _04635_, \oc8051_golden_model_1.P0 [4]);
  and (_09958_, _05332_, \oc8051_golden_model_1.P1 [4]);
  nor (_09959_, _09958_, _09957_);
  and (_09960_, _09959_, _09570_);
  and (_09961_, _09960_, _09956_);
  and (_09962_, _09961_, _09567_);
  and (_09963_, _09962_, _05193_);
  nor (_09964_, _09560_, _09963_);
  nor (_09965_, _09964_, _05501_);
  and (_09966_, _09965_, _09951_);
  and (_09967_, _04635_, \oc8051_golden_model_1.P0 [0]);
  and (_09968_, _05332_, \oc8051_golden_model_1.P1 [0]);
  nor (_09969_, _09968_, _09967_);
  and (_09970_, _05337_, \oc8051_golden_model_1.P3 [0]);
  and (_09971_, _05335_, \oc8051_golden_model_1.P2 [0]);
  or (_09972_, _09971_, _09970_);
  nor (_09973_, _09972_, _09599_);
  and (_09974_, _09973_, _09595_);
  and (_09975_, _09974_, _09598_);
  and (_09976_, _09975_, _09969_);
  and (_09977_, _09976_, _05039_);
  nor (_09978_, _09977_, _09588_);
  and (_09979_, _04635_, \oc8051_golden_model_1.P0 [6]);
  and (_09980_, _05332_, \oc8051_golden_model_1.P1 [6]);
  nor (_09981_, _09980_, _09979_);
  and (_09982_, _05337_, \oc8051_golden_model_1.P3 [6]);
  and (_09983_, _05335_, \oc8051_golden_model_1.P2 [6]);
  or (_09984_, _09983_, _09982_);
  nor (_09985_, _09984_, _09631_);
  and (_09986_, _09985_, _09621_);
  and (_09987_, _09986_, _09630_);
  and (_09988_, _09987_, _09981_);
  and (_09989_, _09988_, _04791_);
  nor (_09990_, _09614_, _09989_);
  nor (_09991_, _09990_, _09978_);
  and (_09992_, _04635_, \oc8051_golden_model_1.P0 [3]);
  and (_09993_, _05332_, \oc8051_golden_model_1.P1 [3]);
  nor (_09994_, _09993_, _09992_);
  and (_09995_, _05337_, \oc8051_golden_model_1.P3 [3]);
  and (_09996_, _05335_, \oc8051_golden_model_1.P2 [3]);
  or (_09997_, _09996_, _09995_);
  nor (_09998_, _09997_, _09657_);
  and (_09999_, _09998_, _09647_);
  and (_10000_, _09999_, _09656_);
  and (_10001_, _10000_, _09994_);
  and (_10002_, _10001_, _04946_);
  nor (_10003_, _10002_, _09640_);
  and (_10004_, _04635_, \oc8051_golden_model_1.P0 [5]);
  and (_10005_, _05332_, \oc8051_golden_model_1.P1 [5]);
  nor (_10006_, _10005_, _10004_);
  and (_10007_, _05337_, \oc8051_golden_model_1.P3 [5]);
  and (_10008_, _05335_, \oc8051_golden_model_1.P2 [5]);
  or (_10009_, _10008_, _10007_);
  nor (_10010_, _10009_, _09670_);
  and (_10011_, _10010_, _09680_);
  and (_10012_, _10011_, _09669_);
  and (_10013_, _10012_, _10006_);
  and (_10014_, _10013_, _04895_);
  nor (_10015_, _09666_, _10014_);
  nor (_10016_, _10015_, _10003_);
  and (_10017_, _10016_, _09991_);
  and (_10018_, _10017_, _09966_);
  and (_10019_, _02937_, \oc8051_golden_model_1.PSW [7]);
  nand (_10020_, _10019_, _10018_);
  and (_10021_, _10020_, _09927_);
  and (_10022_, _10021_, _09924_);
  or (_10023_, _06252_, _02941_);
  or (_10024_, _10023_, _10022_);
  and (_10025_, _10024_, _09800_);
  or (_10026_, _10025_, _02940_);
  nor (_10027_, _03767_, _03455_);
  nand (_10028_, _03448_, _04138_);
  and (_10029_, _10028_, _10027_);
  not (_10030_, _02940_);
  nor (_10031_, _10018_, \oc8051_golden_model_1.PSW [7]);
  or (_10032_, _10031_, _10030_);
  and (_10033_, _10032_, _10029_);
  and (_10034_, _10033_, _10026_);
  and (_10035_, _02962_, _02864_);
  and (_10036_, _07244_, _05258_);
  and (_10037_, _07249_, _07243_);
  nor (_10038_, _10037_, _07241_);
  not (_10039_, _10038_);
  and (_10040_, _07250_, _07243_);
  not (_10041_, _10040_);
  nor (_10042_, _10041_, _07529_);
  nor (_10043_, _10042_, _10039_);
  nor (_10044_, _10043_, _10036_);
  or (_10045_, _10044_, _10035_);
  and (_10046_, _10045_, _07400_);
  or (_10047_, _10046_, _10034_);
  nor (_10048_, _07397_, _10035_);
  and (_10049_, _10044_, _07507_);
  or (_10050_, _10049_, _10048_);
  and (_10051_, _10050_, _10047_);
  and (_10052_, _07335_, _07331_);
  nor (_10053_, _10052_, _07329_);
  not (_10054_, _10053_);
  and (_10055_, _07938_, _07331_);
  not (_10056_, _10055_);
  nor (_10057_, _10056_, _07391_);
  nor (_10058_, _10057_, _10054_);
  or (_10059_, _07507_, _07327_);
  nor (_10060_, _10059_, _10058_);
  or (_10061_, _10060_, _02979_);
  or (_10062_, _10061_, _10051_);
  and (_10063_, _10062_, _09798_);
  or (_10064_, _10063_, _07540_);
  nand (_10065_, _07723_, _04720_);
  and (_10066_, _07735_, _07731_);
  nor (_10067_, _10066_, _07729_);
  and (_10068_, _07999_, _07731_);
  not (_10069_, _10068_);
  nor (_10070_, _10069_, _07794_);
  not (_10071_, _10070_);
  and (_10072_, _10071_, _10067_);
  not (_10073_, _10072_);
  and (_10074_, _10073_, _10065_);
  or (_10075_, _10074_, _07541_);
  and (_10076_, _10075_, _02859_);
  and (_10077_, _10076_, _10064_);
  or (_10078_, _10077_, _09785_);
  and (_10079_, _10078_, _02842_);
  or (_10080_, _05810_, _09779_);
  nor (_10081_, _09773_, _02842_);
  and (_10082_, _10081_, _10080_);
  or (_10083_, _10082_, _02567_);
  or (_10084_, _10083_, _10079_);
  and (_10085_, _10084_, _09782_);
  or (_10086_, _06786_, _02930_);
  or (_10087_, _10086_, _10085_);
  or (_10088_, _10018_, _07288_);
  or (_10089_, _10088_, _03508_);
  and (_10090_, _10089_, _07140_);
  and (_10091_, _10090_, _10087_);
  and (_10092_, _05549_, _04718_);
  nor (_10093_, _10092_, _09773_);
  and (_10094_, _10093_, _02834_);
  or (_10095_, _10094_, _10091_);
  and (_10096_, _10095_, _09778_);
  and (_10097_, _10018_, _07288_);
  and (_10098_, _10097_, _02928_);
  or (_10099_, _10098_, _10096_);
  and (_10100_, _10099_, _07139_);
  nand (_10101_, _05764_, _04718_);
  nor (_10102_, _09773_, _07139_);
  and (_10103_, _10102_, _10101_);
  or (_10104_, _10103_, _03148_);
  or (_10105_, _10104_, _10100_);
  nand (_10106_, _10105_, _09777_);
  nand (_10107_, _10106_, _03138_);
  and (_10108_, _09774_, _04739_);
  or (_10109_, _09853_, _06213_);
  or (_10110_, _10093_, _03023_);
  and (_10111_, _10110_, _10109_);
  or (_10112_, _10111_, _10108_);
  and (_10113_, _10112_, _03043_);
  and (_10114_, _10113_, _10107_);
  or (_10115_, _05763_, _09779_);
  nor (_10116_, _09773_, _03043_);
  and (_10117_, _10116_, _10115_);
  or (_10118_, _10117_, _03143_);
  or (_10119_, _10118_, _10114_);
  or (_10120_, _05771_, _09779_);
  and (_10121_, _10120_, _09774_);
  or (_10122_, _10121_, _07161_);
  and (_10123_, _10122_, _07234_);
  and (_10124_, _10123_, _10119_);
  nor (_10125_, _07240_, _05364_);
  or (_10126_, _10125_, _07305_);
  or (_10127_, _10126_, _10036_);
  nor (_10128_, _10127_, _07234_);
  or (_10129_, _10128_, _10124_);
  and (_10130_, _10129_, _07936_);
  and (_10131_, _07328_, \oc8051_golden_model_1.ACC [7]);
  nor (_10132_, _10131_, _07958_);
  nor (_10133_, _07936_, _07327_);
  and (_10134_, _10133_, _10132_);
  or (_10135_, _10134_, _03133_);
  or (_10136_, _10135_, _10130_);
  nor (_10137_, _07644_, _05364_);
  nor (_10138_, _10137_, _07989_);
  and (_10139_, _10138_, _09788_);
  or (_10140_, _10139_, _03134_);
  and (_10141_, _10140_, _07997_);
  and (_10142_, _10141_, _10136_);
  nor (_10143_, _07728_, _05364_);
  nor (_10144_, _10143_, _08020_);
  and (_10145_, _10065_, _07964_);
  and (_10146_, _10145_, _10144_);
  or (_10147_, _10146_, _07995_);
  or (_10148_, _10147_, _10142_);
  nand (_10149_, _07995_, \oc8051_golden_model_1.ACC [7]);
  and (_10150_, _10149_, _07189_);
  and (_10151_, _10150_, _10148_);
  nand (_10152_, _07223_, _07192_);
  not (_10153_, _07189_);
  nor (_10154_, _07193_, _07191_);
  or (_10155_, _10154_, _07190_);
  and (_10156_, _10155_, _10153_);
  and (_10157_, _10156_, _10152_);
  or (_10158_, _10157_, _10151_);
  and (_10159_, _10158_, _08031_);
  nand (_10160_, _08062_, _07856_);
  nor (_10161_, _08032_, _07855_);
  or (_10162_, _10161_, _07854_);
  and (_10163_, _10162_, _07185_);
  and (_10164_, _10163_, _10160_);
  or (_10165_, _10164_, _02892_);
  or (_10166_, _10165_, _10159_);
  not (_10167_, _08071_);
  not (_10168_, _03359_);
  not (_10169_, _08072_);
  and (_10170_, _08107_, _10169_);
  nor (_10171_, _10170_, _10168_);
  nand (_10172_, _10171_, _10167_);
  and (_10173_, _10172_, _08117_);
  and (_10174_, _10173_, _10166_);
  not (_10175_, _07865_);
  nor (_10176_, _08145_, _07866_);
  nor (_10177_, _10176_, _08117_);
  and (_10178_, _10177_, _10175_);
  nor (_10179_, _10178_, _10174_);
  nor (_10180_, _10179_, _03174_);
  and (_10181_, _09850_, _03174_);
  nor (_10182_, _10181_, _08160_);
  not (_10183_, _10182_);
  nor (_10184_, _10183_, _10180_);
  and (_10185_, _08160_, \oc8051_golden_model_1.ACC [0]);
  or (_10186_, _10185_, _10184_);
  and (_10187_, _10186_, _03183_);
  nor (_10188_, _09883_, _03183_);
  or (_10189_, _10188_, _10187_);
  and (_10190_, _10189_, _02888_);
  and (_10191_, _05246_, _04718_);
  nor (_10192_, _10191_, _09773_);
  nor (_10193_, _10192_, _02888_);
  or (_10194_, _10193_, _10190_);
  or (_10195_, _10194_, _34659_);
  or (_10196_, _34655_, \oc8051_golden_model_1.PSW [7]);
  and (_10197_, _10196_, _35796_);
  and (_35843_[7], _10197_, _10195_);
  and (_35841_[7], \oc8051_golden_model_1.PCON [7], _35796_);
  and (_35844_[7], \oc8051_golden_model_1.SBUF [7], _35796_);
  and (_35845_[7], \oc8051_golden_model_1.SCON [7], _35796_);
  not (_10198_, \oc8051_golden_model_1.SP [7]);
  nor (_10199_, _04638_, _10198_);
  and (_10200_, _05246_, _04638_);
  nor (_10201_, _10200_, _10199_);
  nor (_10202_, _10201_, _02888_);
  and (_10203_, _05772_, _04638_);
  nor (_10204_, _10203_, _10199_);
  nor (_10205_, _10204_, _07150_);
  not (_10206_, _04638_);
  nor (_10207_, _10206_, _04630_);
  nor (_10208_, _10207_, _10199_);
  nor (_10209_, _10208_, _02859_);
  or (_10210_, _10209_, _02841_);
  and (_10211_, _04219_, \oc8051_golden_model_1.SP [4]);
  and (_10212_, _10211_, \oc8051_golden_model_1.SP [5]);
  and (_10213_, _10212_, \oc8051_golden_model_1.SP [6]);
  and (_10214_, _10213_, \oc8051_golden_model_1.SP [0]);
  nor (_10215_, _10214_, \oc8051_golden_model_1.SP [7]);
  and (_10216_, _10214_, \oc8051_golden_model_1.SP [7]);
  nor (_10217_, _10216_, _10215_);
  and (_10218_, _10217_, _02876_);
  not (_10219_, _04135_);
  and (_10220_, _04638_, \oc8051_golden_model_1.ACC [7]);
  nor (_10221_, _10220_, _10199_);
  nor (_10222_, _10221_, _04194_);
  nor (_10223_, _03845_, _10198_);
  or (_10224_, _10223_, _03849_);
  nor (_10225_, _10224_, _10222_);
  nor (_10226_, _10213_, \oc8051_golden_model_1.SP [7]);
  and (_10227_, _10213_, \oc8051_golden_model_1.SP [7]);
  nor (_10228_, _10227_, _10226_);
  nor (_10229_, _10228_, _02603_);
  nor (_10230_, _10229_, _10225_);
  and (_10231_, _10230_, _03006_);
  and (_10232_, _05474_, _04638_);
  nor (_10233_, _10232_, _10199_);
  nor (_10234_, _10233_, _03006_);
  or (_10235_, _10234_, _10231_);
  and (_10236_, _10235_, _02597_);
  not (_10237_, _10228_);
  nor (_10238_, _10237_, _02597_);
  or (_10239_, _10238_, _10236_);
  and (_10240_, _10239_, _07474_);
  not (_10241_, \oc8051_golden_model_1.SP [6]);
  not (_10242_, \oc8051_golden_model_1.SP [5]);
  not (_10243_, \oc8051_golden_model_1.SP [4]);
  and (_10244_, _05415_, _10243_);
  and (_10245_, _10244_, _10242_);
  and (_10246_, _10245_, _10241_);
  and (_10247_, _10246_, _02868_);
  nor (_10248_, _10247_, \oc8051_golden_model_1.SP [7]);
  and (_10249_, _10247_, \oc8051_golden_model_1.SP [7]);
  nor (_10250_, _10249_, _10248_);
  and (_10251_, _10250_, _10206_);
  nor (_10252_, _10251_, _10207_);
  nor (_10253_, _10252_, _07474_);
  or (_10254_, _10253_, _10240_);
  and (_10255_, _10254_, _02992_);
  nor (_10256_, _10221_, _02992_);
  or (_10257_, _10256_, _10255_);
  and (_10258_, _10257_, _03962_);
  or (_10259_, _10258_, _10219_);
  nor (_10260_, _10259_, _10218_);
  nor (_10261_, _10228_, _04135_);
  nor (_10262_, _10261_, _05535_);
  not (_10263_, _10262_);
  nor (_10264_, _10263_, _10260_);
  nor (_10265_, _10264_, _10210_);
  and (_10266_, _05461_, _04638_);
  nor (_10267_, _10199_, _02842_);
  not (_10268_, _10267_);
  nor (_10269_, _10268_, _10266_);
  nor (_10270_, _10269_, _02567_);
  not (_10271_, _10270_);
  nor (_10272_, _10271_, _10265_);
  nor (_10273_, _05740_, _10206_);
  nor (_10274_, _10273_, _10199_);
  nor (_10275_, _10274_, _02839_);
  or (_10276_, _10275_, _02834_);
  or (_10277_, _10276_, _10272_);
  and (_10278_, _05549_, _04638_);
  nor (_10279_, _10278_, _10199_);
  nand (_10280_, _10279_, _02834_);
  and (_10281_, _10280_, _10277_);
  nor (_10282_, _10281_, _02522_);
  and (_10283_, _10237_, _02522_);
  nor (_10284_, _10283_, _10282_);
  and (_10285_, _10284_, _07139_);
  and (_10286_, _05764_, _04638_);
  nor (_10287_, _10286_, _10199_);
  nor (_10288_, _10287_, _07139_);
  or (_10289_, _10288_, _10285_);
  and (_10290_, _10289_, _07150_);
  nor (_10291_, _10290_, _10205_);
  nor (_10292_, _10291_, _03022_);
  nor (_10293_, _10199_, _04740_);
  not (_10294_, _10293_);
  nor (_10295_, _10279_, _03023_);
  and (_10296_, _10295_, _10294_);
  nor (_10297_, _10296_, _10292_);
  nor (_10298_, _10297_, _09463_);
  and (_10299_, _10228_, _02530_);
  or (_10300_, _10293_, _06213_);
  nor (_10301_, _10300_, _10221_);
  or (_10302_, _10301_, _10299_);
  or (_10303_, _10302_, _03042_);
  nor (_10304_, _10303_, _10298_);
  nor (_10305_, _05763_, _10206_);
  nor (_10306_, _10305_, _10199_);
  and (_10307_, _10306_, _03042_);
  nor (_10308_, _10307_, _10304_);
  nor (_10309_, _10308_, _03143_);
  nor (_10310_, _05771_, _10206_);
  or (_10311_, _10199_, _07161_);
  nor (_10312_, _10311_, _10310_);
  or (_10313_, _10312_, _03155_);
  nor (_10314_, _10313_, _10309_);
  nor (_10315_, _10246_, \oc8051_golden_model_1.SP [7]);
  and (_10316_, _10246_, \oc8051_golden_model_1.SP [7]);
  nor (_10317_, _10316_, _10315_);
  and (_10318_, _10317_, _03155_);
  or (_10319_, _10318_, _02528_);
  nor (_10320_, _10319_, _10314_);
  and (_10321_, _10237_, _02528_);
  nor (_10322_, _10321_, _10320_);
  and (_10323_, _10322_, _02891_);
  and (_10324_, _10317_, _02890_);
  or (_10325_, _10324_, _10323_);
  and (_10326_, _10325_, _03179_);
  nor (_10327_, _10233_, _03179_);
  or (_10328_, _10327_, _04150_);
  nor (_10329_, _10328_, _10326_);
  nor (_10330_, _10228_, _03936_);
  nor (_10331_, _10330_, _02887_);
  not (_10332_, _10331_);
  nor (_10333_, _10332_, _10329_);
  nor (_10334_, _10333_, _10202_);
  nand (_10335_, _10334_, _34655_);
  or (_10336_, _34655_, \oc8051_golden_model_1.SP [7]);
  and (_10337_, _10336_, _35796_);
  and (_35846_[7], _10337_, _10335_);
  and (_35847_[7], \oc8051_golden_model_1.TCON [7], _35796_);
  and (_35848_[7], \oc8051_golden_model_1.TH0 [7], _35796_);
  and (_35849_[7], \oc8051_golden_model_1.TH1 [7], _35796_);
  and (_35850_[7], \oc8051_golden_model_1.TL0 [7], _35796_);
  and (_35851_[7], \oc8051_golden_model_1.TL1 [7], _35796_);
  and (_35852_[7], \oc8051_golden_model_1.TMOD [7], _35796_);
  nor (_10338_, _09150_, _09134_);
  nor (_10339_, _10338_, _05364_);
  or (_10340_, _10339_, _34659_);
  or (_10341_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [7]);
  and (_10342_, _10341_, _35796_);
  and (_35854_[7], _10342_, _10340_);
  or (_10343_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [15]);
  and (_10344_, _10343_, _35796_);
  nor (_10345_, _09150_, _07433_);
  nor (_10346_, _10345_, _08295_);
  or (_10347_, _10346_, _34659_);
  and (_35853_[15], _10347_, _10344_);
  and (_10348_, _34659_, \oc8051_golden_model_1.P0INREG [7]);
  or (_10349_, _10348_, _00478_);
  and (_35833_[7], _10349_, _35796_);
  and (_10350_, _34659_, \oc8051_golden_model_1.P1INREG [7]);
  or (_10351_, _10350_, _00553_);
  and (_35835_[7], _10351_, _35796_);
  and (_10352_, _34659_, \oc8051_golden_model_1.P2INREG [7]);
  or (_10353_, _10352_, _00683_);
  and (_35837_[7], _10353_, _35796_);
  and (_10354_, _34659_, \oc8051_golden_model_1.P3INREG [7]);
  or (_10355_, _10354_, _00616_);
  and (_35839_[7], _10355_, _35796_);
  nor (_10356_, _04563_, _04127_);
  nor (_10357_, _10356_, _04564_);
  nor (_10358_, _04563_, _04540_);
  nor (_10359_, _10358_, _04567_);
  and (_10360_, _10359_, _04562_);
  and (_10361_, _10360_, _10357_);
  not (_10362_, _10361_);
  nand (_10363_, _02505_, _02247_);
  not (_10364_, _05785_);
  nor (_10365_, _05085_, _05660_);
  nor (_10366_, _10365_, _05786_);
  nor (_10367_, _05085_, \oc8051_golden_model_1.ACC [0]);
  and (_10368_, _05085_, \oc8051_golden_model_1.ACC [0]);
  nor (_10369_, _10368_, _10367_);
  and (_10370_, _10369_, _05762_);
  and (_10371_, _05085_, _05660_);
  nor (_10372_, _10371_, _10365_);
  and (_10373_, _10372_, _05758_);
  or (_10374_, _05541_, _03838_);
  nor (_10375_, _09611_, _04646_);
  and (_10376_, _04646_, \oc8051_golden_model_1.PSW [7]);
  nor (_10377_, _10376_, _10375_);
  nor (_10378_, _10377_, _04325_);
  and (_10379_, _03868_, _03838_);
  or (_10380_, _05361_, _03872_);
  nor (_10381_, _02603_, _02247_);
  and (_10382_, _02603_, \oc8051_golden_model_1.ACC [0]);
  nor (_10383_, _10382_, _10381_);
  and (_10384_, _10383_, _05361_);
  nor (_10385_, _10384_, _03843_);
  and (_10386_, _10385_, _10380_);
  nor (_10387_, _05085_, _03844_);
  or (_10388_, _10387_, _10386_);
  and (_10389_, _10388_, _05346_);
  nand (_10390_, _09977_, _09588_);
  and (_10391_, _10390_, _02886_);
  or (_10392_, _10391_, _04225_);
  or (_10393_, _10392_, _10389_);
  nor (_10394_, _02597_, \oc8051_golden_model_1.PC [0]);
  nor (_10395_, _10394_, _03868_);
  and (_10396_, _10395_, _10393_);
  or (_10397_, _10396_, _10379_);
  and (_10398_, _10397_, _05305_);
  nor (_10399_, _09977_, _04646_);
  and (_10400_, _10399_, _02879_);
  or (_10401_, _10400_, _02876_);
  or (_10402_, _10401_, _10398_);
  nand (_10403_, _07607_, _02876_);
  and (_10404_, _10403_, _02874_);
  and (_10405_, _10404_, _10402_);
  nor (_10406_, _09978_, _02874_);
  and (_10407_, _10406_, _10390_);
  or (_10408_, _10407_, _10405_);
  and (_10409_, _10408_, _02591_);
  or (_10410_, _02591_, _02247_);
  nand (_10411_, _02971_, _10410_);
  or (_10412_, _10411_, _10409_);
  nand (_10413_, _07607_, _03433_);
  and (_10414_, _10413_, _10412_);
  or (_10415_, _10414_, _03889_);
  or (_10416_, _05945_, _02838_);
  nand (_10417_, _10416_, _07606_);
  or (_10418_, _10417_, _05379_);
  and (_10419_, _10418_, _04325_);
  and (_10420_, _10419_, _10415_);
  or (_10421_, _10420_, _10378_);
  and (_10422_, _10421_, _04134_);
  and (_10423_, _02569_, \oc8051_golden_model_1.PC [0]);
  or (_10424_, _05536_, _10423_);
  or (_10425_, _10424_, _10422_);
  and (_10426_, _10425_, _10374_);
  or (_10427_, _10426_, _05540_);
  or (_10428_, _06164_, _05545_);
  and (_10429_, _10428_, _04193_);
  and (_10430_, _10429_, _10427_);
  and (_10431_, _05302_, _03838_);
  and (_10432_, _05673_, \oc8051_golden_model_1.ACC [0]);
  and (_10433_, _05676_, \oc8051_golden_model_1.B [0]);
  nor (_10434_, _10433_, _10432_);
  and (_10435_, _05681_, \oc8051_golden_model_1.P0INREG [0]);
  and (_10436_, _05663_, \oc8051_golden_model_1.SBUF [0]);
  nor (_10437_, _10436_, _10435_);
  and (_10438_, _10437_, _10434_);
  and (_10439_, _05657_, \oc8051_golden_model_1.SCON [0]);
  and (_10440_, _05667_, \oc8051_golden_model_1.PSW [0]);
  nor (_10441_, _10440_, _10439_);
  and (_10442_, _05683_, \oc8051_golden_model_1.TCON [0]);
  and (_10443_, _05652_, \oc8051_golden_model_1.P1INREG [0]);
  nor (_10444_, _10443_, _10442_);
  and (_10445_, _10444_, _10441_);
  and (_10446_, _10445_, _10438_);
  and (_10447_, _05694_, \oc8051_golden_model_1.PCON [0]);
  and (_10448_, _05691_, \oc8051_golden_model_1.DPH [0]);
  nor (_10449_, _10448_, _10447_);
  and (_10450_, _10449_, _10446_);
  and (_10451_, _05711_, \oc8051_golden_model_1.DPL [0]);
  and (_10452_, _05715_, \oc8051_golden_model_1.TL1 [0]);
  nor (_10453_, _10452_, _10451_);
  and (_10454_, _05700_, \oc8051_golden_model_1.TH0 [0]);
  and (_10455_, _05720_, \oc8051_golden_model_1.TMOD [0]);
  nor (_10456_, _10455_, _10454_);
  and (_10457_, _10456_, _10453_);
  and (_10458_, _05717_, \oc8051_golden_model_1.TH1 [0]);
  not (_10459_, _10458_);
  and (_10460_, _05730_, \oc8051_golden_model_1.IE [0]);
  and (_10461_, _05732_, \oc8051_golden_model_1.IP [0]);
  nor (_10462_, _10461_, _10460_);
  and (_10463_, _05724_, \oc8051_golden_model_1.P2INREG [0]);
  and (_10464_, _05727_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_10465_, _10464_, _10463_);
  and (_10466_, _10465_, _10462_);
  and (_10467_, _10466_, _10459_);
  and (_10468_, _05709_, \oc8051_golden_model_1.SP [0]);
  and (_10469_, _05705_, \oc8051_golden_model_1.TL0 [0]);
  nor (_10470_, _10469_, _10468_);
  and (_10471_, _10470_, _10467_);
  and (_10472_, _10471_, _10457_);
  and (_10473_, _10472_, _10450_);
  not (_10474_, _10473_);
  nor (_10475_, _10474_, _10431_);
  nor (_10476_, _10475_, _04193_);
  or (_10477_, _10476_, _05749_);
  or (_10478_, _10477_, _10430_);
  and (_10479_, _05749_, _02837_);
  nor (_10480_, _10479_, _02835_);
  and (_10481_, _10480_, _10478_);
  and (_10482_, _05660_, _02835_);
  or (_10483_, _10482_, _02522_);
  or (_10484_, _10483_, _10481_);
  and (_10485_, _02522_, _02247_);
  nor (_10486_, _10485_, _05758_);
  and (_10487_, _10486_, _10484_);
  or (_10488_, _10487_, _10373_);
  and (_10489_, _10488_, _05769_);
  or (_10490_, _10489_, _10370_);
  and (_10491_, _10490_, _05768_);
  and (_10492_, _10371_, _05271_);
  or (_10493_, _10492_, _10491_);
  and (_10494_, _10493_, _04129_);
  and (_10495_, _10368_, _03909_);
  or (_10496_, _10495_, _02530_);
  or (_10497_, _10496_, _10494_);
  and (_10498_, _02530_, _02247_);
  nor (_10499_, _10498_, _05781_);
  and (_10500_, _10499_, _10497_);
  or (_10501_, _10500_, _10366_);
  and (_10502_, _10501_, _10364_);
  nor (_10503_, _10367_, _10364_);
  or (_10504_, _10503_, _02528_);
  or (_10505_, _10504_, _10502_);
  nand (_10506_, _02528_, _02247_);
  and (_10507_, _10506_, _09723_);
  and (_10508_, _10507_, _10505_);
  or (_10509_, _03927_, _03872_);
  and (_10510_, _10509_, _09725_);
  or (_10511_, _10510_, _10508_);
  or (_10512_, _05945_, _05809_);
  and (_10513_, _10512_, _10511_);
  or (_10514_, _10513_, _03929_);
  nand (_10515_, _05085_, _03929_);
  and (_10516_, _10515_, _06185_);
  and (_10517_, _10516_, _10514_);
  and (_10518_, _03034_, _02247_);
  or (_10519_, _10518_, _02505_);
  or (_10520_, _10519_, _10517_);
  and (_10521_, _10520_, _10363_);
  or (_10522_, _10521_, _02801_);
  or (_10523_, _10375_, _02802_);
  and (_10524_, _10523_, _05257_);
  and (_10525_, _10524_, _10522_);
  and (_10526_, _06154_, _03872_);
  or (_10527_, _10526_, _10525_);
  and (_10528_, _10527_, _06161_);
  and (_10529_, _05945_, _03941_);
  or (_10530_, _10529_, _03943_);
  or (_10531_, _10530_, _10528_);
  nand (_10532_, _05085_, _03943_);
  and (_10533_, _10532_, _04562_);
  and (_10534_, _10533_, _10531_);
  or (_10535_, _10534_, _10362_);
  and (_10536_, _04555_, _04548_);
  nor (_10537_, _10536_, _04556_);
  and (_10538_, _04555_, _03955_);
  and (_10539_, _10538_, _10537_);
  nor (_10540_, _10361_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_10541_, _10540_, _10539_);
  and (_10542_, _10541_, _10535_);
  nand (_10543_, _08921_, _03034_);
  or (_10544_, _09097_, _03034_);
  and (_10545_, _10544_, _10543_);
  and (_10546_, _10545_, _04555_);
  and (_10547_, _10546_, _10539_);
  or (_35855_, _10547_, _10542_);
  nor (_10548_, _04554_, _04128_);
  not (_10549_, _10548_);
  not (_10550_, _03955_);
  and (_10551_, _10548_, _04548_);
  and (_10552_, _10548_, _04551_);
  or (_10553_, _10552_, _10551_);
  or (_10554_, _10553_, _10550_);
  or (_10556_, _10554_, _10549_);
  or (_10557_, _10361_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_10558_, _10557_, _10556_);
  nor (_10559_, _05352_, _05250_);
  and (_10560_, _10559_, _06154_);
  not (_10561_, _10559_);
  or (_10562_, _10561_, _09722_);
  nor (_10563_, _05037_, _02543_);
  and (_10564_, _05037_, _02543_);
  nor (_10565_, _10564_, _10563_);
  and (_10567_, _10565_, _05762_);
  not (_10568_, _09950_);
  nand (_10569_, _09949_, _09533_);
  and (_10570_, _10569_, _02873_);
  and (_10571_, _10570_, _10568_);
  nor (_10572_, _09949_, _04637_);
  or (_10573_, _10572_, _05305_);
  nor (_10574_, _05467_, _05086_);
  nor (_10575_, _10574_, _03844_);
  nand (_10576_, _10559_, _09132_);
  nor (_10578_, _02603_, \oc8051_golden_model_1.PC [1]);
  and (_10579_, _02603_, \oc8051_golden_model_1.ACC [1]);
  nor (_10580_, _10579_, _10578_);
  and (_10581_, _10580_, _05361_);
  nor (_10582_, _10581_, _03843_);
  and (_10583_, _10582_, _10576_);
  or (_10584_, _10583_, _02886_);
  or (_10585_, _10584_, _10575_);
  or (_10586_, _10569_, _05346_);
  and (_10587_, _10586_, _10585_);
  or (_10589_, _10587_, _04225_);
  nor (_10590_, _02597_, _02220_);
  nor (_10591_, _10590_, _03868_);
  and (_10592_, _10591_, _10589_);
  and (_10593_, _04021_, _03868_);
  or (_10594_, _10593_, _02879_);
  or (_10595_, _10594_, _10592_);
  and (_10596_, _10595_, _10573_);
  or (_10597_, _10596_, _02876_);
  nand (_10598_, _07595_, _02876_);
  and (_10600_, _10598_, _02874_);
  and (_10601_, _10600_, _10597_);
  or (_10602_, _10601_, _10571_);
  and (_10603_, _10602_, _02591_);
  or (_10604_, _02591_, \oc8051_golden_model_1.PC [1]);
  nand (_10605_, _02971_, _10604_);
  or (_10606_, _10605_, _10603_);
  nand (_10607_, _07595_, _03433_);
  and (_10608_, _10607_, _10606_);
  or (_10609_, _10608_, _03889_);
  or (_10611_, _05900_, _02838_);
  nand (_10612_, _10611_, _07594_);
  or (_10613_, _10612_, _05379_);
  and (_10614_, _10613_, _04325_);
  and (_10615_, _10614_, _10609_);
  nor (_10616_, _09556_, _04637_);
  and (_10617_, _04637_, \oc8051_golden_model_1.PSW [7]);
  nor (_10618_, _10617_, _10616_);
  nor (_10619_, _10618_, _04325_);
  or (_10620_, _10619_, _02569_);
  or (_10622_, _10620_, _10615_);
  and (_10623_, _02569_, \oc8051_golden_model_1.PC [1]);
  nor (_10624_, _10623_, _05536_);
  and (_10625_, _10624_, _10622_);
  nor (_10626_, _04020_, _05541_);
  or (_10627_, _10626_, _05540_);
  or (_10628_, _10627_, _10625_);
  or (_10629_, _06163_, _05545_);
  and (_10630_, _10629_, _04193_);
  and (_10631_, _10630_, _10628_);
  nor (_10632_, _05549_, _04020_);
  and (_10633_, _05663_, \oc8051_golden_model_1.SBUF [1]);
  and (_10634_, _05667_, \oc8051_golden_model_1.PSW [1]);
  or (_10635_, _10634_, _10633_);
  and (_10636_, _05683_, \oc8051_golden_model_1.TCON [1]);
  and (_10637_, _05673_, \oc8051_golden_model_1.ACC [1]);
  or (_10638_, _10637_, _10636_);
  or (_10639_, _10638_, _10635_);
  and (_10640_, _05657_, \oc8051_golden_model_1.SCON [1]);
  and (_10641_, _05676_, \oc8051_golden_model_1.B [1]);
  or (_10642_, _10641_, _10640_);
  and (_10643_, _05681_, \oc8051_golden_model_1.P0INREG [1]);
  and (_10644_, _05652_, \oc8051_golden_model_1.P1INREG [1]);
  or (_10645_, _10644_, _10643_);
  or (_10646_, _10645_, _10642_);
  or (_10647_, _10646_, _10639_);
  and (_10648_, _05691_, \oc8051_golden_model_1.DPH [1]);
  and (_10649_, _05694_, \oc8051_golden_model_1.PCON [1]);
  or (_10650_, _10649_, _10648_);
  or (_10651_, _10650_, _10647_);
  and (_10652_, _05715_, \oc8051_golden_model_1.TL1 [1]);
  and (_10653_, _05705_, \oc8051_golden_model_1.TL0 [1]);
  or (_10654_, _10653_, _10652_);
  and (_10655_, _05711_, \oc8051_golden_model_1.DPL [1]);
  and (_10656_, _05720_, \oc8051_golden_model_1.TMOD [1]);
  or (_10657_, _10656_, _10655_);
  or (_10658_, _10657_, _10654_);
  and (_10659_, _05717_, \oc8051_golden_model_1.TH1 [1]);
  and (_10660_, _05724_, \oc8051_golden_model_1.P2INREG [1]);
  and (_10661_, _05732_, \oc8051_golden_model_1.IP [1]);
  or (_10662_, _10661_, _10660_);
  and (_10663_, _05730_, \oc8051_golden_model_1.IE [1]);
  and (_10664_, _05727_, \oc8051_golden_model_1.P3INREG [1]);
  or (_10665_, _10664_, _10663_);
  or (_10666_, _10665_, _10662_);
  or (_10667_, _10666_, _10659_);
  and (_10668_, _05709_, \oc8051_golden_model_1.SP [1]);
  and (_10669_, _05700_, \oc8051_golden_model_1.TH0 [1]);
  or (_10670_, _10669_, _10668_);
  or (_10671_, _10670_, _10667_);
  or (_10672_, _10671_, _10658_);
  or (_10673_, _10672_, _10651_);
  or (_10674_, _10673_, _10632_);
  and (_10675_, _10674_, _04192_);
  or (_10676_, _10675_, _05749_);
  or (_10677_, _10676_, _10631_);
  and (_10678_, _05749_, _03687_);
  nor (_10679_, _10678_, _02835_);
  and (_10680_, _10679_, _10677_);
  and (_10681_, _05703_, _02835_);
  or (_10682_, _10681_, _02522_);
  or (_10683_, _10682_, _10680_);
  and (_10684_, _02522_, \oc8051_golden_model_1.PC [1]);
  nor (_10685_, _10684_, _05758_);
  and (_10686_, _10685_, _10683_);
  and (_10687_, _05037_, _03720_);
  nor (_10688_, _05037_, _03720_);
  nor (_10689_, _10688_, _10687_);
  and (_10690_, _10689_, _05758_);
  or (_10691_, _10690_, _10686_);
  and (_10692_, _10691_, _05769_);
  or (_10693_, _10692_, _10567_);
  and (_10694_, _10693_, _05768_);
  and (_10695_, _10688_, _05271_);
  or (_10696_, _10695_, _10694_);
  and (_10697_, _10696_, _04129_);
  and (_10698_, _10563_, _03909_);
  or (_10699_, _10698_, _02530_);
  or (_10700_, _10699_, _10697_);
  and (_10701_, _02530_, \oc8051_golden_model_1.PC [1]);
  nor (_10702_, _10701_, _05781_);
  and (_10703_, _10702_, _10700_);
  nor (_10704_, _10687_, _05786_);
  or (_10705_, _10704_, _05785_);
  or (_10706_, _10705_, _10703_);
  nand (_10707_, _10564_, _05785_);
  and (_10708_, _10707_, _05790_);
  and (_10709_, _10708_, _10706_);
  nand (_10710_, _02528_, _02220_);
  nand (_10711_, _09722_, _10710_);
  or (_10712_, _10711_, _10709_);
  nand (_10713_, _10712_, _10562_);
  nand (_10714_, _10713_, _04105_);
  and (_10715_, _03014_, _02504_);
  not (_10716_, _10715_);
  or (_10717_, _10561_, _04105_);
  and (_10718_, _10717_, _10716_);
  and (_10719_, _10718_, _10714_);
  or (_10720_, _06165_, _05946_);
  and (_10721_, _10720_, _10715_);
  or (_10722_, _10721_, _03589_);
  or (_10723_, _10722_, _10719_);
  or (_10724_, _10720_, _03590_);
  and (_10725_, _10724_, _05808_);
  and (_10726_, _10725_, _10723_);
  nor (_10727_, _10574_, _05808_);
  or (_10728_, _10727_, _03034_);
  or (_10729_, _10728_, _10726_);
  nand (_10730_, _03034_, _08894_);
  and (_10731_, _10730_, _09742_);
  and (_10732_, _10731_, _10729_);
  and (_10733_, _02505_, _02220_);
  or (_10734_, _02801_, _10733_);
  or (_10735_, _10734_, _10732_);
  or (_10736_, _10616_, _02802_);
  and (_10737_, _10736_, _05257_);
  and (_10738_, _10737_, _10735_);
  or (_10739_, _10738_, _10560_);
  nor (_10740_, _04139_, _03604_);
  and (_10741_, _10740_, _10739_);
  nor (_10742_, _06165_, _05946_);
  not (_10743_, _10740_);
  and (_10744_, _10743_, _10742_);
  or (_10745_, _10744_, _03943_);
  or (_10746_, _10745_, _10741_);
  or (_10747_, _10574_, _06160_);
  and (_10748_, _10747_, _04562_);
  and (_10749_, _10748_, _10746_);
  or (_10750_, _10749_, _10362_);
  and (_10751_, _10750_, _10558_);
  nand (_10752_, _08859_, _03034_);
  or (_10753_, _09043_, _03034_);
  and (_10754_, _10753_, _10752_);
  and (_10755_, _10754_, _04555_);
  and (_10756_, _10755_, _10539_);
  or (_35856_, _10756_, _10751_);
  nor (_10757_, _06165_, _06167_);
  nor (_10758_, _10757_, _07355_);
  or (_10759_, _10758_, _10740_);
  and (_10760_, _05946_, _06036_);
  nor (_10761_, _05946_, _06036_);
  or (_10762_, _10761_, _10760_);
  and (_10763_, _10762_, _03927_);
  nor (_10764_, _05134_, _06964_);
  and (_10765_, _05134_, _06964_);
  nor (_10766_, _10765_, _10764_);
  and (_10767_, _10766_, _05762_);
  and (_10768_, _05134_, _03262_);
  nor (_10769_, _05134_, _03262_);
  nor (_10770_, _10769_, _10768_);
  and (_10771_, _10770_, _05758_);
  nand (_10772_, _04449_, _05536_);
  nor (_10773_, _09938_, _04642_);
  or (_10774_, _10773_, _05305_);
  and (_10775_, _05352_, _04449_);
  nor (_10776_, _05352_, _04449_);
  or (_10777_, _10776_, _10775_);
  or (_10778_, _10777_, _05361_);
  nor (_10779_, _02620_, _02603_);
  and (_10780_, _02603_, \oc8051_golden_model_1.ACC [2]);
  nor (_10781_, _10780_, _10779_);
  nand (_10782_, _10781_, _05361_);
  and (_10783_, _10782_, _10778_);
  and (_10784_, _10783_, _03844_);
  and (_10785_, _05134_, _05037_);
  and (_10786_, _10785_, _05466_);
  nor (_10787_, _05467_, _05134_);
  nor (_10788_, _10787_, _10786_);
  nor (_10789_, _10788_, _03844_);
  or (_10790_, _10789_, _10784_);
  or (_10791_, _10790_, _02886_);
  nand (_10792_, _09938_, _09508_);
  or (_10793_, _10792_, _05346_);
  and (_10794_, _10793_, _10791_);
  or (_10795_, _10794_, _04225_);
  nor (_10796_, _02614_, _02597_);
  nor (_10797_, _10796_, _03868_);
  and (_10798_, _10797_, _10795_);
  and (_10799_, _04450_, _03868_);
  or (_10800_, _10799_, _02879_);
  or (_10801_, _10800_, _10798_);
  and (_10802_, _10801_, _10774_);
  or (_10803_, _10802_, _02876_);
  nand (_10804_, _07577_, _02876_);
  and (_10805_, _10804_, _02874_);
  and (_10806_, _10805_, _10803_);
  not (_10807_, _09939_);
  and (_10808_, _10792_, _10807_);
  and (_10809_, _10808_, _02873_);
  or (_10810_, _10809_, _10806_);
  and (_10811_, _10810_, _02591_);
  or (_10812_, _02620_, _02591_);
  nand (_10813_, _02971_, _10812_);
  or (_10814_, _10813_, _10811_);
  nand (_10815_, _07577_, _03433_);
  and (_10816_, _10815_, _10814_);
  or (_10817_, _10816_, _03889_);
  and (_10818_, _06167_, _02763_);
  nand (_10819_, _07576_, _03889_);
  or (_10820_, _10819_, _10818_);
  and (_10821_, _10820_, _10817_);
  or (_10822_, _10821_, _03888_);
  nor (_10823_, _09531_, _04642_);
  and (_10824_, _04642_, \oc8051_golden_model_1.PSW [7]);
  nor (_10825_, _10824_, _10823_);
  nand (_10826_, _10825_, _03888_);
  and (_10827_, _10826_, _04134_);
  and (_10828_, _10827_, _10822_);
  and (_10829_, _02614_, _02569_);
  or (_10830_, _05536_, _10829_);
  or (_10831_, _10830_, _10828_);
  and (_10832_, _10831_, _10772_);
  or (_10833_, _10832_, _05540_);
  or (_10834_, _06167_, _05545_);
  and (_10835_, _10834_, _04193_);
  and (_10836_, _10835_, _10833_);
  nor (_10837_, _05549_, _04449_);
  not (_10838_, _10837_);
  and (_10839_, _05667_, \oc8051_golden_model_1.PSW [2]);
  and (_10840_, _05673_, \oc8051_golden_model_1.ACC [2]);
  nor (_10841_, _10840_, _10839_);
  and (_10842_, _05681_, \oc8051_golden_model_1.P0INREG [2]);
  and (_10843_, _05676_, \oc8051_golden_model_1.B [2]);
  nor (_10844_, _10843_, _10842_);
  and (_10845_, _10844_, _10841_);
  and (_10846_, _05657_, \oc8051_golden_model_1.SCON [2]);
  and (_10847_, _05663_, \oc8051_golden_model_1.SBUF [2]);
  nor (_10848_, _10847_, _10846_);
  and (_10849_, _05683_, \oc8051_golden_model_1.TCON [2]);
  and (_10850_, _05652_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_10851_, _10850_, _10849_);
  and (_10852_, _10851_, _10848_);
  and (_10853_, _10852_, _10845_);
  and (_10854_, _05691_, \oc8051_golden_model_1.DPH [2]);
  and (_10855_, _05694_, \oc8051_golden_model_1.PCON [2]);
  nor (_10856_, _10855_, _10854_);
  and (_10857_, _10856_, _10853_);
  and (_10858_, _05720_, \oc8051_golden_model_1.TMOD [2]);
  and (_10859_, _05705_, \oc8051_golden_model_1.TL0 [2]);
  nor (_10860_, _10859_, _10858_);
  and (_10861_, _05700_, \oc8051_golden_model_1.TH0 [2]);
  and (_10862_, _05715_, \oc8051_golden_model_1.TL1 [2]);
  nor (_10863_, _10862_, _10861_);
  and (_10864_, _10863_, _10860_);
  and (_10865_, _05709_, \oc8051_golden_model_1.SP [2]);
  not (_10866_, _10865_);
  and (_10867_, _05724_, \oc8051_golden_model_1.P2INREG [2]);
  and (_10868_, _05732_, \oc8051_golden_model_1.IP [2]);
  nor (_10869_, _10868_, _10867_);
  and (_10870_, _05730_, \oc8051_golden_model_1.IE [2]);
  and (_10871_, _05727_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_10872_, _10871_, _10870_);
  and (_10873_, _10872_, _10869_);
  and (_10874_, _10873_, _10866_);
  and (_10875_, _05711_, \oc8051_golden_model_1.DPL [2]);
  and (_10876_, _05717_, \oc8051_golden_model_1.TH1 [2]);
  nor (_10877_, _10876_, _10875_);
  and (_10878_, _10877_, _10874_);
  and (_10879_, _10878_, _10864_);
  and (_10880_, _10879_, _10857_);
  and (_10881_, _10880_, _10838_);
  nor (_10882_, _10881_, _04193_);
  or (_10883_, _10882_, _05749_);
  or (_10884_, _10883_, _10836_);
  and (_10885_, _05749_, _03356_);
  nor (_10886_, _10885_, _02835_);
  and (_10887_, _10886_, _10884_);
  and (_10888_, _05693_, _02835_);
  or (_10889_, _10888_, _02522_);
  or (_10890_, _10889_, _10887_);
  and (_10891_, _02620_, _02522_);
  nor (_10892_, _10891_, _05758_);
  and (_10893_, _10892_, _10890_);
  or (_10894_, _10893_, _10771_);
  and (_10895_, _10894_, _05769_);
  or (_10896_, _10895_, _10767_);
  and (_10897_, _10896_, _05768_);
  and (_10898_, _10769_, _05271_);
  or (_10899_, _10898_, _10897_);
  and (_10900_, _10899_, _04129_);
  and (_10901_, _10764_, _03909_);
  or (_10902_, _10901_, _02530_);
  or (_10903_, _10902_, _10900_);
  and (_10904_, _02620_, _02530_);
  nor (_10905_, _10904_, _05781_);
  and (_10906_, _10905_, _10903_);
  nor (_10907_, _10768_, _05786_);
  or (_10908_, _10907_, _05785_);
  or (_10909_, _10908_, _10906_);
  nand (_10910_, _10765_, _05785_);
  and (_10911_, _10910_, _05790_);
  and (_10912_, _10911_, _10909_);
  nand (_10913_, _02614_, _02528_);
  nand (_10914_, _09723_, _10913_);
  or (_10915_, _10914_, _10912_);
  or (_10916_, _10777_, _09723_);
  and (_10917_, _10916_, _05809_);
  and (_10918_, _10917_, _10915_);
  or (_10919_, _10918_, _10763_);
  and (_10920_, _10919_, _05808_);
  nor (_10921_, _10788_, _05808_);
  or (_10922_, _10921_, _03034_);
  or (_10923_, _10922_, _10920_);
  nand (_10924_, _08892_, _03034_);
  and (_10925_, _10924_, _09742_);
  and (_10926_, _10925_, _10923_);
  and (_10927_, _02614_, _02505_);
  or (_10928_, _02801_, _10927_);
  or (_10929_, _10928_, _10926_);
  or (_10930_, _10823_, _02802_);
  and (_10931_, _10930_, _05257_);
  and (_10932_, _10931_, _10929_);
  or (_10933_, _05250_, _04450_);
  nor (_10934_, _05257_, _07267_);
  and (_10935_, _10934_, _10933_);
  or (_10936_, _10935_, _10743_);
  or (_10937_, _10936_, _10932_);
  and (_10938_, _10937_, _10759_);
  or (_10939_, _10938_, _03943_);
  nor (_10940_, _05135_, _05086_);
  nor (_10941_, _10940_, _05136_);
  or (_10942_, _10941_, _06160_);
  and (_10943_, _10942_, _04562_);
  and (_10944_, _10943_, _10939_);
  or (_10945_, _10944_, _10362_);
  nor (_10946_, _10361_, \oc8051_golden_model_1.IRAM[0] [2]);
  nor (_10947_, _10946_, _10539_);
  and (_10948_, _10947_, _10945_);
  nand (_10949_, _08852_, _03034_);
  or (_10950_, _09036_, _03034_);
  and (_10951_, _10950_, _10949_);
  and (_10952_, _10951_, _04555_);
  and (_10953_, _10952_, _10539_);
  or (_35857_, _10953_, _10948_);
  or (_10954_, _10361_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_10955_, _10954_, _10556_);
  or (_10956_, _07267_, _07266_);
  nor (_10957_, _05257_, _05252_);
  and (_10958_, _10957_, _10956_);
  nor (_10959_, _10760_, _05991_);
  or (_10960_, _10959_, _06038_);
  and (_10961_, _10960_, _03927_);
  and (_10962_, _04992_, _02625_);
  nor (_10963_, _04992_, _02625_);
  nor (_10964_, _10963_, _10962_);
  and (_10965_, _10964_, _05762_);
  nor (_10966_, _04992_, _03128_);
  and (_10967_, _04992_, _03128_);
  nor (_10968_, _10967_, _10966_);
  and (_10969_, _10968_, _05758_);
  nand (_10970_, _04275_, _05536_);
  and (_10971_, _04695_, \oc8051_golden_model_1.PSW [7]);
  nor (_10972_, _09663_, _04695_);
  nor (_10973_, _10972_, _10971_);
  nor (_10974_, _10973_, _04325_);
  not (_10975_, _10003_);
  nand (_10976_, _10002_, _09640_);
  and (_10977_, _10976_, _02873_);
  and (_10978_, _10977_, _10975_);
  nor (_10979_, _10002_, _04695_);
  or (_10980_, _10979_, _05305_);
  or (_10981_, _10976_, _05346_);
  nor (_10982_, _10786_, _04992_);
  nor (_10983_, _10982_, _05469_);
  nor (_10984_, _10983_, _03844_);
  nor (_10985_, _10775_, _04275_);
  or (_10986_, _10985_, _05354_);
  or (_10987_, _10986_, _05361_);
  nor (_10988_, _02661_, _02603_);
  and (_10989_, _02603_, \oc8051_golden_model_1.ACC [3]);
  nor (_10990_, _10989_, _10988_);
  and (_10991_, _10990_, _05361_);
  nor (_10992_, _10991_, _03843_);
  and (_10993_, _10992_, _10987_);
  or (_10994_, _10993_, _02886_);
  or (_10995_, _10994_, _10984_);
  and (_10996_, _10995_, _10981_);
  or (_10997_, _10996_, _04225_);
  nor (_10998_, _02640_, _02597_);
  nor (_10999_, _10998_, _03868_);
  and (_11000_, _10999_, _10997_);
  and (_11001_, _07266_, _03868_);
  or (_11002_, _11001_, _02879_);
  or (_11003_, _11002_, _11000_);
  and (_11004_, _11003_, _10980_);
  or (_11005_, _11004_, _02876_);
  nand (_11006_, _07566_, _02876_);
  and (_11007_, _11006_, _02874_);
  and (_11008_, _11007_, _11005_);
  or (_11009_, _11008_, _10978_);
  and (_11010_, _11009_, _02591_);
  or (_11011_, _02661_, _02591_);
  nand (_11012_, _02971_, _11011_);
  or (_11013_, _11012_, _11010_);
  nand (_11014_, _07566_, _03433_);
  and (_11015_, _11014_, _11013_);
  or (_11016_, _11015_, _03889_);
  and (_11017_, _06166_, _02763_);
  nand (_11018_, _07565_, _03889_);
  or (_11019_, _11018_, _11017_);
  and (_11020_, _11019_, _04325_);
  and (_11021_, _11020_, _11016_);
  or (_11022_, _11021_, _10974_);
  and (_11023_, _11022_, _04134_);
  and (_11024_, _02640_, _02569_);
  or (_11025_, _05536_, _11024_);
  or (_11026_, _11025_, _11023_);
  and (_11027_, _11026_, _10970_);
  or (_11028_, _11027_, _05540_);
  or (_11029_, _06166_, _05545_);
  and (_11030_, _11029_, _04193_);
  and (_11031_, _11030_, _11028_);
  nor (_11032_, _05549_, _04275_);
  and (_11033_, _05681_, \oc8051_golden_model_1.P0INREG [3]);
  and (_11034_, _05652_, \oc8051_golden_model_1.P1INREG [3]);
  nor (_11035_, _11034_, _11033_);
  and (_11036_, _05657_, \oc8051_golden_model_1.SCON [3]);
  and (_11037_, _05667_, \oc8051_golden_model_1.PSW [3]);
  nor (_11038_, _11037_, _11036_);
  and (_11039_, _11038_, _11035_);
  and (_11040_, _05683_, \oc8051_golden_model_1.TCON [3]);
  and (_11041_, _05673_, \oc8051_golden_model_1.ACC [3]);
  nor (_11042_, _11041_, _11040_);
  and (_11043_, _05663_, \oc8051_golden_model_1.SBUF [3]);
  and (_11044_, _05676_, \oc8051_golden_model_1.B [3]);
  nor (_11045_, _11044_, _11043_);
  and (_11046_, _11045_, _11042_);
  and (_11047_, _11046_, _11039_);
  and (_11048_, _05691_, \oc8051_golden_model_1.DPH [3]);
  and (_11049_, _05694_, \oc8051_golden_model_1.PCON [3]);
  nor (_11050_, _11049_, _11048_);
  and (_11051_, _11050_, _11047_);
  and (_11052_, _05711_, \oc8051_golden_model_1.DPL [3]);
  and (_11053_, _05720_, \oc8051_golden_model_1.TMOD [3]);
  nor (_11054_, _11053_, _11052_);
  and (_11055_, _05705_, \oc8051_golden_model_1.TL0 [3]);
  and (_11056_, _05717_, \oc8051_golden_model_1.TH1 [3]);
  nor (_11057_, _11056_, _11055_);
  and (_11058_, _11057_, _11054_);
  and (_11059_, _05709_, \oc8051_golden_model_1.SP [3]);
  not (_11060_, _11059_);
  and (_11061_, _05724_, \oc8051_golden_model_1.P2INREG [3]);
  and (_11062_, _05732_, \oc8051_golden_model_1.IP [3]);
  nor (_11063_, _11062_, _11061_);
  and (_11064_, _05730_, \oc8051_golden_model_1.IE [3]);
  and (_11065_, _05727_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_11066_, _11065_, _11064_);
  and (_11067_, _11066_, _11063_);
  and (_11068_, _11067_, _11060_);
  and (_11069_, _05700_, \oc8051_golden_model_1.TH0 [3]);
  and (_11070_, _05715_, \oc8051_golden_model_1.TL1 [3]);
  nor (_11071_, _11070_, _11069_);
  and (_11072_, _11071_, _11068_);
  and (_11073_, _11072_, _11058_);
  and (_11074_, _11073_, _11051_);
  not (_11075_, _11074_);
  nor (_11076_, _11075_, _11032_);
  nor (_11077_, _11076_, _04193_);
  or (_11078_, _11077_, _05749_);
  or (_11079_, _11078_, _11031_);
  nor (_11080_, _05748_, _02794_);
  nor (_11081_, _11080_, _02835_);
  and (_11082_, _11081_, _11079_);
  and (_11083_, _05654_, _02835_);
  or (_11084_, _11083_, _02522_);
  or (_11085_, _11084_, _11082_);
  and (_11086_, _02661_, _02522_);
  nor (_11087_, _11086_, _05758_);
  and (_11088_, _11087_, _11085_);
  or (_11089_, _11088_, _10969_);
  and (_11090_, _11089_, _05769_);
  or (_11091_, _11090_, _10965_);
  and (_11092_, _11091_, _05768_);
  and (_11093_, _10966_, _05271_);
  or (_11094_, _11093_, _11092_);
  and (_11095_, _11094_, _04129_);
  and (_11096_, _10963_, _03909_);
  or (_11097_, _11096_, _02530_);
  or (_11098_, _11097_, _11095_);
  and (_11099_, _02661_, _02530_);
  nor (_11100_, _11099_, _05781_);
  and (_11101_, _11100_, _11098_);
  nor (_11102_, _10967_, _05786_);
  or (_11103_, _11102_, _05785_);
  or (_11104_, _11103_, _11101_);
  nand (_11105_, _10962_, _05785_);
  and (_11106_, _11105_, _05790_);
  and (_11107_, _11106_, _11104_);
  nand (_11108_, _02640_, _02528_);
  nand (_11109_, _09723_, _11108_);
  or (_11110_, _11109_, _11107_);
  or (_11111_, _10986_, _09723_);
  and (_11112_, _11111_, _05809_);
  and (_11113_, _11112_, _11110_);
  or (_11114_, _11113_, _10961_);
  and (_11115_, _11114_, _05808_);
  nor (_11116_, _10983_, _05808_);
  or (_11117_, _11116_, _03034_);
  or (_11118_, _11117_, _11115_);
  nand (_11119_, _08887_, _03034_);
  and (_11120_, _11119_, _09742_);
  and (_11121_, _11120_, _11118_);
  and (_11122_, _02640_, _02505_);
  or (_11123_, _02801_, _11122_);
  or (_11124_, _11123_, _11121_);
  or (_11125_, _10972_, _02802_);
  and (_11126_, _11125_, _05257_);
  and (_11127_, _11126_, _11124_);
  or (_11128_, _11127_, _10958_);
  and (_11129_, _11128_, _06161_);
  or (_11130_, _07355_, _06166_);
  nor (_11131_, _06169_, _06161_);
  and (_11132_, _11131_, _11130_);
  or (_11133_, _11132_, _03943_);
  or (_11134_, _11133_, _11129_);
  nor (_11135_, _05136_, _04993_);
  nor (_11136_, _11135_, _05137_);
  or (_11137_, _11136_, _06160_);
  and (_11138_, _11137_, _04562_);
  and (_11139_, _11138_, _11134_);
  or (_11140_, _11139_, _10362_);
  and (_11141_, _11140_, _10955_);
  nand (_11142_, _08845_, _03034_);
  or (_11143_, _09030_, _03034_);
  and (_11144_, _11143_, _11142_);
  and (_11145_, _11144_, _04555_);
  and (_11146_, _11145_, _10539_);
  or (_35858_, _11146_, _11141_);
  or (_11147_, _10361_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_11148_, _11147_, _10556_);
  or (_11149_, _05252_, _05249_);
  nor (_11150_, _05257_, _05253_);
  and (_11151_, _11150_, _11149_);
  and (_11152_, _05239_, _06864_);
  nor (_11153_, _05239_, _06864_);
  nor (_11154_, _11153_, _11152_);
  and (_11155_, _11154_, _05762_);
  nor (_11156_, _05617_, _05239_);
  and (_11157_, _05617_, _05239_);
  nor (_11158_, _11157_, _11156_);
  and (_11159_, _11158_, _05758_);
  nand (_11160_, _05192_, _05536_);
  nor (_11161_, _09583_, _09559_);
  and (_11162_, _09559_, \oc8051_golden_model_1.PSW [7]);
  nor (_11163_, _11162_, _11161_);
  nor (_11164_, _11163_, _04325_);
  nor (_11165_, _09559_, _09963_);
  or (_11166_, _11165_, _05305_);
  nand (_11167_, _09560_, _09963_);
  or (_11168_, _11167_, _05346_);
  nor (_11169_, _05354_, _05192_);
  and (_11170_, _05354_, _05192_);
  or (_11171_, _11170_, _11169_);
  or (_11172_, _11171_, _05361_);
  and (_11173_, _02603_, \oc8051_golden_model_1.ACC [4]);
  nor (_11174_, _09067_, _02603_);
  nor (_11175_, _11174_, _11173_);
  nand (_11176_, _11175_, _05361_);
  and (_11177_, _11176_, _11172_);
  or (_11178_, _11177_, _03840_);
  or (_11179_, _06171_, _05371_);
  and (_11180_, _11179_, _11178_);
  or (_11181_, _11180_, _03843_);
  and (_11182_, _05469_, _05239_);
  nor (_11183_, _05469_, _05239_);
  nor (_11184_, _11183_, _11182_);
  nand (_11185_, _11184_, _03843_);
  and (_11186_, _11185_, _11181_);
  or (_11187_, _11186_, _02886_);
  and (_11188_, _11187_, _11168_);
  or (_11189_, _11188_, _04225_);
  nor (_11190_, _09066_, _02597_);
  nor (_11191_, _11190_, _03868_);
  and (_11192_, _11191_, _11189_);
  and (_11193_, _05249_, _03868_);
  or (_11194_, _11193_, _02879_);
  or (_11195_, _11194_, _11192_);
  and (_11196_, _11195_, _11166_);
  or (_11197_, _11196_, _02876_);
  nand (_11198_, _07638_, _02876_);
  and (_11199_, _11198_, _02874_);
  and (_11200_, _11199_, _11197_);
  not (_11201_, _09964_);
  and (_11202_, _11167_, _11201_);
  and (_11203_, _11202_, _02873_);
  or (_11204_, _11203_, _11200_);
  and (_11205_, _11204_, _02591_);
  or (_11206_, _09067_, _02591_);
  nand (_11207_, _11206_, _02971_);
  or (_11208_, _11207_, _11205_);
  nand (_11209_, _07638_, _03433_);
  and (_11210_, _11209_, _11208_);
  or (_11211_, _11210_, _03889_);
  and (_11212_, _06171_, _02763_);
  nand (_11213_, _07637_, _03889_);
  or (_11214_, _11213_, _11212_);
  and (_11215_, _11214_, _04325_);
  and (_11216_, _11215_, _11211_);
  or (_11217_, _11216_, _11164_);
  and (_11218_, _11217_, _04134_);
  and (_11219_, _09066_, _02569_);
  or (_11220_, _11219_, _05536_);
  or (_11221_, _11220_, _11218_);
  and (_11222_, _11221_, _11160_);
  or (_11223_, _11222_, _05540_);
  or (_11224_, _06171_, _05545_);
  and (_11225_, _11224_, _04193_);
  and (_11226_, _11225_, _11223_);
  nor (_11227_, _05549_, _05192_);
  not (_11228_, _11227_);
  and (_11229_, _05652_, \oc8051_golden_model_1.P1INREG [4]);
  and (_11230_, _05657_, \oc8051_golden_model_1.SCON [4]);
  nor (_11231_, _11230_, _11229_);
  and (_11232_, _05681_, \oc8051_golden_model_1.P0INREG [4]);
  and (_11233_, _05673_, \oc8051_golden_model_1.ACC [4]);
  nor (_11234_, _11233_, _11232_);
  and (_11235_, _11234_, _11231_);
  and (_11236_, _05663_, \oc8051_golden_model_1.SBUF [4]);
  and (_11237_, _05676_, \oc8051_golden_model_1.B [4]);
  nor (_11238_, _11237_, _11236_);
  and (_11239_, _05683_, \oc8051_golden_model_1.TCON [4]);
  and (_11240_, _05667_, \oc8051_golden_model_1.PSW [4]);
  nor (_11241_, _11240_, _11239_);
  and (_11242_, _11241_, _11238_);
  and (_11243_, _11242_, _11235_);
  and (_11244_, _05694_, \oc8051_golden_model_1.PCON [4]);
  and (_11245_, _05691_, \oc8051_golden_model_1.DPH [4]);
  nor (_11246_, _11245_, _11244_);
  and (_11247_, _11246_, _11243_);
  and (_11248_, _05711_, \oc8051_golden_model_1.DPL [4]);
  and (_11249_, _05705_, \oc8051_golden_model_1.TL0 [4]);
  nor (_11250_, _11249_, _11248_);
  and (_11251_, _05700_, \oc8051_golden_model_1.TH0 [4]);
  and (_11252_, _05717_, \oc8051_golden_model_1.TH1 [4]);
  nor (_11253_, _11252_, _11251_);
  and (_11254_, _11253_, _11250_);
  and (_11255_, _05709_, \oc8051_golden_model_1.SP [4]);
  not (_11256_, _11255_);
  and (_11257_, _05724_, \oc8051_golden_model_1.P2INREG [4]);
  and (_11258_, _05732_, \oc8051_golden_model_1.IP [4]);
  nor (_11259_, _11258_, _11257_);
  and (_11260_, _05730_, \oc8051_golden_model_1.IE [4]);
  and (_11261_, _05727_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_11262_, _11261_, _11260_);
  and (_11263_, _11262_, _11259_);
  and (_11264_, _11263_, _11256_);
  and (_11265_, _05715_, \oc8051_golden_model_1.TL1 [4]);
  and (_11266_, _05720_, \oc8051_golden_model_1.TMOD [4]);
  nor (_11267_, _11266_, _11265_);
  and (_11268_, _11267_, _11264_);
  and (_11269_, _11268_, _11254_);
  and (_11270_, _11269_, _11247_);
  and (_11271_, _11270_, _11228_);
  nor (_11272_, _11271_, _04193_);
  or (_11273_, _11272_, _05749_);
  or (_11274_, _11273_, _11226_);
  and (_11275_, _05749_, _03647_);
  nor (_11276_, _11275_, _02835_);
  and (_11277_, _11276_, _11274_);
  and (_11278_, _05618_, _02835_);
  or (_11279_, _11278_, _02522_);
  or (_11280_, _11279_, _11277_);
  and (_11281_, _09067_, _02522_);
  nor (_11282_, _11281_, _05758_);
  and (_11283_, _11282_, _11280_);
  or (_11284_, _11283_, _11159_);
  and (_11285_, _11284_, _05769_);
  or (_11286_, _11285_, _11155_);
  and (_11287_, _11286_, _05768_);
  and (_11288_, _11156_, _05271_);
  or (_11289_, _11288_, _11287_);
  and (_11290_, _11289_, _04129_);
  and (_11291_, _11153_, _03909_);
  or (_11292_, _11291_, _02530_);
  or (_11293_, _11292_, _11290_);
  and (_11294_, _09067_, _02530_);
  nor (_11295_, _11294_, _05781_);
  and (_11296_, _11295_, _11293_);
  nor (_11297_, _11157_, _05786_);
  or (_11298_, _11297_, _05785_);
  or (_11299_, _11298_, _11296_);
  nand (_11300_, _11152_, _05785_);
  and (_11301_, _11300_, _05790_);
  and (_11302_, _11301_, _11299_);
  nand (_11303_, _09066_, _02528_);
  nand (_11304_, _11303_, _09723_);
  or (_11305_, _11304_, _11302_);
  or (_11306_, _11171_, _09723_);
  and (_11307_, _11306_, _10716_);
  and (_11308_, _11307_, _11305_);
  and (_11309_, _06038_, _06128_);
  nor (_11310_, _06038_, _06128_);
  or (_11311_, _11310_, _11309_);
  or (_11312_, _11311_, _03589_);
  and (_11313_, _11312_, _03927_);
  or (_11314_, _11313_, _11308_);
  or (_11315_, _11311_, _03590_);
  and (_11316_, _11315_, _05808_);
  and (_11317_, _11316_, _11314_);
  nor (_11318_, _11184_, _05808_);
  or (_11319_, _11318_, _03034_);
  or (_11320_, _11319_, _11317_);
  nand (_11321_, _08883_, _03034_);
  and (_11322_, _11321_, _09742_);
  and (_11323_, _11322_, _11320_);
  and (_11324_, _09066_, _02505_);
  or (_11325_, _11324_, _02801_);
  or (_11326_, _11325_, _11323_);
  or (_11327_, _11161_, _02802_);
  and (_11328_, _11327_, _05257_);
  and (_11329_, _11328_, _11326_);
  or (_11330_, _11329_, _11151_);
  and (_11331_, _11330_, _10740_);
  or (_11332_, _06169_, _06171_);
  nor (_11333_, _10740_, _07337_);
  and (_11334_, _11333_, _11332_);
  or (_11335_, _11334_, _03943_);
  or (_11336_, _11335_, _11331_);
  nor (_11337_, _05240_, _05137_);
  nor (_11338_, _11337_, _05241_);
  or (_11339_, _11338_, _06160_);
  and (_11340_, _11339_, _04562_);
  and (_11341_, _11340_, _11336_);
  or (_11342_, _11341_, _10362_);
  and (_11343_, _11342_, _11148_);
  nand (_11344_, _08841_, _03034_);
  or (_11345_, _09026_, _03034_);
  and (_11346_, _11345_, _11344_);
  and (_11347_, _11346_, _04555_);
  and (_11348_, _11347_, _10539_);
  or (_35859_, _11348_, _11343_);
  or (_11349_, _10361_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_11350_, _11349_, _10556_);
  nor (_11351_, _05253_, _05248_);
  nor (_11352_, _11351_, _05254_);
  and (_11353_, _11352_, _06154_);
  nor (_11354_, _04944_, _06858_);
  and (_11355_, _04944_, _06858_);
  nor (_11356_, _11355_, _11354_);
  and (_11357_, _11356_, _05762_);
  nand (_11358_, _04894_, _05536_);
  nor (_11359_, _09688_, _09665_);
  and (_11360_, _09665_, \oc8051_golden_model_1.PSW [7]);
  nor (_11361_, _11360_, _11359_);
  nor (_11362_, _11361_, _04325_);
  nor (_11363_, _09665_, _10014_);
  or (_11364_, _11363_, _05305_);
  nand (_11365_, _09666_, _10014_);
  or (_11366_, _11365_, _05346_);
  or (_11367_, _06170_, _05371_);
  nor (_11368_, _11170_, _04894_);
  or (_11369_, _11368_, _05355_);
  and (_11370_, _11369_, _09132_);
  and (_11371_, _02603_, \oc8051_golden_model_1.ACC [5]);
  nor (_11372_, _09062_, _02603_);
  or (_11373_, _11372_, _11371_);
  and (_11374_, _11373_, _05361_);
  or (_11375_, _11374_, _03840_);
  or (_11376_, _11375_, _11370_);
  and (_11377_, _11376_, _11367_);
  or (_11378_, _11377_, _03843_);
  nor (_11379_, _11182_, _04944_);
  nor (_11380_, _11379_, _05470_);
  nand (_11381_, _11380_, _03843_);
  and (_11382_, _11381_, _11378_);
  or (_11383_, _11382_, _02886_);
  and (_11384_, _11383_, _11366_);
  or (_11385_, _11384_, _04225_);
  nor (_11386_, _09061_, _02597_);
  nor (_11387_, _11386_, _03868_);
  and (_11388_, _11387_, _11385_);
  and (_11389_, _05248_, _03868_);
  or (_11390_, _11389_, _02879_);
  or (_11391_, _11390_, _11388_);
  and (_11392_, _11391_, _11364_);
  or (_11393_, _11392_, _02876_);
  nand (_11394_, _07621_, _02876_);
  and (_11395_, _11394_, _02874_);
  and (_11396_, _11395_, _11393_);
  not (_11397_, _10015_);
  and (_11398_, _11365_, _11397_);
  and (_11399_, _11398_, _02873_);
  or (_11400_, _11399_, _11396_);
  and (_11401_, _11400_, _02591_);
  or (_11402_, _09062_, _02591_);
  nand (_11403_, _11402_, _02971_);
  or (_11404_, _11403_, _11401_);
  nand (_11405_, _07621_, _03433_);
  and (_11406_, _11405_, _11404_);
  or (_11407_, _11406_, _03889_);
  and (_11408_, _06170_, _02763_);
  nand (_11409_, _07620_, _03889_);
  or (_11410_, _11409_, _11408_);
  and (_11411_, _11410_, _04325_);
  and (_11412_, _11411_, _11407_);
  or (_11413_, _11412_, _11362_);
  and (_11414_, _11413_, _04134_);
  and (_11415_, _09061_, _02569_);
  or (_11416_, _11415_, _05536_);
  or (_11417_, _11416_, _11414_);
  and (_11418_, _11417_, _11358_);
  or (_11419_, _11418_, _05540_);
  or (_11420_, _06170_, _05545_);
  and (_11421_, _11420_, _04193_);
  and (_11422_, _11421_, _11419_);
  nor (_11423_, _05549_, _04894_);
  not (_11424_, _11423_);
  and (_11425_, _05667_, \oc8051_golden_model_1.PSW [5]);
  and (_11426_, _05673_, \oc8051_golden_model_1.ACC [5]);
  nor (_11427_, _11426_, _11425_);
  and (_11428_, _05681_, \oc8051_golden_model_1.P0INREG [5]);
  and (_11429_, _05657_, \oc8051_golden_model_1.SCON [5]);
  nor (_11430_, _11429_, _11428_);
  and (_11431_, _11430_, _11427_);
  and (_11432_, _05663_, \oc8051_golden_model_1.SBUF [5]);
  and (_11433_, _05676_, \oc8051_golden_model_1.B [5]);
  nor (_11434_, _11433_, _11432_);
  and (_11435_, _05683_, \oc8051_golden_model_1.TCON [5]);
  and (_11436_, _05652_, \oc8051_golden_model_1.P1INREG [5]);
  nor (_11437_, _11436_, _11435_);
  and (_11438_, _11437_, _11434_);
  and (_11439_, _11438_, _11431_);
  and (_11440_, _05694_, \oc8051_golden_model_1.PCON [5]);
  and (_11441_, _05691_, \oc8051_golden_model_1.DPH [5]);
  nor (_11442_, _11441_, _11440_);
  and (_11443_, _11442_, _11439_);
  and (_11444_, _05711_, \oc8051_golden_model_1.DPL [5]);
  and (_11445_, _05715_, \oc8051_golden_model_1.TL1 [5]);
  nor (_11446_, _11445_, _11444_);
  and (_11447_, _05705_, \oc8051_golden_model_1.TL0 [5]);
  and (_11448_, _05717_, \oc8051_golden_model_1.TH1 [5]);
  nor (_11449_, _11448_, _11447_);
  and (_11450_, _11449_, _11446_);
  and (_11451_, _05700_, \oc8051_golden_model_1.TH0 [5]);
  not (_11452_, _11451_);
  and (_11453_, _05724_, \oc8051_golden_model_1.P2INREG [5]);
  and (_11454_, _05727_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_11455_, _11454_, _11453_);
  and (_11456_, _05730_, \oc8051_golden_model_1.IE [5]);
  and (_11457_, _05732_, \oc8051_golden_model_1.IP [5]);
  nor (_11458_, _11457_, _11456_);
  and (_11459_, _11458_, _11455_);
  and (_11460_, _11459_, _11452_);
  and (_11461_, _05709_, \oc8051_golden_model_1.SP [5]);
  and (_11462_, _05720_, \oc8051_golden_model_1.TMOD [5]);
  nor (_11463_, _11462_, _11461_);
  and (_11464_, _11463_, _11460_);
  and (_11465_, _11464_, _11450_);
  and (_11466_, _11465_, _11443_);
  and (_11467_, _11466_, _11424_);
  nor (_11468_, _11467_, _04193_);
  or (_11469_, _11468_, _05749_);
  or (_11470_, _11469_, _11422_);
  and (_11471_, _05749_, _03220_);
  nor (_11472_, _11471_, _02835_);
  and (_11473_, _11472_, _11470_);
  and (_11474_, _05671_, _02835_);
  or (_11475_, _11474_, _02522_);
  or (_11476_, _11475_, _11473_);
  and (_11477_, _09062_, _02522_);
  nor (_11478_, _11477_, _05758_);
  and (_11479_, _11478_, _11476_);
  and (_11480_, _05649_, _04944_);
  nor (_11481_, _05649_, _04944_);
  nor (_11482_, _11481_, _11480_);
  and (_11483_, _11482_, _05758_);
  or (_11484_, _11483_, _11479_);
  and (_11485_, _11484_, _05769_);
  or (_11486_, _11485_, _11357_);
  and (_11487_, _11486_, _05768_);
  and (_11488_, _11481_, _05271_);
  or (_11489_, _11488_, _11487_);
  and (_11490_, _11489_, _04129_);
  and (_11491_, _11354_, _03909_);
  or (_11492_, _11491_, _02530_);
  or (_11493_, _11492_, _11490_);
  and (_11494_, _09062_, _02530_);
  nor (_11495_, _11494_, _05781_);
  and (_11496_, _11495_, _11493_);
  nor (_11497_, _11480_, _05786_);
  or (_11498_, _11497_, _05785_);
  or (_11499_, _11498_, _11496_);
  nand (_11500_, _11355_, _05785_);
  and (_11501_, _11500_, _05790_);
  and (_11502_, _11501_, _11499_);
  and (_11503_, _05797_, _09721_);
  nand (_11504_, _09061_, _02528_);
  nand (_11505_, _11504_, _11503_);
  or (_11506_, _11505_, _11502_);
  and (_11507_, _11369_, _05801_);
  or (_11508_, _11507_, _09723_);
  and (_11509_, _11508_, _11506_);
  and (_11510_, _11369_, _03587_);
  or (_11511_, _11510_, _10715_);
  or (_11512_, _11511_, _11509_);
  nor (_11513_, _11309_, _06083_);
  or (_11514_, _11513_, _06130_);
  or (_11515_, _11514_, _10716_);
  and (_11516_, _11515_, _11512_);
  and (_11517_, _11516_, _03590_);
  and (_11518_, _11514_, _03589_);
  or (_11519_, _11518_, _11517_);
  and (_11520_, _11519_, _05808_);
  nor (_11521_, _11380_, _05808_);
  or (_11522_, _11521_, _03034_);
  or (_11523_, _11522_, _11520_);
  nand (_11524_, _08878_, _03034_);
  and (_11525_, _11524_, _09742_);
  and (_11526_, _11525_, _11523_);
  and (_11527_, _09061_, _02505_);
  or (_11528_, _11527_, _02801_);
  or (_11529_, _11528_, _11526_);
  or (_11530_, _11359_, _02802_);
  and (_11531_, _11530_, _05257_);
  and (_11532_, _11531_, _11529_);
  or (_11533_, _11532_, _11353_);
  and (_11534_, _11533_, _06161_);
  or (_11535_, _07337_, _06170_);
  nor (_11536_, _06173_, _06161_);
  and (_11537_, _11536_, _11535_);
  or (_11538_, _11537_, _03943_);
  or (_11539_, _11538_, _11534_);
  nor (_11540_, _05241_, _04945_);
  nor (_11541_, _11540_, _05242_);
  or (_11542_, _11541_, _06160_);
  and (_11543_, _11542_, _04562_);
  and (_11544_, _11543_, _11539_);
  or (_11545_, _11544_, _10362_);
  and (_11546_, _11545_, _11350_);
  nor (_11547_, _09022_, _03034_);
  and (_11548_, _08834_, _03034_);
  or (_11549_, _11548_, _11547_);
  and (_11550_, _11549_, _04555_);
  and (_11551_, _11550_, _10539_);
  or (_35860_, _11551_, _11546_);
  or (_11552_, _10361_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_11553_, _11552_, _10556_);
  nor (_11554_, _04837_, _06807_);
  and (_11555_, _04837_, _06807_);
  nor (_11556_, _11555_, _11554_);
  and (_11557_, _11556_, _05762_);
  and (_11558_, _05585_, _04837_);
  nor (_11559_, _05585_, _04837_);
  nor (_11560_, _11559_, _11558_);
  and (_11561_, _11560_, _05758_);
  nor (_11562_, _09613_, _09989_);
  or (_11563_, _11562_, _05305_);
  nand (_11564_, _09614_, _09989_);
  or (_11565_, _11564_, _05346_);
  nor (_11566_, _05470_, _04837_);
  nor (_11567_, _11566_, _05471_);
  nand (_11568_, _11567_, _03843_);
  or (_11569_, _06162_, _05371_);
  and (_11570_, _05361_, _05371_);
  and (_11571_, _02603_, \oc8051_golden_model_1.ACC [6]);
  nor (_11572_, _09055_, _02603_);
  nor (_11573_, _11572_, _11571_);
  nand (_11574_, _11573_, _11570_);
  nor (_11575_, _05355_, _04790_);
  or (_11576_, _11575_, _05356_);
  or (_11577_, _11576_, _05361_);
  and (_11578_, _11577_, _11574_);
  and (_11579_, _11578_, _11569_);
  or (_11580_, _11579_, _03843_);
  and (_11581_, _11580_, _11568_);
  or (_11582_, _11581_, _02886_);
  and (_11583_, _11582_, _11565_);
  or (_11584_, _11583_, _04225_);
  nor (_11585_, _09054_, _02597_);
  nor (_11586_, _11585_, _03868_);
  and (_11587_, _11586_, _11584_);
  and (_11588_, _07235_, _03868_);
  or (_11589_, _11588_, _02879_);
  or (_11590_, _11589_, _11587_);
  and (_11591_, _11590_, _11563_);
  or (_11592_, _11591_, _02876_);
  nand (_11593_, _07552_, _02876_);
  and (_11594_, _11593_, _02874_);
  and (_11595_, _11594_, _11592_);
  not (_11596_, _09990_);
  and (_11597_, _11564_, _11596_);
  and (_11598_, _11597_, _02873_);
  or (_11599_, _11598_, _11595_);
  and (_11600_, _11599_, _02591_);
  or (_11601_, _09055_, _02591_);
  nand (_11602_, _11601_, _02971_);
  or (_11603_, _11602_, _11600_);
  nand (_11604_, _07552_, _03433_);
  and (_11605_, _11604_, _11603_);
  or (_11606_, _11605_, _03889_);
  and (_11607_, _06162_, _02763_);
  nand (_11608_, _07551_, _03889_);
  or (_11609_, _11608_, _11607_);
  and (_11610_, _11609_, _04325_);
  and (_11611_, _11610_, _11606_);
  nor (_11612_, _09637_, _09613_);
  and (_11613_, _09613_, \oc8051_golden_model_1.PSW [7]);
  nor (_11614_, _11613_, _11612_);
  nor (_11615_, _11614_, _04325_);
  or (_11616_, _11615_, _02569_);
  or (_11617_, _11616_, _11611_);
  and (_11618_, _09055_, _02569_);
  nor (_11619_, _11618_, _05536_);
  and (_11620_, _11619_, _11617_);
  nor (_11621_, _04790_, _05541_);
  or (_11622_, _11621_, _05540_);
  or (_11623_, _11622_, _11620_);
  or (_11624_, _06162_, _05545_);
  and (_11625_, _11624_, _04193_);
  and (_11626_, _11625_, _11623_);
  nor (_11627_, _05549_, _04790_);
  not (_11628_, _11627_);
  and (_11629_, _05681_, \oc8051_golden_model_1.P0INREG [6]);
  and (_11630_, _05676_, \oc8051_golden_model_1.B [6]);
  nor (_11631_, _11630_, _11629_);
  and (_11632_, _05683_, \oc8051_golden_model_1.TCON [6]);
  and (_11633_, _05667_, \oc8051_golden_model_1.PSW [6]);
  nor (_11634_, _11633_, _11632_);
  and (_11635_, _11634_, _11631_);
  and (_11636_, _05657_, \oc8051_golden_model_1.SCON [6]);
  and (_11637_, _05673_, \oc8051_golden_model_1.ACC [6]);
  nor (_11638_, _11637_, _11636_);
  and (_11639_, _05652_, \oc8051_golden_model_1.P1INREG [6]);
  and (_11640_, _05663_, \oc8051_golden_model_1.SBUF [6]);
  nor (_11641_, _11640_, _11639_);
  and (_11642_, _11641_, _11638_);
  and (_11643_, _11642_, _11635_);
  and (_11644_, _05691_, \oc8051_golden_model_1.DPH [6]);
  and (_11645_, _05694_, \oc8051_golden_model_1.PCON [6]);
  nor (_11646_, _11645_, _11644_);
  and (_11647_, _11646_, _11643_);
  and (_11648_, _05709_, \oc8051_golden_model_1.SP [6]);
  and (_11649_, _05720_, \oc8051_golden_model_1.TMOD [6]);
  nor (_11650_, _11649_, _11648_);
  and (_11651_, _05711_, \oc8051_golden_model_1.DPL [6]);
  and (_11652_, _05715_, \oc8051_golden_model_1.TL1 [6]);
  nor (_11653_, _11652_, _11651_);
  and (_11654_, _11653_, _11650_);
  and (_11655_, _05700_, \oc8051_golden_model_1.TH0 [6]);
  not (_11656_, _11655_);
  and (_11657_, _05724_, \oc8051_golden_model_1.P2INREG [6]);
  and (_11658_, _05727_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_11659_, _11658_, _11657_);
  and (_11660_, _05730_, \oc8051_golden_model_1.IE [6]);
  and (_11661_, _05732_, \oc8051_golden_model_1.IP [6]);
  nor (_11662_, _11661_, _11660_);
  and (_11663_, _11662_, _11659_);
  and (_11664_, _11663_, _11656_);
  and (_11665_, _05705_, \oc8051_golden_model_1.TL0 [6]);
  and (_11666_, _05717_, \oc8051_golden_model_1.TH1 [6]);
  nor (_11667_, _11666_, _11665_);
  and (_11668_, _11667_, _11664_);
  and (_11669_, _11668_, _11654_);
  and (_11670_, _11669_, _11647_);
  and (_11671_, _11670_, _11628_);
  nor (_11672_, _11671_, _04193_);
  or (_11673_, _11672_, _05749_);
  or (_11674_, _11673_, _11626_);
  and (_11675_, _05749_, _02924_);
  nor (_11676_, _11675_, _02835_);
  and (_11677_, _11676_, _11674_);
  not (_11678_, _05585_);
  and (_11679_, _11678_, _02835_);
  or (_11680_, _11679_, _02522_);
  or (_11681_, _11680_, _11677_);
  and (_11682_, _09055_, _02522_);
  nor (_11683_, _11682_, _05758_);
  and (_11684_, _11683_, _11681_);
  or (_11685_, _11684_, _11561_);
  and (_11686_, _11685_, _05769_);
  or (_11687_, _11686_, _11557_);
  and (_11688_, _11687_, _05768_);
  and (_11689_, _11559_, _05271_);
  or (_11690_, _11689_, _11688_);
  and (_11691_, _11690_, _04129_);
  and (_11692_, _11554_, _03909_);
  or (_11693_, _11692_, _02530_);
  or (_11694_, _11693_, _11691_);
  and (_11695_, _09055_, _02530_);
  nor (_11696_, _11695_, _05781_);
  and (_11697_, _11696_, _11694_);
  nor (_11698_, _11558_, _05786_);
  or (_11699_, _11698_, _05785_);
  or (_11700_, _11699_, _11697_);
  nand (_11701_, _11555_, _05785_);
  and (_11702_, _11701_, _05790_);
  and (_11703_, _11702_, _11700_);
  nand (_11704_, _09054_, _02528_);
  nand (_11705_, _11704_, _09723_);
  or (_11706_, _11705_, _11703_);
  or (_11707_, _11576_, _09723_);
  and (_11708_, _11707_, _10716_);
  and (_11709_, _11708_, _11706_);
  nor (_11710_, _06130_, _05855_);
  or (_11711_, _11710_, _06131_);
  or (_11712_, _11711_, _03589_);
  and (_11713_, _11712_, _03927_);
  or (_11714_, _11713_, _11709_);
  or (_11715_, _11711_, _03590_);
  and (_11716_, _11715_, _05808_);
  and (_11717_, _11716_, _11714_);
  nor (_11718_, _11567_, _05808_);
  or (_11719_, _11718_, _03034_);
  or (_11720_, _11719_, _11717_);
  nand (_11721_, _08869_, _03034_);
  and (_11722_, _11721_, _09742_);
  and (_11723_, _11722_, _11720_);
  and (_11724_, _09054_, _02505_);
  or (_11725_, _11724_, _02801_);
  or (_11726_, _11725_, _11723_);
  or (_11727_, _11612_, _02802_);
  and (_11728_, _11727_, _05257_);
  and (_11729_, _11728_, _11726_);
  or (_11730_, _05254_, _07235_);
  nor (_11731_, _07236_, _05257_);
  and (_11732_, _11731_, _11730_);
  or (_11733_, _11732_, _04139_);
  or (_11734_, _11733_, _11729_);
  nor (_11735_, _06173_, _06162_);
  nor (_11736_, _11735_, _06174_);
  nor (_11737_, _11736_, _04140_);
  nor (_11738_, _11737_, _03604_);
  and (_11739_, _11738_, _11734_);
  and (_11740_, _11736_, _03604_);
  or (_11741_, _11740_, _03943_);
  or (_11742_, _11741_, _11739_);
  nor (_11743_, _05242_, _04838_);
  nor (_11744_, _11743_, _05243_);
  or (_11745_, _11744_, _06160_);
  and (_11746_, _11745_, _04562_);
  and (_11747_, _11746_, _11742_);
  or (_11748_, _11747_, _10362_);
  and (_11749_, _11748_, _11553_);
  or (_11750_, _08826_, _06185_);
  or (_11751_, _09015_, _03034_);
  and (_11752_, _11751_, _11750_);
  and (_11753_, _11752_, _04555_);
  and (_11754_, _11753_, _10539_);
  or (_35861_, _11754_, _11749_);
  or (_11755_, _10361_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_11756_, _11755_, _10556_);
  or (_11757_, _10362_, _06182_);
  and (_11758_, _11757_, _11756_);
  and (_11759_, _10539_, _06209_);
  or (_35862_, _11759_, _11758_);
  and (_11760_, _04564_, _04127_);
  and (_11761_, _11760_, _10359_);
  or (_11762_, _11761_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_11763_, _04215_);
  or (_11764_, _10553_, _11763_);
  or (_11765_, _11764_, _10549_);
  and (_11766_, _11765_, _11762_);
  not (_11767_, _11761_);
  or (_11768_, _11767_, _10534_);
  and (_11769_, _11768_, _11766_);
  and (_11770_, _04555_, _04215_);
  and (_11771_, _11770_, _10537_);
  and (_11772_, _11771_, _10546_);
  or (_35911_, _11772_, _11769_);
  or (_11773_, _11761_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_11774_, _11773_, _11765_);
  or (_11775_, _11767_, _10749_);
  and (_11776_, _11775_, _11774_);
  and (_11777_, _11771_, _10755_);
  or (_35912_, _11777_, _11776_);
  or (_11778_, _11761_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_11779_, _11778_, _11765_);
  or (_11780_, _11767_, _10944_);
  and (_11781_, _11780_, _11779_);
  and (_11782_, _11771_, _10952_);
  or (_35913_, _11782_, _11781_);
  or (_11783_, _11761_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_11784_, _11783_, _11765_);
  or (_11785_, _11767_, _11139_);
  and (_11786_, _11785_, _11784_);
  and (_11787_, _11771_, _11145_);
  or (_35914_, _11787_, _11786_);
  or (_11788_, _11761_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_11789_, _11788_, _11765_);
  or (_11790_, _11767_, _11341_);
  and (_11791_, _11790_, _11789_);
  and (_11792_, _11771_, _11347_);
  or (_35915_, _11792_, _11791_);
  or (_11793_, _11761_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_11794_, _11793_, _11765_);
  or (_11795_, _11767_, _11544_);
  and (_11796_, _11795_, _11794_);
  and (_11797_, _11771_, _11550_);
  or (_35916_, _11797_, _11796_);
  or (_11798_, _11761_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_11799_, _11798_, _11765_);
  or (_11800_, _11767_, _11747_);
  and (_11801_, _11800_, _11799_);
  and (_11802_, _11771_, _11753_);
  or (_35917_, _11802_, _11801_);
  or (_11803_, _11761_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_11804_, _11803_, _11765_);
  or (_11805_, _11767_, _06182_);
  and (_11806_, _11805_, _11804_);
  and (_11807_, _11771_, _06209_);
  or (_35918_, _11807_, _11806_);
  nor (_11808_, _04384_, _04211_);
  nor (_11809_, _11808_, _04541_);
  and (_11810_, _04212_, _03949_);
  and (_11811_, _11810_, _11809_);
  or (_11812_, _11811_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_11813_, _05373_);
  or (_11814_, _10553_, _11813_);
  or (_11815_, _11814_, _10549_);
  and (_11816_, _11815_, _11812_);
  and (_11817_, _10532_, _04210_);
  and (_11818_, _11817_, _10531_);
  not (_11819_, _11811_);
  or (_11820_, _11819_, _11818_);
  and (_11821_, _11820_, _11816_);
  and (_11822_, _05373_, _04555_);
  and (_11823_, _11822_, _10537_);
  and (_11824_, _11823_, _10546_);
  or (_35919_, _11824_, _11821_);
  or (_11825_, _11811_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_11826_, _11825_, _11815_);
  not (_11827_, _10359_);
  nand (_11828_, _10356_, _03949_);
  or (_11829_, _11828_, _11827_);
  or (_11830_, _11829_, _10749_);
  and (_11831_, _11830_, _11826_);
  and (_11832_, _11823_, _10755_);
  or (_35920_, _11832_, _11831_);
  or (_11833_, _11811_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_11834_, _11833_, _11815_);
  or (_11835_, _11829_, _10944_);
  and (_11836_, _11835_, _11834_);
  and (_11837_, _11823_, _10952_);
  or (_35921_, _11837_, _11836_);
  or (_11838_, _11811_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_11839_, _11838_, _11815_);
  and (_11840_, _11137_, _04210_);
  and (_11841_, _11840_, _11134_);
  or (_11842_, _11819_, _11841_);
  and (_11843_, _11842_, _11839_);
  and (_11844_, _11823_, _11145_);
  or (_35922_, _11844_, _11843_);
  or (_11845_, _11811_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_11846_, _11845_, _11815_);
  and (_11847_, _11339_, _04210_);
  and (_11848_, _11847_, _11336_);
  or (_11849_, _11819_, _11848_);
  and (_11850_, _11849_, _11846_);
  and (_11851_, _11823_, _11347_);
  or (_35923_, _11851_, _11850_);
  or (_11852_, _11811_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_11853_, _11852_, _11815_);
  and (_11854_, _11542_, _04210_);
  and (_11855_, _11854_, _11539_);
  or (_11856_, _11819_, _11855_);
  and (_11857_, _11856_, _11853_);
  and (_11858_, _11823_, _11550_);
  or (_35924_, _11858_, _11857_);
  or (_11859_, _11811_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_11860_, _11859_, _11815_);
  and (_11861_, _11745_, _04210_);
  and (_11862_, _11861_, _11742_);
  or (_11863_, _11819_, _11862_);
  and (_11864_, _11863_, _11860_);
  and (_11865_, _11823_, _11753_);
  or (_35925_, _11865_, _11864_);
  or (_11866_, _11811_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_11867_, _11866_, _11815_);
  or (_11868_, _11829_, _06182_);
  and (_11869_, _11868_, _11867_);
  and (_11870_, _11823_, _06209_);
  or (_35926_, _11870_, _11869_);
  and (_11871_, _10359_, _04565_);
  or (_11872_, _11871_, \oc8051_golden_model_1.IRAM[3] [0]);
  not (_11873_, _03954_);
  or (_11874_, _10553_, _11873_);
  or (_11875_, _11874_, _10549_);
  and (_11876_, _11875_, _11872_);
  not (_11877_, _11871_);
  or (_11878_, _11877_, _10534_);
  and (_11879_, _11878_, _11876_);
  and (_11880_, _04555_, _03954_);
  and (_11881_, _11880_, _10537_);
  and (_11882_, _11881_, _10546_);
  or (_35927_, _11882_, _11879_);
  or (_11883_, _11871_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_11884_, _11883_, _11875_);
  or (_11885_, _11877_, _10749_);
  and (_11886_, _11885_, _11884_);
  and (_11887_, _11881_, _10755_);
  or (_35928_, _11887_, _11886_);
  or (_11888_, _11871_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_11889_, _11888_, _11875_);
  or (_11890_, _11877_, _10944_);
  and (_11891_, _11890_, _11889_);
  and (_11892_, _11881_, _10952_);
  or (_35929_, _11892_, _11891_);
  or (_11893_, _11871_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_11894_, _11893_, _11875_);
  or (_11895_, _11877_, _11139_);
  and (_11896_, _11895_, _11894_);
  and (_11897_, _11881_, _11145_);
  or (_35930_, _11897_, _11896_);
  or (_11898_, _11871_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_11899_, _11898_, _11875_);
  or (_11900_, _11877_, _11341_);
  and (_11901_, _11900_, _11899_);
  and (_11902_, _11881_, _11347_);
  or (_35931_, _11902_, _11901_);
  or (_11903_, _11871_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_11904_, _11903_, _11875_);
  or (_11905_, _11877_, _11544_);
  and (_11906_, _11905_, _11904_);
  and (_11907_, _11881_, _11550_);
  or (_35932_, _11907_, _11906_);
  or (_11908_, _11877_, _11747_);
  or (_11909_, _11871_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_11910_, _11909_, _11875_);
  and (_11911_, _11910_, _11908_);
  and (_11912_, _11881_, _11753_);
  or (_35933_, _11912_, _11911_);
  or (_11913_, _11871_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_11914_, _11913_, _11875_);
  or (_11915_, _11877_, _06182_);
  and (_11916_, _11915_, _11914_);
  and (_11917_, _11881_, _06209_);
  or (_35934_, _11917_, _11916_);
  and (_11918_, _10358_, _04384_);
  and (_11919_, _11918_, _10357_);
  not (_11920_, _11919_);
  or (_11921_, _11920_, _10534_);
  not (_11922_, _04551_);
  and (_11923_, _10536_, _11922_);
  and (_11924_, _11923_, _03955_);
  nor (_11925_, _11919_, \oc8051_golden_model_1.IRAM[4] [0]);
  nor (_11926_, _11925_, _11924_);
  and (_11927_, _11926_, _11921_);
  and (_11928_, _11924_, _10546_);
  or (_35935_, _11928_, _11927_);
  or (_11929_, _11920_, _10749_);
  nor (_11930_, _11919_, \oc8051_golden_model_1.IRAM[4] [1]);
  nor (_11931_, _11930_, _11924_);
  and (_11932_, _11931_, _11929_);
  and (_11933_, _11924_, _10755_);
  or (_35936_, _11933_, _11932_);
  and (_11934_, _10551_, _11922_);
  nand (_11935_, _11934_, _03955_);
  nor (_11936_, _04211_, _03949_);
  nor (_11937_, _11936_, _04212_);
  and (_11938_, _04541_, _04384_);
  and (_11939_, _11938_, _11937_);
  or (_11940_, _11939_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_11941_, _11940_, _11935_);
  or (_11942_, _11920_, _10944_);
  and (_11943_, _11942_, _11941_);
  and (_11944_, _11924_, _10952_);
  or (_35937_, _11944_, _11943_);
  or (_11945_, _11939_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_11946_, _11945_, _11935_);
  not (_11947_, _11939_);
  or (_11948_, _11947_, _11841_);
  and (_11949_, _11948_, _11946_);
  and (_11950_, _11924_, _11145_);
  or (_35938_, _11950_, _11949_);
  or (_11951_, _11939_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_11952_, _11951_, _11935_);
  or (_11953_, _11947_, _11848_);
  and (_11954_, _11953_, _11952_);
  and (_11955_, _11924_, _11347_);
  or (_35939_, _11955_, _11954_);
  or (_11956_, _11939_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_11957_, _11956_, _11935_);
  or (_11958_, _11947_, _11855_);
  and (_11959_, _11958_, _11957_);
  and (_11960_, _11924_, _11550_);
  or (_35940_, _11960_, _11959_);
  or (_11961_, _11939_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_11962_, _11961_, _11935_);
  or (_11963_, _11947_, _11862_);
  and (_11964_, _11963_, _11962_);
  and (_11965_, _11924_, _11753_);
  or (_35941_, _11965_, _11964_);
  or (_11966_, _11939_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_11967_, _11966_, _11935_);
  or (_11968_, _11920_, _06182_);
  and (_11969_, _11968_, _11967_);
  and (_11970_, _11924_, _06209_);
  or (_35942_, _11970_, _11969_);
  and (_11971_, _11918_, _11760_);
  or (_11972_, _11971_, \oc8051_golden_model_1.IRAM[5] [0]);
  nand (_11973_, _11934_, _04215_);
  and (_11974_, _11973_, _11972_);
  not (_11975_, _11971_);
  or (_11976_, _11975_, _10534_);
  and (_11977_, _11976_, _11974_);
  and (_11978_, _11923_, _04215_);
  and (_11979_, _11978_, _10546_);
  or (_35943_, _11979_, _11977_);
  or (_11980_, _11971_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_11981_, _11980_, _11973_);
  or (_11982_, _11975_, _10749_);
  and (_11983_, _11982_, _11981_);
  and (_11984_, _11978_, _10755_);
  or (_35944_, _11984_, _11983_);
  or (_11985_, _11971_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_11986_, _11985_, _11973_);
  or (_11987_, _11975_, _10944_);
  and (_11988_, _11987_, _11986_);
  and (_11989_, _11978_, _10952_);
  or (_35945_, _11989_, _11988_);
  or (_11990_, _11971_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_11991_, _11990_, _11973_);
  or (_11992_, _11975_, _11139_);
  and (_11993_, _11992_, _11991_);
  and (_11994_, _11978_, _11145_);
  or (_35946_, _11994_, _11993_);
  or (_11995_, _11971_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_11996_, _11995_, _11973_);
  or (_11997_, _11975_, _11341_);
  and (_11998_, _11997_, _11996_);
  and (_11999_, _11978_, _11347_);
  or (_35947_, _11999_, _11998_);
  or (_12000_, _11975_, _11544_);
  or (_12001_, _11971_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_12002_, _12001_, _11973_);
  and (_12003_, _12002_, _12000_);
  and (_12004_, _11978_, _11550_);
  or (_35948_, _12004_, _12003_);
  or (_12005_, _11971_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_12006_, _12005_, _11973_);
  or (_12007_, _11975_, _11747_);
  and (_12008_, _12007_, _12006_);
  and (_12009_, _11978_, _11753_);
  or (_35949_, _12009_, _12008_);
  or (_12010_, _11971_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_12011_, _12010_, _11973_);
  or (_12012_, _11975_, _06182_);
  and (_12013_, _12012_, _12011_);
  and (_12014_, _11978_, _06209_);
  or (_35950_, _12014_, _12013_);
  not (_12015_, _11918_);
  nor (_12016_, _12015_, _11828_);
  not (_12017_, _12016_);
  or (_12018_, _12017_, _10534_);
  and (_12019_, _11934_, _05373_);
  not (_12020_, _12019_);
  or (_12021_, _12016_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_12022_, _12021_, _12020_);
  and (_12023_, _12022_, _12018_);
  and (_12024_, _12019_, _10546_);
  or (_35951_, _12024_, _12023_);
  or (_12025_, _12017_, _10749_);
  or (_12026_, _12016_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_12027_, _12026_, _12020_);
  and (_12028_, _12027_, _12025_);
  and (_12029_, _12019_, _10755_);
  or (_35952_, _12029_, _12028_);
  and (_12030_, _11938_, _11810_);
  or (_12031_, _12030_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_12032_, _12031_, _12020_);
  or (_12033_, _12017_, _10944_);
  and (_12034_, _12033_, _12032_);
  and (_12035_, _12019_, _10952_);
  or (_35953_, _12035_, _12034_);
  or (_12036_, _12030_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_12037_, _12036_, _12020_);
  not (_12038_, _12030_);
  or (_12039_, _12038_, _11841_);
  and (_12040_, _12039_, _12037_);
  and (_12041_, _12019_, _11145_);
  or (_35954_, _12041_, _12040_);
  or (_12042_, _12030_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_12043_, _12042_, _12020_);
  or (_12044_, _12038_, _11848_);
  and (_12045_, _12044_, _12043_);
  and (_12046_, _12019_, _11347_);
  or (_35955_, _12046_, _12045_);
  or (_12047_, _12030_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_12048_, _12047_, _12020_);
  or (_12049_, _12038_, _11855_);
  and (_12050_, _12049_, _12048_);
  and (_12051_, _12019_, _11550_);
  or (_35956_, _12051_, _12050_);
  or (_12052_, _12030_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_12053_, _12052_, _12020_);
  or (_12054_, _12038_, _11862_);
  and (_12055_, _12054_, _12053_);
  and (_12056_, _12019_, _11753_);
  or (_35957_, _12056_, _12055_);
  or (_12057_, _12030_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_12058_, _12057_, _12020_);
  or (_12059_, _12017_, _06182_);
  and (_12060_, _12059_, _12058_);
  and (_12061_, _12019_, _06209_);
  or (_35958_, _12061_, _12060_);
  and (_12062_, _11918_, _04565_);
  not (_12063_, _12062_);
  or (_12064_, _12063_, _10534_);
  and (_12065_, _11923_, _03954_);
  nor (_12066_, _12062_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_12067_, _12066_, _12065_);
  and (_12068_, _12067_, _12064_);
  and (_12069_, _12065_, _10546_);
  or (_35959_, _12069_, _12068_);
  or (_12070_, _12063_, _10749_);
  nor (_12071_, _12062_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_12072_, _12071_, _12065_);
  and (_12073_, _12072_, _12070_);
  and (_12074_, _12065_, _10755_);
  or (_35960_, _12074_, _12073_);
  nand (_12075_, _11934_, _03954_);
  and (_12076_, _11938_, _04213_);
  or (_12077_, _12076_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_12078_, _12077_, _12075_);
  or (_12079_, _12063_, _10944_);
  and (_12080_, _12079_, _12078_);
  and (_12081_, _12065_, _10952_);
  or (_35961_, _12081_, _12080_);
  or (_12082_, _12076_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_12083_, _12082_, _12075_);
  not (_12084_, _12076_);
  or (_12085_, _12084_, _11841_);
  and (_12086_, _12085_, _12083_);
  and (_12087_, _12065_, _11145_);
  or (_35962_, _12087_, _12086_);
  or (_12088_, _12076_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_12089_, _12088_, _12075_);
  or (_12090_, _12084_, _11848_);
  and (_12091_, _12090_, _12089_);
  and (_12092_, _12065_, _11347_);
  or (_35963_, _12092_, _12091_);
  or (_12093_, _12076_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_12094_, _12093_, _12075_);
  or (_12095_, _12084_, _11855_);
  and (_12096_, _12095_, _12094_);
  and (_12097_, _12065_, _11550_);
  or (_35964_, _12097_, _12096_);
  or (_12098_, _12076_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_12099_, _12098_, _12075_);
  or (_12100_, _12084_, _11862_);
  and (_12101_, _12100_, _12099_);
  and (_12102_, _12065_, _11753_);
  or (_35965_, _12102_, _12101_);
  or (_12103_, _12076_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_12104_, _12103_, _12075_);
  or (_12105_, _12063_, _06182_);
  and (_12106_, _12105_, _12104_);
  and (_12107_, _12065_, _06209_);
  or (_35966_, _12107_, _12106_);
  and (_12108_, _04567_, _04540_);
  and (_12109_, _12108_, _10357_);
  not (_12110_, _12109_);
  or (_12111_, _12110_, _10534_);
  not (_12112_, _04548_);
  and (_12113_, _04556_, _12112_);
  and (_12114_, _12113_, _03955_);
  not (_12115_, _12114_);
  or (_12116_, _12109_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_12117_, _12116_, _12115_);
  and (_12118_, _12117_, _12111_);
  and (_12119_, _12114_, _10546_);
  or (_35967_, _12119_, _12118_);
  or (_12120_, _12110_, _10749_);
  or (_12121_, _12109_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_12122_, _12121_, _12115_);
  and (_12123_, _12122_, _12120_);
  and (_12124_, _12114_, _10755_);
  or (_35968_, _12124_, _12123_);
  or (_12125_, _12109_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_12126_, _12125_, _12115_);
  or (_12127_, _12110_, _10944_);
  and (_12128_, _12127_, _12126_);
  and (_12129_, _12114_, _10952_);
  or (_35969_, _12129_, _12128_);
  or (_12130_, _12109_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_12131_, _12130_, _12115_);
  or (_12132_, _12110_, _11139_);
  and (_12133_, _12132_, _12131_);
  and (_12134_, _12114_, _11145_);
  or (_35970_, _12134_, _12133_);
  or (_12135_, _12109_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_12136_, _12135_, _12115_);
  or (_12137_, _12110_, _11341_);
  and (_12138_, _12137_, _12136_);
  and (_12139_, _12114_, _11347_);
  or (_35971_, _12139_, _12138_);
  or (_12140_, _12109_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_12141_, _12140_, _12115_);
  or (_12142_, _12110_, _11544_);
  and (_12143_, _12142_, _12141_);
  and (_12144_, _12114_, _11550_);
  or (_35972_, _12144_, _12143_);
  or (_12145_, _12109_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_12146_, _12145_, _12115_);
  or (_12147_, _12110_, _11747_);
  and (_12148_, _12147_, _12146_);
  and (_12149_, _12114_, _11753_);
  or (_35973_, _12149_, _12148_);
  or (_12150_, _12109_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_12151_, _12150_, _12115_);
  or (_12152_, _12110_, _06182_);
  and (_12153_, _12152_, _12151_);
  and (_12154_, _12114_, _06209_);
  or (_35974_, _12154_, _12153_);
  and (_12155_, _12108_, _11760_);
  or (_12156_, _12155_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_12157_, _10552_, _04216_);
  and (_12158_, _12157_, _12156_);
  not (_12159_, _12155_);
  or (_12160_, _12159_, _10534_);
  and (_12161_, _12160_, _12158_);
  and (_12162_, _12113_, _04215_);
  and (_12163_, _12162_, _10546_);
  or (_35975_, _12163_, _12161_);
  or (_12164_, _12159_, _10749_);
  or (_12165_, _12155_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_12166_, _12165_, _12157_);
  and (_12167_, _12166_, _12164_);
  and (_12168_, _12162_, _10755_);
  or (_35976_, _12168_, _12167_);
  or (_12169_, _12159_, _10944_);
  or (_12170_, _12155_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_12171_, _12170_, _12157_);
  and (_12172_, _12171_, _12169_);
  and (_12173_, _12162_, _10952_);
  or (_35977_, _12173_, _12172_);
  or (_12174_, _12155_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_12175_, _12174_, _12157_);
  or (_12176_, _12159_, _11139_);
  and (_12177_, _12176_, _12175_);
  and (_12178_, _12162_, _11145_);
  or (_35978_, _12178_, _12177_);
  or (_12179_, _12155_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_12180_, _12179_, _12157_);
  or (_12181_, _12159_, _11341_);
  and (_12182_, _12181_, _12180_);
  and (_12183_, _12162_, _11347_);
  or (_35979_, _12183_, _12182_);
  or (_12184_, _12155_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_12185_, _12184_, _12157_);
  or (_12186_, _12159_, _11544_);
  and (_12187_, _12186_, _12185_);
  and (_12188_, _12162_, _11550_);
  or (_35980_, _12188_, _12187_);
  or (_12189_, _12155_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_12190_, _12189_, _12157_);
  or (_12191_, _12159_, _11747_);
  and (_12192_, _12191_, _12190_);
  and (_12193_, _12162_, _11753_);
  or (_35981_, _12193_, _12192_);
  or (_12194_, _12155_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_12195_, _12194_, _12157_);
  or (_12196_, _12159_, _06182_);
  and (_12197_, _12196_, _12195_);
  and (_12198_, _12162_, _06209_);
  or (_35982_, _12198_, _12197_);
  not (_12199_, _12108_);
  nor (_12200_, _12199_, _11828_);
  not (_12201_, _12200_);
  or (_12202_, _12201_, _10534_);
  and (_12203_, _12113_, _05373_);
  not (_12204_, _12203_);
  or (_12205_, _12200_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_12206_, _12205_, _12204_);
  and (_12207_, _12206_, _12202_);
  and (_12208_, _12203_, _10546_);
  or (_35863_, _12208_, _12207_);
  or (_12209_, _12201_, _10749_);
  or (_12210_, _12200_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_12211_, _12210_, _12204_);
  and (_12212_, _12211_, _12209_);
  and (_12213_, _12203_, _10755_);
  or (_35864_, _12213_, _12212_);
  and (_12214_, _11808_, _04540_);
  and (_12215_, _12214_, _11810_);
  or (_12216_, _12215_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_12217_, _12216_, _12204_);
  or (_12218_, _12201_, _10944_);
  and (_12219_, _12218_, _12217_);
  and (_12220_, _12203_, _10952_);
  or (_35865_, _12220_, _12219_);
  or (_12221_, _12215_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_12222_, _12221_, _12204_);
  or (_12223_, _12201_, _11139_);
  and (_12224_, _12223_, _12222_);
  and (_12225_, _12203_, _11145_);
  or (_35866_, _12225_, _12224_);
  or (_12226_, _12215_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_12227_, _12226_, _12204_);
  or (_12228_, _12201_, _11341_);
  and (_12229_, _12228_, _12227_);
  and (_12230_, _12203_, _11347_);
  or (_35867_, _12230_, _12229_);
  or (_12231_, _12215_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_12232_, _12231_, _12204_);
  or (_12233_, _12201_, _11544_);
  and (_12234_, _12233_, _12232_);
  and (_12235_, _12203_, _11550_);
  or (_35868_, _12235_, _12234_);
  or (_12236_, _12215_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_12237_, _12236_, _12204_);
  or (_12238_, _12201_, _11747_);
  and (_12239_, _12238_, _12237_);
  and (_12240_, _12203_, _11753_);
  or (_35869_, _12240_, _12239_);
  or (_12241_, _12215_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_12242_, _12241_, _12204_);
  or (_12243_, _12201_, _06182_);
  and (_12244_, _12243_, _12242_);
  and (_12245_, _12203_, _06209_);
  or (_35870_, _12245_, _12244_);
  and (_12246_, _12108_, _04565_);
  not (_12247_, _12246_);
  or (_12248_, _12247_, _10534_);
  and (_12249_, _12113_, _03954_);
  not (_12250_, _12249_);
  or (_12251_, _12246_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_12252_, _12251_, _12250_);
  and (_12253_, _12252_, _12248_);
  and (_12254_, _12249_, _10546_);
  or (_35871_, _12254_, _12253_);
  or (_12255_, _12247_, _10749_);
  or (_12256_, _12246_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_12257_, _12256_, _12250_);
  and (_12258_, _12257_, _12255_);
  and (_12259_, _12249_, _10755_);
  or (_35872_, _12259_, _12258_);
  or (_12260_, _12246_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_12261_, _12260_, _12250_);
  or (_12262_, _12247_, _10944_);
  and (_12263_, _12262_, _12261_);
  and (_12264_, _12249_, _10952_);
  or (_35873_, _12264_, _12263_);
  or (_12265_, _12246_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_12266_, _12265_, _12250_);
  or (_12267_, _12247_, _11139_);
  and (_12268_, _12267_, _12266_);
  and (_12269_, _12249_, _11145_);
  or (_35874_, _12269_, _12268_);
  or (_12270_, _12246_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_12271_, _12270_, _12250_);
  or (_12272_, _12247_, _11341_);
  and (_12273_, _12272_, _12271_);
  and (_12274_, _12249_, _11347_);
  or (_35875_, _12274_, _12273_);
  or (_12275_, _12246_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_12276_, _12275_, _12250_);
  or (_12277_, _12247_, _11544_);
  and (_12278_, _12277_, _12276_);
  and (_12279_, _12249_, _11550_);
  or (_35876_, _12279_, _12278_);
  or (_12280_, _12246_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_12281_, _12280_, _12250_);
  or (_12282_, _12247_, _11747_);
  and (_12283_, _12282_, _12281_);
  and (_12284_, _12249_, _11753_);
  or (_35877_, _12284_, _12283_);
  or (_12285_, _12246_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_12286_, _12285_, _12250_);
  or (_12287_, _12247_, _06182_);
  and (_12288_, _12287_, _12286_);
  and (_12289_, _12249_, _06209_);
  or (_35878_, _12289_, _12288_);
  nand (_12290_, _10357_, _04568_);
  or (_12291_, _12290_, _10534_);
  and (_12292_, _04557_, _03955_);
  not (_12293_, _12292_);
  nand (_12294_, _12290_, _03829_);
  and (_12295_, _12294_, _12293_);
  and (_12296_, _12295_, _12291_);
  and (_12297_, _12292_, _10546_);
  or (_35879_, _12297_, _12296_);
  or (_12298_, _12290_, _10749_);
  nand (_12299_, _12290_, _04011_);
  and (_12300_, _12299_, _12293_);
  and (_12301_, _12300_, _12298_);
  and (_12302_, _12292_, _10755_);
  or (_35880_, _12302_, _12301_);
  and (_12303_, _11937_, _04543_);
  or (_12304_, _12303_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_12305_, _12304_, _12293_);
  or (_12306_, _12290_, _10944_);
  and (_12307_, _12306_, _12305_);
  and (_12308_, _12292_, _10952_);
  or (_35881_, _12308_, _12307_);
  or (_12309_, _12303_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_12310_, _12309_, _12293_);
  or (_12311_, _12290_, _11139_);
  and (_12312_, _12311_, _12310_);
  and (_12313_, _12292_, _11145_);
  or (_35882_, _12313_, _12312_);
  or (_12314_, _12303_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_12315_, _12314_, _12293_);
  or (_12316_, _12290_, _11341_);
  and (_12317_, _12316_, _12315_);
  and (_12318_, _12292_, _11347_);
  or (_35883_, _12318_, _12317_);
  or (_12319_, _12303_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_12320_, _12319_, _12293_);
  or (_12321_, _12290_, _11544_);
  and (_12322_, _12321_, _12320_);
  and (_12323_, _12292_, _11550_);
  or (_35884_, _12323_, _12322_);
  or (_12324_, _12303_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_12325_, _12324_, _12293_);
  or (_12326_, _12290_, _11747_);
  and (_12327_, _12326_, _12325_);
  and (_12328_, _12292_, _11753_);
  or (_35885_, _12328_, _12327_);
  or (_12329_, _12303_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_12330_, _12329_, _12293_);
  or (_12331_, _12290_, _06182_);
  and (_12332_, _12331_, _12330_);
  and (_12333_, _12292_, _06209_);
  or (_35886_, _12333_, _12332_);
  and (_12334_, _11936_, _04127_);
  and (_12335_, _12334_, _04543_);
  or (_12336_, _12335_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_12337_, _04557_, _04215_);
  not (_12338_, _12337_);
  and (_12339_, _12338_, _12336_);
  nand (_12340_, _11760_, _04568_);
  or (_12341_, _12340_, _10534_);
  and (_12342_, _12341_, _12339_);
  and (_12343_, _12337_, _10546_);
  or (_35887_, _12343_, _12342_);
  or (_12344_, _12335_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_12345_, _12344_, _12338_);
  or (_12346_, _12340_, _10749_);
  and (_12347_, _12346_, _12345_);
  and (_12348_, _12337_, _10755_);
  or (_35888_, _12348_, _12347_);
  or (_12349_, _12335_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_12350_, _12349_, _12338_);
  or (_12351_, _12340_, _10944_);
  and (_12352_, _12351_, _12350_);
  and (_12353_, _12337_, _10952_);
  or (_35889_, _12353_, _12352_);
  or (_12354_, _12335_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_12355_, _12354_, _12338_);
  or (_12356_, _12340_, _11139_);
  and (_12357_, _12356_, _12355_);
  and (_12358_, _12337_, _11145_);
  or (_35890_, _12358_, _12357_);
  or (_12359_, _12335_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_12360_, _12359_, _12338_);
  or (_12361_, _12340_, _11341_);
  and (_12362_, _12361_, _12360_);
  and (_12363_, _12337_, _11347_);
  or (_35891_, _12363_, _12362_);
  or (_12364_, _12335_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_12365_, _12364_, _12338_);
  or (_12366_, _12340_, _11544_);
  and (_12367_, _12366_, _12365_);
  and (_12368_, _12337_, _11550_);
  or (_35892_, _12368_, _12367_);
  or (_12369_, _12335_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_12370_, _12369_, _12338_);
  or (_12371_, _12340_, _11747_);
  and (_12372_, _12371_, _12370_);
  and (_12373_, _12337_, _11753_);
  or (_35893_, _12373_, _12372_);
  or (_12374_, _12335_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_12375_, _12374_, _12338_);
  or (_12376_, _12340_, _06182_);
  and (_12377_, _12376_, _12375_);
  and (_12378_, _12337_, _06209_);
  or (_35894_, _12378_, _12377_);
  not (_12379_, _04568_);
  nor (_12380_, _11828_, _12379_);
  not (_12381_, _12380_);
  or (_12382_, _12381_, _10534_);
  and (_12383_, _05373_, _04557_);
  not (_12384_, _12383_);
  or (_12385_, _12380_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_12386_, _12385_, _12384_);
  and (_12387_, _12386_, _12382_);
  and (_12388_, _12383_, _10546_);
  or (_35895_, _12388_, _12387_);
  or (_12389_, _12381_, _10749_);
  or (_12390_, _12380_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_12391_, _12390_, _12384_);
  and (_12392_, _12391_, _12389_);
  and (_12393_, _12383_, _10755_);
  or (_35896_, _12393_, _12392_);
  and (_12394_, _11810_, _04543_);
  or (_12395_, _12394_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_12396_, _12395_, _12384_);
  or (_12397_, _12381_, _10944_);
  and (_12398_, _12397_, _12396_);
  and (_12399_, _12383_, _10952_);
  or (_35897_, _12399_, _12398_);
  or (_12400_, _12394_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_12401_, _12400_, _12384_);
  or (_12402_, _12381_, _11139_);
  and (_12403_, _12402_, _12401_);
  and (_12404_, _12383_, _11145_);
  or (_35898_, _12404_, _12403_);
  or (_12405_, _12394_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_12406_, _12405_, _12384_);
  or (_12407_, _12381_, _11341_);
  and (_12408_, _12407_, _12406_);
  and (_12409_, _12383_, _11347_);
  or (_35899_, _12409_, _12408_);
  or (_12410_, _12394_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_12411_, _12410_, _12384_);
  or (_12412_, _12381_, _11544_);
  and (_12413_, _12412_, _12411_);
  and (_12414_, _12383_, _11550_);
  or (_35900_, _12414_, _12413_);
  or (_12415_, _12394_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_12416_, _12415_, _12384_);
  or (_12417_, _12381_, _11747_);
  and (_12418_, _12417_, _12416_);
  and (_12419_, _12383_, _11753_);
  or (_35901_, _12419_, _12418_);
  or (_12420_, _12394_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_12421_, _12420_, _12384_);
  or (_12422_, _12381_, _06182_);
  and (_12423_, _12422_, _12421_);
  and (_12424_, _12383_, _06209_);
  or (_35902_, _12424_, _12423_);
  or (_12425_, _10534_, _04570_);
  or (_12426_, _04569_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_12427_, _12426_, _04559_);
  and (_12428_, _12427_, _12425_);
  and (_12429_, _10546_, _04558_);
  or (_35903_, _12429_, _12428_);
  or (_12430_, _10749_, _04570_);
  or (_12431_, _04569_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_12432_, _12431_, _04559_);
  and (_12433_, _12432_, _12430_);
  and (_12434_, _10755_, _04558_);
  or (_35904_, _12434_, _12433_);
  or (_12435_, _04544_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_12436_, _12435_, _04559_);
  or (_12437_, _10944_, _04570_);
  and (_12438_, _12437_, _12436_);
  and (_12439_, _10952_, _04558_);
  or (_35905_, _12439_, _12438_);
  or (_12440_, _04544_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_12441_, _12440_, _04559_);
  or (_12442_, _11139_, _04570_);
  and (_12443_, _12442_, _12441_);
  and (_12444_, _11145_, _04558_);
  or (_35906_, _12444_, _12443_);
  or (_12445_, _11341_, _04570_);
  or (_12446_, _04544_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_12447_, _12446_, _04559_);
  and (_12448_, _12447_, _12445_);
  and (_12449_, _11347_, _04558_);
  or (_35907_, _12449_, _12448_);
  or (_12450_, _04544_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_12451_, _12450_, _04559_);
  or (_12452_, _11544_, _04570_);
  and (_12453_, _12452_, _12451_);
  and (_12454_, _11550_, _04558_);
  or (_35908_, _12454_, _12453_);
  or (_12455_, _04544_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_12456_, _12455_, _04559_);
  or (_12458_, _11747_, _04570_);
  and (_12459_, _12458_, _12456_);
  and (_12460_, _11753_, _04558_);
  or (_35909_, _12460_, _12459_);
  nor (_12461_, _34655_, _06798_);
  and (_12462_, _06164_, _04721_);
  nor (_12463_, _04721_, _06798_);
  or (_12464_, _12463_, _02842_);
  or (_12465_, _12464_, _12462_);
  and (_12466_, _04721_, _03838_);
  or (_12467_, _12466_, _12463_);
  or (_12468_, _12467_, _02859_);
  nor (_12469_, _05321_, _06798_);
  and (_12470_, _10390_, _05321_);
  or (_12471_, _12470_, _12469_);
  and (_12472_, _12471_, _02884_);
  nor (_12473_, _05085_, _06220_);
  or (_12474_, _12473_, _12463_);
  or (_12475_, _12474_, _03006_);
  and (_12476_, _04721_, \oc8051_golden_model_1.ACC [0]);
  or (_12478_, _12476_, _12463_);
  and (_12479_, _12478_, _03845_);
  nor (_12480_, _03845_, _06798_);
  or (_12481_, _12480_, _02948_);
  or (_12482_, _12481_, _12479_);
  and (_12483_, _12482_, _02976_);
  or (_12484_, _12483_, _02877_);
  and (_12485_, _12484_, _12475_);
  and (_12486_, _12467_, _02946_);
  or (_12487_, _12486_, _02880_);
  or (_12488_, _12487_, _12485_);
  or (_12489_, _12488_, _12472_);
  or (_12490_, _12476_, _02992_);
  and (_12491_, _12490_, _02987_);
  or (_12492_, _12491_, _12463_);
  and (_12493_, _12492_, _06246_);
  and (_12494_, _12493_, _12489_);
  and (_12495_, _12474_, _02871_);
  or (_12496_, _12495_, _06252_);
  or (_12497_, _12496_, _12494_);
  nor (_12498_, _06734_, _06732_);
  nor (_12499_, _12498_, _06735_);
  or (_12500_, _12499_, _06258_);
  and (_12501_, _12500_, _02986_);
  and (_12502_, _12501_, _12497_);
  nor (_12503_, _10377_, _06773_);
  or (_12504_, _12503_, _12469_);
  and (_12505_, _12504_, _02866_);
  or (_12506_, _12505_, _05535_);
  or (_12507_, _12506_, _12502_);
  and (_12508_, _12507_, _12468_);
  or (_12509_, _12508_, _02841_);
  and (_12510_, _12509_, _12465_);
  or (_12511_, _12510_, _02567_);
  nor (_12512_, _10475_, _06220_);
  or (_12513_, _12463_, _02839_);
  or (_12514_, _12513_, _12512_);
  and (_12515_, _12514_, _06792_);
  and (_12516_, _12515_, _12511_);
  nand (_12517_, _07133_, _02696_);
  nor (_12518_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_12519_, _12518_, _06713_);
  or (_12520_, _07133_, _12519_);
  and (_12521_, _12520_, _06786_);
  and (_12522_, _12521_, _12517_);
  or (_12523_, _12522_, _08207_);
  or (_12524_, _12523_, _12516_);
  and (_12525_, _10372_, _04721_);
  or (_12526_, _12463_, _07139_);
  or (_12527_, _12526_, _12525_);
  and (_12528_, _04721_, _05660_);
  or (_12529_, _12528_, _12463_);
  or (_12530_, _12529_, _07140_);
  and (_12531_, _12530_, _07150_);
  and (_12532_, _12531_, _12527_);
  and (_12533_, _12532_, _12524_);
  and (_12534_, _10369_, _04721_);
  or (_12535_, _12534_, _12463_);
  and (_12536_, _12535_, _03148_);
  or (_12537_, _12536_, _12533_);
  and (_12538_, _12537_, _03138_);
  nand (_12539_, _12529_, _03022_);
  nor (_12540_, _12539_, _12473_);
  or (_12541_, _12463_, _05085_);
  and (_12542_, _12478_, _03137_);
  and (_12543_, _12542_, _12541_);
  or (_12544_, _12543_, _03042_);
  or (_12545_, _12544_, _12540_);
  or (_12546_, _12545_, _12538_);
  nor (_12547_, _10365_, _06220_);
  or (_12548_, _12463_, _03043_);
  or (_12549_, _12548_, _12547_);
  and (_12550_, _12549_, _07161_);
  and (_12551_, _12550_, _12546_);
  nor (_12552_, _10367_, _06220_);
  or (_12553_, _12552_, _12463_);
  and (_12554_, _12553_, _03143_);
  or (_12555_, _12554_, _03174_);
  or (_12556_, _12555_, _12551_);
  or (_12557_, _12474_, _03179_);
  and (_12558_, _12557_, _03183_);
  and (_12559_, _12558_, _12556_);
  and (_12560_, _12463_, _02799_);
  or (_12561_, _12560_, _02887_);
  or (_12562_, _12561_, _12559_);
  or (_12563_, _12474_, _02888_);
  and (_12564_, _12563_, _34655_);
  and (_12565_, _12564_, _12562_);
  or (_12566_, _12565_, _12461_);
  and (_35828_[0], _12566_, _35796_);
  nor (_12567_, _34655_, _06793_);
  nand (_12568_, _04721_, _03720_);
  or (_12569_, _04721_, \oc8051_golden_model_1.B [1]);
  and (_12570_, _12569_, _02834_);
  and (_12571_, _12570_, _12568_);
  and (_12572_, _10574_, _04721_);
  not (_12573_, _12572_);
  and (_12574_, _12573_, _12569_);
  or (_12575_, _12574_, _03006_);
  nand (_12576_, _04721_, _02543_);
  and (_12577_, _12576_, _12569_);
  and (_12578_, _12577_, _03845_);
  nor (_12579_, _03845_, _06793_);
  or (_12580_, _12579_, _02948_);
  or (_12581_, _12580_, _12578_);
  and (_12582_, _12581_, _02976_);
  and (_12583_, _12582_, _12575_);
  nor (_12584_, _04721_, _06793_);
  nor (_12585_, _06220_, _04020_);
  or (_12586_, _12585_, _12584_);
  and (_12587_, _12586_, _02946_);
  nor (_12588_, _05321_, _06793_);
  and (_12589_, _10569_, _05321_);
  or (_12590_, _12589_, _12588_);
  and (_12591_, _12590_, _02884_);
  or (_12592_, _12591_, _12587_);
  or (_12593_, _12592_, _02880_);
  or (_12594_, _12593_, _12583_);
  or (_12595_, _12577_, _02992_);
  and (_12596_, _12595_, _12594_);
  or (_12597_, _12596_, _02877_);
  and (_12598_, _10572_, _05321_);
  or (_12599_, _12598_, _12588_);
  or (_12600_, _12599_, _02987_);
  and (_12601_, _12600_, _06246_);
  and (_12602_, _12601_, _12597_);
  and (_12603_, _12589_, _10568_);
  or (_12604_, _12603_, _12588_);
  and (_12605_, _12604_, _02871_);
  or (_12606_, _12605_, _06252_);
  or (_12607_, _12606_, _12602_);
  nor (_12608_, _06737_, _06680_);
  nor (_12609_, _12608_, _06738_);
  or (_12610_, _12609_, _06258_);
  and (_12611_, _12610_, _02986_);
  and (_12612_, _12611_, _12607_);
  nor (_12613_, _10618_, _06773_);
  or (_12614_, _12613_, _12588_);
  and (_12615_, _12614_, _02866_);
  or (_12616_, _12615_, _05535_);
  or (_12617_, _12616_, _12612_);
  or (_12618_, _12586_, _02859_);
  and (_12619_, _12618_, _12617_);
  or (_12620_, _12619_, _02841_);
  and (_12621_, _06163_, _04721_);
  or (_12622_, _12584_, _02842_);
  or (_12623_, _12622_, _12621_);
  and (_12624_, _12623_, _02839_);
  and (_12625_, _12624_, _12620_);
  or (_12626_, _10674_, _06220_);
  and (_12627_, _12569_, _02567_);
  and (_12628_, _12627_, _12626_);
  or (_12629_, _12628_, _06786_);
  or (_12630_, _12629_, _12625_);
  and (_12631_, _07133_, _07080_);
  nor (_12632_, _07128_, _07127_);
  or (_12633_, _12632_, _07129_);
  nor (_12634_, _12633_, _07133_);
  or (_12635_, _12634_, _12631_);
  or (_12636_, _12635_, _06792_);
  and (_12637_, _12636_, _07140_);
  and (_12638_, _12637_, _12630_);
  or (_12639_, _12638_, _12571_);
  and (_12640_, _12639_, _03910_);
  or (_12641_, _10688_, _06220_);
  and (_12642_, _12569_, _03022_);
  and (_12643_, _12642_, _12641_);
  or (_12644_, _10565_, _06220_);
  and (_12645_, _12569_, _03148_);
  and (_12646_, _12645_, _12644_);
  or (_12647_, _10689_, _06220_);
  and (_12648_, _12569_, _03051_);
  and (_12649_, _12648_, _12647_);
  or (_12650_, _12649_, _12646_);
  or (_12651_, _12650_, _12643_);
  or (_12652_, _12651_, _12640_);
  and (_12653_, _12652_, _06213_);
  or (_12654_, _12584_, _05038_);
  and (_12655_, _12577_, _03137_);
  and (_12656_, _12655_, _12654_);
  or (_12657_, _12656_, _12653_);
  and (_12658_, _12657_, _03144_);
  or (_12659_, _12568_, _05038_);
  and (_12660_, _12569_, _03042_);
  and (_12661_, _12660_, _12659_);
  or (_12662_, _12576_, _05038_);
  and (_12663_, _12569_, _03143_);
  and (_12664_, _12663_, _12662_);
  or (_12665_, _12664_, _03174_);
  or (_12666_, _12665_, _12661_);
  or (_12667_, _12666_, _12658_);
  or (_12668_, _12574_, _03179_);
  and (_12669_, _12668_, _03183_);
  and (_12670_, _12669_, _12667_);
  and (_12671_, _12599_, _02799_);
  or (_12672_, _12671_, _02887_);
  or (_12673_, _12672_, _12670_);
  or (_12674_, _12584_, _02888_);
  or (_12675_, _12674_, _12572_);
  and (_12676_, _12675_, _34655_);
  and (_12677_, _12676_, _12673_);
  or (_12678_, _12677_, _12567_);
  and (_35828_[1], _12678_, _35796_);
  nor (_12679_, _34655_, _06951_);
  nor (_12680_, _04721_, _06951_);
  nor (_12681_, _06220_, _04449_);
  or (_12682_, _12681_, _12680_);
  or (_12683_, _12682_, _02859_);
  and (_12684_, _04721_, \oc8051_golden_model_1.ACC [2]);
  or (_12685_, _12684_, _12680_);
  or (_12686_, _12685_, _02992_);
  nor (_12687_, _10788_, _06220_);
  or (_12688_, _12687_, _12680_);
  or (_12689_, _12688_, _03006_);
  and (_12690_, _12685_, _03845_);
  nor (_12691_, _03845_, _06951_);
  or (_12692_, _12691_, _02948_);
  or (_12693_, _12692_, _12690_);
  and (_12694_, _12693_, _02976_);
  and (_12695_, _12694_, _12689_);
  nor (_12696_, _05321_, _06951_);
  and (_12697_, _10792_, _05321_);
  or (_12698_, _12697_, _12696_);
  and (_12699_, _12698_, _02884_);
  and (_12700_, _12682_, _02946_);
  or (_12701_, _12700_, _02880_);
  or (_12702_, _12701_, _12699_);
  or (_12703_, _12702_, _12695_);
  and (_12704_, _12703_, _12686_);
  or (_12705_, _12704_, _02877_);
  and (_12706_, _10773_, _05321_);
  or (_12707_, _12706_, _12696_);
  or (_12708_, _12707_, _02987_);
  and (_12709_, _12708_, _06246_);
  and (_12710_, _12709_, _12705_);
  or (_12711_, _12696_, _10807_);
  and (_12712_, _12711_, _02871_);
  and (_12713_, _12712_, _12698_);
  or (_12714_, _12713_, _06252_);
  or (_12715_, _12714_, _12710_);
  nor (_12716_, _06740_, _06635_);
  nor (_12717_, _12716_, _06741_);
  or (_12718_, _12717_, _06258_);
  and (_12719_, _12718_, _02986_);
  and (_12720_, _12719_, _12715_);
  nor (_12721_, _10825_, _06773_);
  or (_12722_, _12721_, _12696_);
  and (_12723_, _12722_, _02866_);
  or (_12724_, _12723_, _05535_);
  or (_12725_, _12724_, _12720_);
  and (_12726_, _12725_, _12683_);
  or (_12727_, _12726_, _02841_);
  and (_12728_, _06167_, _04721_);
  or (_12729_, _12680_, _02842_);
  or (_12730_, _12729_, _12728_);
  and (_12731_, _12730_, _12727_);
  or (_12732_, _12731_, _02567_);
  nor (_12733_, _10881_, _06220_);
  or (_12734_, _12680_, _02839_);
  or (_12735_, _12734_, _12733_);
  and (_12736_, _12735_, _06792_);
  and (_12737_, _12736_, _12732_);
  not (_12738_, _07133_);
  or (_12739_, _12738_, _07070_);
  nor (_12740_, _07129_, _07081_);
  not (_12741_, _12740_);
  and (_12742_, _12741_, _07073_);
  nor (_12743_, _12741_, _07073_);
  nor (_12744_, _12743_, _12742_);
  or (_12745_, _12744_, _07133_);
  and (_12746_, _12745_, _06786_);
  and (_12747_, _12746_, _12739_);
  or (_12748_, _12747_, _08207_);
  or (_12749_, _12748_, _12737_);
  and (_12750_, _10770_, _04721_);
  or (_12751_, _12680_, _07139_);
  or (_12752_, _12751_, _12750_);
  and (_12753_, _04721_, _05693_);
  or (_12754_, _12753_, _12680_);
  or (_12755_, _12754_, _07140_);
  and (_12756_, _12755_, _07150_);
  and (_12757_, _12756_, _12752_);
  and (_12758_, _12757_, _12749_);
  and (_12759_, _10766_, _04721_);
  or (_12760_, _12759_, _12680_);
  and (_12761_, _12760_, _03148_);
  or (_12762_, _12761_, _12758_);
  and (_12763_, _12762_, _03138_);
  or (_12764_, _12680_, _05135_);
  and (_12765_, _12685_, _03137_);
  and (_12766_, _12754_, _03022_);
  or (_12767_, _12766_, _12765_);
  and (_12768_, _12767_, _12764_);
  or (_12769_, _12768_, _03042_);
  or (_12770_, _12769_, _12763_);
  nor (_12771_, _10768_, _06220_);
  or (_12772_, _12680_, _03043_);
  or (_12773_, _12772_, _12771_);
  and (_12774_, _12773_, _07161_);
  and (_12775_, _12774_, _12770_);
  nor (_12776_, _10765_, _06220_);
  or (_12777_, _12776_, _12680_);
  and (_12778_, _12777_, _03143_);
  or (_12779_, _12778_, _03174_);
  or (_12780_, _12779_, _12775_);
  or (_12781_, _12688_, _03179_);
  and (_12782_, _12781_, _03183_);
  and (_12783_, _12782_, _12780_);
  and (_12784_, _12707_, _02799_);
  or (_12785_, _12784_, _02887_);
  or (_12786_, _12785_, _12783_);
  and (_12787_, _10941_, _04721_);
  or (_12788_, _12680_, _02888_);
  or (_12789_, _12788_, _12787_);
  and (_12790_, _12789_, _34655_);
  and (_12791_, _12790_, _12786_);
  or (_12792_, _12791_, _12679_);
  and (_35828_[2], _12792_, _35796_);
  nor (_12793_, _34655_, _06876_);
  nor (_12794_, _04721_, _06876_);
  nor (_12795_, _06220_, _04275_);
  or (_12796_, _12795_, _12794_);
  or (_12797_, _12796_, _02859_);
  nor (_12798_, _10983_, _06220_);
  or (_12799_, _12798_, _12794_);
  or (_12800_, _12799_, _03006_);
  and (_12801_, _04721_, \oc8051_golden_model_1.ACC [3]);
  or (_12802_, _12801_, _12794_);
  and (_12803_, _12802_, _03845_);
  nor (_12804_, _03845_, _06876_);
  or (_12805_, _12804_, _02948_);
  or (_12806_, _12805_, _12803_);
  and (_12807_, _12806_, _02976_);
  and (_12808_, _12807_, _12800_);
  and (_12809_, _12796_, _02946_);
  nor (_12810_, _05321_, _06876_);
  and (_12811_, _10976_, _05321_);
  or (_12812_, _12811_, _12810_);
  and (_12813_, _12812_, _02884_);
  or (_12814_, _12813_, _12809_);
  or (_12815_, _12814_, _02880_);
  or (_12816_, _12815_, _12808_);
  or (_12817_, _12802_, _02992_);
  and (_12818_, _12817_, _12816_);
  or (_12819_, _12818_, _02877_);
  and (_12820_, _10979_, _05321_);
  or (_12821_, _12820_, _12810_);
  or (_12822_, _12821_, _02987_);
  and (_12823_, _12822_, _06246_);
  and (_12824_, _12823_, _12819_);
  and (_12825_, _12811_, _10975_);
  or (_12826_, _12825_, _12810_);
  and (_12827_, _12826_, _02871_);
  or (_12828_, _12827_, _06252_);
  or (_12829_, _12828_, _12824_);
  nor (_12830_, _06743_, _06577_);
  nor (_12831_, _12830_, _06744_);
  or (_12832_, _12831_, _06258_);
  and (_12833_, _12832_, _02986_);
  and (_12834_, _12833_, _12829_);
  nor (_12835_, _10973_, _06773_);
  or (_12836_, _12835_, _12810_);
  and (_12837_, _12836_, _02866_);
  or (_12838_, _12837_, _05535_);
  or (_12839_, _12838_, _12834_);
  and (_12840_, _12839_, _12797_);
  or (_12841_, _12840_, _02841_);
  and (_12842_, _06166_, _04721_);
  or (_12843_, _12794_, _02842_);
  or (_12844_, _12843_, _12842_);
  and (_12845_, _12844_, _12841_);
  or (_12846_, _12845_, _02567_);
  nor (_12847_, _11076_, _06220_);
  or (_12848_, _12794_, _02839_);
  or (_12849_, _12848_, _12847_);
  and (_12850_, _12849_, _06792_);
  and (_12851_, _12850_, _12846_);
  nor (_12852_, _12742_, _07072_);
  nor (_12853_, _12852_, _07065_);
  and (_12854_, _12852_, _07065_);
  or (_12855_, _12854_, _12853_);
  or (_12856_, _12855_, _07133_);
  or (_12857_, _12738_, _07062_);
  and (_12858_, _12857_, _06786_);
  and (_12859_, _12858_, _12856_);
  or (_12860_, _12859_, _08207_);
  or (_12861_, _12860_, _12851_);
  and (_12862_, _10968_, _04721_);
  or (_12863_, _12794_, _07139_);
  or (_12864_, _12863_, _12862_);
  and (_12865_, _04721_, _05654_);
  or (_12866_, _12865_, _12794_);
  or (_12867_, _12866_, _07140_);
  and (_12868_, _12867_, _07150_);
  and (_12869_, _12868_, _12864_);
  and (_12870_, _12869_, _12861_);
  and (_12871_, _10964_, _04721_);
  or (_12872_, _12871_, _12794_);
  and (_12873_, _12872_, _03148_);
  or (_12874_, _12873_, _12870_);
  and (_12875_, _12874_, _03138_);
  or (_12876_, _12794_, _04993_);
  and (_12877_, _12802_, _03137_);
  and (_12878_, _12866_, _03022_);
  or (_12879_, _12878_, _12877_);
  and (_12880_, _12879_, _12876_);
  or (_12881_, _12880_, _03042_);
  or (_12882_, _12881_, _12875_);
  nor (_12883_, _10967_, _06220_);
  or (_12884_, _12794_, _03043_);
  or (_12885_, _12884_, _12883_);
  and (_12886_, _12885_, _07161_);
  and (_12887_, _12886_, _12882_);
  nor (_12888_, _10962_, _06220_);
  or (_12889_, _12888_, _12794_);
  and (_12890_, _12889_, _03143_);
  or (_12891_, _12890_, _03174_);
  or (_12892_, _12891_, _12887_);
  or (_12893_, _12799_, _03179_);
  and (_12894_, _12893_, _03183_);
  and (_12895_, _12894_, _12892_);
  and (_12896_, _12821_, _02799_);
  or (_12897_, _12896_, _02887_);
  or (_12898_, _12897_, _12895_);
  and (_12899_, _11136_, _04721_);
  or (_12900_, _12794_, _02888_);
  or (_12901_, _12900_, _12899_);
  and (_12902_, _12901_, _34655_);
  and (_12903_, _12902_, _12898_);
  or (_12904_, _12903_, _12793_);
  and (_35828_[3], _12904_, _35796_);
  nor (_12905_, _34655_, _06930_);
  nor (_12906_, _04721_, _06930_);
  nor (_12907_, _11271_, _06220_);
  or (_12908_, _12907_, _12906_);
  and (_12909_, _12908_, _02567_);
  nor (_12910_, _05192_, _06220_);
  or (_12911_, _12910_, _12906_);
  or (_12912_, _12911_, _02859_);
  nor (_12913_, _11184_, _06220_);
  or (_12914_, _12913_, _12906_);
  or (_12915_, _12914_, _03006_);
  and (_12916_, _04721_, \oc8051_golden_model_1.ACC [4]);
  or (_12917_, _12916_, _12906_);
  and (_12918_, _12917_, _03845_);
  nor (_12919_, _03845_, _06930_);
  or (_12920_, _12919_, _02948_);
  or (_12921_, _12920_, _12918_);
  and (_12922_, _12921_, _02976_);
  and (_12923_, _12922_, _12915_);
  and (_12924_, _12911_, _02946_);
  nor (_12925_, _05321_, _06930_);
  and (_12926_, _11167_, _05321_);
  or (_12927_, _12926_, _12925_);
  and (_12928_, _12927_, _02884_);
  or (_12929_, _12928_, _12924_);
  or (_12930_, _12929_, _02880_);
  or (_12931_, _12930_, _12923_);
  or (_12932_, _12917_, _02992_);
  and (_12933_, _12932_, _12931_);
  or (_12934_, _12933_, _02877_);
  and (_12935_, _11165_, _05321_);
  or (_12936_, _12935_, _12925_);
  or (_12937_, _12936_, _02987_);
  and (_12938_, _12937_, _06246_);
  and (_12939_, _12938_, _12934_);
  or (_12940_, _12925_, _11201_);
  and (_12941_, _12940_, _12927_);
  and (_12942_, _12941_, _02871_);
  or (_12943_, _12942_, _06252_);
  or (_12944_, _12943_, _12939_);
  nor (_12945_, _06748_, _06746_);
  nor (_12946_, _12945_, _06749_);
  or (_12947_, _12946_, _06258_);
  and (_12948_, _12947_, _02986_);
  and (_12949_, _12948_, _12944_);
  nor (_12950_, _11163_, _06773_);
  or (_12951_, _12950_, _12925_);
  and (_12952_, _12951_, _02866_);
  or (_12953_, _12952_, _05535_);
  or (_12954_, _12953_, _12949_);
  and (_12955_, _12954_, _12912_);
  or (_12956_, _12955_, _02841_);
  and (_12957_, _06171_, _04721_);
  or (_12958_, _12906_, _02842_);
  or (_12959_, _12958_, _12957_);
  and (_12960_, _12959_, _02839_);
  and (_12961_, _12960_, _12956_);
  or (_12962_, _12961_, _12909_);
  and (_12963_, _12962_, _06792_);
  nand (_12964_, _07133_, _07100_);
  nor (_12965_, _12852_, _07063_);
  or (_12966_, _12965_, _07064_);
  nand (_12967_, _12966_, _07103_);
  or (_12968_, _12966_, _07103_);
  and (_12969_, _12968_, _12967_);
  or (_12970_, _12969_, _07133_);
  and (_12971_, _12970_, _06786_);
  and (_12972_, _12971_, _12964_);
  or (_12973_, _12972_, _08207_);
  or (_12974_, _12973_, _12963_);
  and (_12975_, _11158_, _04721_);
  or (_12976_, _12906_, _07139_);
  or (_12977_, _12976_, _12975_);
  and (_12978_, _05618_, _04721_);
  or (_12979_, _12978_, _12906_);
  or (_12980_, _12979_, _07140_);
  and (_12981_, _12980_, _07150_);
  and (_12982_, _12981_, _12977_);
  and (_12983_, _12982_, _12974_);
  and (_12984_, _11154_, _04721_);
  or (_12985_, _12984_, _12906_);
  and (_12986_, _12985_, _03148_);
  or (_12987_, _12986_, _12983_);
  and (_12988_, _12987_, _03138_);
  or (_12989_, _12906_, _05240_);
  and (_12990_, _12917_, _03137_);
  and (_12991_, _12979_, _03022_);
  or (_12992_, _12991_, _12990_);
  and (_12993_, _12992_, _12989_);
  or (_12994_, _12993_, _03042_);
  or (_12995_, _12994_, _12988_);
  nor (_12996_, _11157_, _06220_);
  or (_12997_, _12906_, _03043_);
  or (_12998_, _12997_, _12996_);
  and (_12999_, _12998_, _07161_);
  and (_13000_, _12999_, _12995_);
  nor (_13001_, _11152_, _06220_);
  or (_13002_, _13001_, _12906_);
  and (_13003_, _13002_, _03143_);
  or (_13004_, _13003_, _03174_);
  or (_13005_, _13004_, _13000_);
  or (_13006_, _12914_, _03179_);
  and (_13007_, _13006_, _03183_);
  and (_13008_, _13007_, _13005_);
  and (_13009_, _12936_, _02799_);
  or (_13010_, _13009_, _02887_);
  or (_13011_, _13010_, _13008_);
  and (_13012_, _11338_, _04721_);
  or (_13013_, _12906_, _02888_);
  or (_13014_, _13013_, _13012_);
  and (_13015_, _13014_, _34655_);
  and (_13016_, _13015_, _13011_);
  or (_13017_, _13016_, _12905_);
  and (_35828_[4], _13017_, _35796_);
  nor (_13018_, _34655_, _06919_);
  nor (_13019_, _04721_, _06919_);
  nor (_13020_, _11467_, _06220_);
  or (_13021_, _13020_, _13019_);
  and (_13022_, _13021_, _02567_);
  nor (_13023_, _11380_, _06220_);
  or (_13024_, _13023_, _13019_);
  or (_13025_, _13024_, _03006_);
  and (_13026_, _04721_, \oc8051_golden_model_1.ACC [5]);
  or (_13027_, _13026_, _13019_);
  and (_13028_, _13027_, _03845_);
  nor (_13029_, _03845_, _06919_);
  or (_13030_, _13029_, _02948_);
  or (_13031_, _13030_, _13028_);
  and (_13032_, _13031_, _02976_);
  and (_13033_, _13032_, _13025_);
  nor (_13034_, _04894_, _06220_);
  or (_13035_, _13034_, _13019_);
  and (_13036_, _13035_, _02946_);
  nor (_13037_, _05321_, _06919_);
  and (_13038_, _11365_, _05321_);
  or (_13039_, _13038_, _13037_);
  and (_13040_, _13039_, _02884_);
  or (_13041_, _13040_, _13036_);
  or (_13042_, _13041_, _02880_);
  or (_13043_, _13042_, _13033_);
  or (_13044_, _13027_, _02992_);
  and (_13045_, _13044_, _13043_);
  or (_13046_, _13045_, _02877_);
  and (_13047_, _11363_, _05321_);
  or (_13048_, _13047_, _13037_);
  or (_13049_, _13048_, _02987_);
  and (_13050_, _13049_, _06246_);
  and (_13051_, _13050_, _13046_);
  or (_13052_, _13037_, _11397_);
  and (_13053_, _13052_, _02871_);
  and (_13054_, _13053_, _13039_);
  or (_13055_, _13054_, _06252_);
  or (_13056_, _13055_, _13051_);
  or (_13057_, _06449_, _06450_);
  and (_13058_, _13057_, _06750_);
  nor (_13059_, _13058_, _06751_);
  or (_13060_, _13059_, _06258_);
  and (_13061_, _13060_, _02986_);
  and (_13062_, _13061_, _13056_);
  nor (_13063_, _11361_, _06773_);
  or (_13064_, _13063_, _13037_);
  and (_13065_, _13064_, _02866_);
  or (_13066_, _13065_, _05535_);
  or (_13067_, _13066_, _13062_);
  or (_13068_, _13035_, _02859_);
  and (_13069_, _13068_, _13067_);
  or (_13070_, _13069_, _02841_);
  and (_13071_, _06170_, _04721_);
  or (_13072_, _13019_, _02842_);
  or (_13073_, _13072_, _13071_);
  and (_13074_, _13073_, _02839_);
  and (_13075_, _13074_, _13070_);
  or (_13076_, _13075_, _13022_);
  and (_13077_, _13076_, _06792_);
  or (_13078_, _12738_, _07110_);
  not (_13079_, _07102_);
  and (_13080_, _12967_, _13079_);
  nor (_13081_, _13080_, _07113_);
  and (_13082_, _13080_, _07113_);
  or (_13083_, _13082_, _13081_);
  or (_13084_, _13083_, _07133_);
  and (_13085_, _13084_, _06786_);
  and (_13086_, _13085_, _13078_);
  or (_13087_, _13086_, _08207_);
  or (_13088_, _13087_, _13077_);
  and (_13089_, _11482_, _04721_);
  or (_13090_, _13019_, _07139_);
  or (_13091_, _13090_, _13089_);
  and (_13092_, _05671_, _04721_);
  or (_13093_, _13092_, _13019_);
  or (_13094_, _13093_, _07140_);
  and (_13095_, _13094_, _07150_);
  and (_13096_, _13095_, _13091_);
  and (_13097_, _13096_, _13088_);
  and (_13098_, _11356_, _04721_);
  or (_13099_, _13098_, _13019_);
  and (_13100_, _13099_, _03148_);
  or (_13101_, _13100_, _13097_);
  and (_13102_, _13101_, _03138_);
  or (_13103_, _13019_, _04945_);
  and (_13104_, _13027_, _03137_);
  and (_13105_, _13093_, _03022_);
  or (_13106_, _13105_, _13104_);
  and (_13107_, _13106_, _13103_);
  or (_13108_, _13107_, _03042_);
  or (_13109_, _13108_, _13102_);
  nor (_13110_, _11480_, _06220_);
  or (_13111_, _13019_, _03043_);
  or (_13112_, _13111_, _13110_);
  and (_13113_, _13112_, _07161_);
  and (_13114_, _13113_, _13109_);
  nor (_13115_, _11355_, _06220_);
  or (_13116_, _13115_, _13019_);
  and (_13117_, _13116_, _03143_);
  or (_13118_, _13117_, _03174_);
  or (_13119_, _13118_, _13114_);
  or (_13120_, _13024_, _03179_);
  and (_13121_, _13120_, _03183_);
  and (_13122_, _13121_, _13119_);
  and (_13123_, _13048_, _02799_);
  or (_13124_, _13123_, _02887_);
  or (_13125_, _13124_, _13122_);
  and (_13126_, _11541_, _04721_);
  or (_13127_, _13019_, _02888_);
  or (_13128_, _13127_, _13126_);
  and (_13129_, _13128_, _34655_);
  and (_13130_, _13129_, _13125_);
  or (_13131_, _13130_, _13018_);
  and (_35828_[5], _13131_, _35796_);
  not (_13132_, \oc8051_golden_model_1.B [6]);
  nor (_13133_, _34655_, _13132_);
  nor (_13134_, _04721_, _13132_);
  nor (_13135_, _11671_, _06220_);
  or (_13136_, _13135_, _13134_);
  and (_13137_, _13136_, _02567_);
  nor (_13138_, _11567_, _06220_);
  or (_13139_, _13138_, _13134_);
  or (_13140_, _13139_, _03006_);
  and (_13141_, _04721_, \oc8051_golden_model_1.ACC [6]);
  or (_13142_, _13141_, _13134_);
  and (_13143_, _13142_, _03845_);
  nor (_13144_, _03845_, _13132_);
  or (_13145_, _13144_, _02948_);
  or (_13146_, _13145_, _13143_);
  and (_13147_, _13146_, _02976_);
  and (_13148_, _13147_, _13140_);
  nor (_13149_, _04790_, _06220_);
  or (_13150_, _13149_, _13134_);
  and (_13151_, _13150_, _02946_);
  nor (_13152_, _05321_, _13132_);
  and (_13153_, _11564_, _05321_);
  or (_13154_, _13153_, _13152_);
  and (_13155_, _13154_, _02884_);
  or (_13156_, _13155_, _13151_);
  or (_13157_, _13156_, _02880_);
  or (_13158_, _13157_, _13148_);
  or (_13159_, _13142_, _02992_);
  and (_13160_, _13159_, _13158_);
  or (_13161_, _13160_, _02877_);
  and (_13162_, _11562_, _05321_);
  or (_13163_, _13162_, _13152_);
  or (_13164_, _13163_, _02987_);
  and (_13165_, _13164_, _06246_);
  and (_13166_, _13165_, _13161_);
  or (_13167_, _13152_, _11596_);
  and (_13168_, _13167_, _02871_);
  and (_13169_, _13168_, _13154_);
  or (_13170_, _13169_, _06252_);
  or (_13171_, _13170_, _13166_);
  nor (_13172_, _06765_, _06752_);
  nor (_13173_, _13172_, _06766_);
  or (_13174_, _13173_, _06258_);
  and (_13175_, _13174_, _02986_);
  and (_13176_, _13175_, _13171_);
  nor (_13177_, _11614_, _06773_);
  or (_13178_, _13177_, _13152_);
  and (_13179_, _13178_, _02866_);
  or (_13180_, _13179_, _05535_);
  or (_13181_, _13180_, _13176_);
  or (_13182_, _13150_, _02859_);
  and (_13183_, _13182_, _13181_);
  or (_13184_, _13183_, _02841_);
  and (_13185_, _06162_, _04721_);
  or (_13186_, _13134_, _02842_);
  or (_13187_, _13186_, _13185_);
  and (_13188_, _13187_, _02839_);
  and (_13189_, _13188_, _13184_);
  or (_13190_, _13189_, _13137_);
  and (_13191_, _13190_, _06792_);
  nor (_13192_, _13080_, _07111_);
  or (_13193_, _13192_, _07112_);
  and (_13194_, _13193_, _07094_);
  nor (_13195_, _13193_, _07094_);
  or (_13196_, _13195_, _13194_);
  or (_13197_, _13196_, _07133_);
  nand (_13198_, _07133_, _07052_);
  and (_13199_, _13198_, _06786_);
  and (_13200_, _13199_, _13197_);
  or (_13201_, _13200_, _08207_);
  or (_13202_, _13201_, _13191_);
  and (_13203_, _11560_, _04721_);
  or (_13204_, _13134_, _07139_);
  or (_13205_, _13204_, _13203_);
  and (_13206_, _11678_, _04721_);
  or (_13207_, _13206_, _13134_);
  or (_13208_, _13207_, _07140_);
  and (_13209_, _13208_, _07150_);
  and (_13210_, _13209_, _13205_);
  and (_13211_, _13210_, _13202_);
  and (_13212_, _11556_, _04721_);
  or (_13213_, _13212_, _13134_);
  and (_13214_, _13213_, _03148_);
  or (_13215_, _13214_, _13211_);
  and (_13216_, _13215_, _03138_);
  or (_13217_, _13134_, _04838_);
  and (_13218_, _13142_, _03137_);
  and (_13219_, _13207_, _03022_);
  or (_13220_, _13219_, _13218_);
  and (_13221_, _13220_, _13217_);
  or (_13222_, _13221_, _03042_);
  or (_13223_, _13222_, _13216_);
  nor (_13224_, _11558_, _06220_);
  or (_13225_, _13134_, _03043_);
  or (_13226_, _13225_, _13224_);
  and (_13227_, _13226_, _07161_);
  and (_13228_, _13227_, _13223_);
  nor (_13229_, _11555_, _06220_);
  or (_13230_, _13229_, _13134_);
  and (_13231_, _13230_, _03143_);
  or (_13232_, _13231_, _03174_);
  or (_13233_, _13232_, _13228_);
  or (_13234_, _13139_, _03179_);
  and (_13235_, _13234_, _03183_);
  and (_13236_, _13235_, _13233_);
  and (_13237_, _13163_, _02799_);
  or (_13238_, _13237_, _02887_);
  or (_13239_, _13238_, _13236_);
  and (_13240_, _11744_, _04721_);
  or (_13241_, _13134_, _02888_);
  or (_13242_, _13241_, _13240_);
  and (_13243_, _13242_, _34655_);
  and (_13244_, _13243_, _13239_);
  or (_13245_, _13244_, _13133_);
  and (_35828_[6], _13245_, _35796_);
  nor (_13246_, _34655_, _02696_);
  nand (_13247_, _08115_, _05364_);
  and (_13248_, _05945_, _02696_);
  nor (_13249_, _08051_, _13248_);
  not (_13250_, _13249_);
  nand (_13251_, _13250_, _03571_);
  nand (_13252_, _07964_, _07780_);
  nand (_13253_, _07921_, _09271_);
  or (_13254_, _10368_, _03136_);
  and (_13255_, _13254_, _07312_);
  and (_13256_, _07883_, _07212_);
  nor (_13257_, _04731_, _02696_);
  and (_13258_, _10372_, _04731_);
  nor (_13259_, _13258_, _13257_);
  nand (_13260_, _13259_, _03051_);
  not (_13261_, _03521_);
  or (_13262_, _13249_, _13261_);
  and (_13263_, _04731_, _03838_);
  nor (_13264_, _13263_, _13257_);
  nand (_13265_, _13264_, _05535_);
  nand (_13266_, _07780_, _07540_);
  or (_13267_, _07402_, _03838_);
  nor (_13268_, _05313_, _02696_);
  and (_13269_, _10390_, _05313_);
  nor (_13270_, _13269_, _13268_);
  nand (_13271_, _13270_, _02884_);
  and (_13272_, _13271_, _07474_);
  nor (_13273_, _07607_, _03401_);
  or (_13274_, _07411_, _06164_);
  not (_13275_, _07421_);
  and (_13276_, _13275_, _03838_);
  or (_13277_, _07423_, \oc8051_golden_model_1.ACC [0]);
  nand (_13278_, _07423_, \oc8051_golden_model_1.ACC [0]);
  and (_13279_, _13278_, _13277_);
  and (_13280_, _13279_, _07421_);
  or (_13281_, _13280_, _07410_);
  or (_13282_, _13281_, _13276_);
  and (_13283_, _13282_, _03401_);
  and (_13284_, _13283_, _13274_);
  or (_13285_, _13284_, _13273_);
  and (_13286_, _13285_, _07437_);
  and (_13287_, _07441_, xram_data_in_reg[0]);
  or (_13288_, _13287_, _03840_);
  or (_13289_, _13288_, _13286_);
  or (_13290_, _06164_, _05371_);
  and (_13291_, _13290_, _03006_);
  and (_13292_, _13291_, _13289_);
  nor (_13293_, _05085_, _07319_);
  nor (_13294_, _13293_, _13257_);
  nor (_13295_, _13294_, _03006_);
  or (_13296_, _13295_, _02884_);
  or (_13297_, _13296_, _13292_);
  and (_13298_, _13297_, _13272_);
  nor (_13299_, _13264_, _07474_);
  or (_13300_, _13299_, _07403_);
  or (_13301_, _13300_, _13298_);
  and (_13302_, _13301_, _13267_);
  or (_13303_, _13302_, _03873_);
  or (_13304_, _06164_, _07481_);
  and (_13305_, _13304_, _02992_);
  and (_13306_, _13305_, _13303_);
  nor (_13307_, _07607_, _02992_);
  or (_13308_, _13307_, _07485_);
  or (_13309_, _13308_, _13306_);
  nand (_13310_, _07485_, _06864_);
  and (_13311_, _13310_, _13309_);
  or (_13312_, _13311_, _02877_);
  or (_13313_, _13257_, _02987_);
  and (_13314_, _13313_, _06246_);
  and (_13315_, _13314_, _13312_);
  nor (_13316_, _13294_, _06246_);
  or (_13317_, _13316_, _06252_);
  or (_13318_, _13317_, _13315_);
  not (_13319_, _06713_);
  nand (_13320_, _13319_, _06252_);
  and (_13321_, _13320_, _07399_);
  and (_13322_, _13321_, _13318_);
  nand (_13323_, _07521_, _07507_);
  and (_13324_, _13323_, _09326_);
  or (_13325_, _13324_, _13322_);
  nand (_13326_, _07397_, _07386_);
  and (_13327_, _13326_, _02991_);
  and (_13328_, _13327_, _13325_);
  nand (_13329_, _07697_, _07541_);
  and (_13330_, _13329_, _09325_);
  or (_13331_, _13330_, _13328_);
  and (_13332_, _13331_, _13266_);
  or (_13333_, _13332_, _07721_);
  or (_13334_, _02833_, _02571_);
  and (_13335_, _13334_, _02986_);
  and (_13336_, _13335_, _13333_);
  nor (_13337_, _10377_, _07806_);
  nor (_13338_, _13337_, _13268_);
  nor (_13339_, _13338_, _02986_);
  or (_13340_, _13339_, _05535_);
  or (_13341_, _13340_, _13336_);
  and (_13342_, _13341_, _13265_);
  or (_13343_, _13342_, _02841_);
  and (_13344_, _06164_, _04731_);
  nor (_13345_, _13344_, _13257_);
  nand (_13346_, _13345_, _02841_);
  and (_13347_, _13346_, _02839_);
  and (_13348_, _13347_, _13343_);
  nor (_13349_, _10475_, _07319_);
  nor (_13350_, _13349_, _13257_);
  nor (_13351_, _13350_, _02839_);
  or (_13352_, _13351_, _06786_);
  or (_13353_, _13352_, _13348_);
  nand (_13354_, _07133_, _06786_);
  and (_13355_, _13354_, _13353_);
  and (_13356_, _13355_, _02609_);
  and (_13357_, _02833_, _02542_);
  or (_13358_, _13357_, _02834_);
  or (_13359_, _13358_, _13356_);
  and (_13360_, _04731_, _05660_);
  nor (_13361_, _13360_, _13257_);
  nand (_13362_, _13361_, _02834_);
  and (_13363_, _13362_, _07831_);
  and (_13364_, _13363_, _13359_);
  and (_13365_, _07830_, _02833_);
  or (_13366_, _13365_, _07843_);
  or (_13367_, _13366_, _13364_);
  and (_13368_, _03872_, _02696_);
  nor (_13369_, _13368_, _07212_);
  or (_13370_, _07842_, _13369_);
  and (_13371_, _02959_, _02523_);
  and (_13372_, _02956_, _02523_);
  nor (_13373_, _13372_, _13371_);
  and (_13374_, _13373_, _03518_);
  and (_13375_, _13374_, _13370_);
  and (_13376_, _13375_, _13367_);
  and (_13377_, _02962_, _02523_);
  not (_13378_, _13369_);
  nor (_13379_, _13374_, _13378_);
  or (_13380_, _13379_, _13377_);
  or (_13381_, _13380_, _13376_);
  and (_13382_, _03014_, _02523_);
  not (_13383_, _13382_);
  nand (_13384_, _13378_, _13377_);
  and (_13385_, _13384_, _13383_);
  and (_13386_, _13385_, _13381_);
  and (_13387_, _13382_, _13249_);
  or (_13388_, _13387_, _03521_);
  or (_13389_, _13388_, _13386_);
  and (_13390_, _13389_, _13262_);
  or (_13392_, _13390_, _03146_);
  or (_13393_, _10369_, _03147_);
  and (_13394_, _13393_, _07861_);
  and (_13395_, _13394_, _13392_);
  and (_13396_, _07860_, _09272_);
  or (_13397_, _13396_, _03051_);
  or (_13398_, _13397_, _13395_);
  and (_13399_, _13398_, _13260_);
  or (_13400_, _13399_, _03148_);
  or (_13401_, _13257_, _07150_);
  and (_13403_, _13401_, _07882_);
  and (_13404_, _13403_, _13400_);
  or (_13405_, _13404_, _13256_);
  and (_13406_, _13405_, _07891_);
  and (_13407_, _07890_, _08051_);
  or (_13408_, _13407_, _03135_);
  or (_13409_, _13408_, _13406_);
  and (_13410_, _13409_, _13255_);
  and (_13411_, _08132_, _07311_);
  or (_13412_, _13411_, _13410_);
  and (_13414_, _13412_, _03023_);
  and (_13415_, _02855_, _02532_);
  or (_13416_, _13415_, _03757_);
  nor (_13417_, _13361_, _13293_);
  and (_13418_, _13417_, _03022_);
  or (_13419_, _13418_, _13416_);
  or (_13420_, _13419_, _13414_);
  and (_13421_, _02845_, _02532_);
  not (_13422_, _13421_);
  nand (_13423_, _13416_, _13368_);
  and (_13425_, _13423_, _13422_);
  and (_13426_, _13425_, _13420_);
  nor (_13427_, _13422_, _13368_);
  or (_13428_, _13427_, _07915_);
  or (_13429_, _13428_, _13426_);
  nand (_13430_, _07915_, _13248_);
  and (_13431_, _13430_, _03142_);
  and (_13432_, _13431_, _13429_);
  not (_13433_, _08812_);
  not (_13434_, _07921_);
  nand (_13436_, _10367_, _13434_);
  and (_13437_, _13436_, _13433_);
  or (_13438_, _13437_, _13432_);
  and (_13439_, _13438_, _13253_);
  nor (_13440_, _13439_, _03042_);
  nor (_13441_, _10365_, _07319_);
  nor (_13442_, _13441_, _13257_);
  and (_13443_, _13442_, _03042_);
  or (_13444_, _13443_, _07931_);
  nor (_13445_, _13444_, _13440_);
  or (_13447_, _07234_, _07521_);
  nand (_13448_, _13447_, _07936_);
  or (_13449_, _13448_, _13445_);
  nand (_13450_, _07229_, _07386_);
  and (_13451_, _13450_, _03134_);
  and (_13452_, _13451_, _13449_);
  nand (_13453_, _07997_, _07697_);
  and (_13454_, _13453_, _07966_);
  or (_13455_, _13454_, _13452_);
  and (_13456_, _13455_, _13252_);
  or (_13458_, _13456_, _07995_);
  nand (_13459_, _07995_, _07288_);
  and (_13460_, _13459_, _07189_);
  and (_13461_, _13460_, _13458_);
  and (_13462_, _03014_, _02509_);
  and (_13463_, _10153_, _13369_);
  or (_13464_, _13463_, _13462_);
  or (_13465_, _13464_, _13461_);
  nand (_13466_, _13462_, _13250_);
  and (_13467_, _13466_, _13465_);
  or (_13469_, _13467_, _03571_);
  and (_13470_, _13469_, _13251_);
  or (_13471_, _13470_, _02892_);
  nand (_13472_, _09290_, _02892_);
  and (_13473_, _13472_, _08117_);
  and (_13474_, _13473_, _13471_);
  and (_13475_, _08070_, _09272_);
  or (_13476_, _13475_, _08115_);
  or (_13477_, _13476_, _13474_);
  and (_13478_, _13477_, _13247_);
  or (_13480_, _13478_, _03174_);
  nand (_13481_, _13294_, _03174_);
  and (_13482_, _13481_, _08156_);
  and (_13483_, _13482_, _13480_);
  nor (_13484_, _08160_, _02696_);
  nor (_13485_, _13484_, _09732_);
  or (_13486_, _13485_, _13483_);
  nand (_13487_, _08160_, _02543_);
  and (_13488_, _13487_, _03183_);
  and (_13489_, _13488_, _13486_);
  and (_13491_, _13257_, _02799_);
  or (_13492_, _13491_, _02887_);
  or (_13493_, _13492_, _13489_);
  nand (_13494_, _13294_, _02887_);
  and (_13495_, _13494_, _08178_);
  and (_13496_, _13495_, _13493_);
  nor (_13497_, _08184_, _02696_);
  nor (_13498_, _13497_, _09755_);
  or (_13499_, _13498_, _13496_);
  nand (_13500_, _08184_, _02543_);
  and (_13502_, _13500_, _34655_);
  and (_13503_, _13502_, _13499_);
  or (_13504_, _13503_, _13246_);
  and (_35827_[0], _13504_, _35796_);
  nor (_13505_, _34655_, _02543_);
  nand (_13506_, _08115_, _02696_);
  nand (_13507_, _07921_, _07782_);
  nand (_13508_, _07210_, _07309_);
  or (_13509_, _07891_, _08048_);
  nor (_13510_, _04731_, _02543_);
  and (_13512_, _10689_, _04731_);
  nor (_13513_, _13512_, _13510_);
  nand (_13514_, _13513_, _03051_);
  nor (_13515_, _07319_, _04020_);
  nor (_13516_, _13515_, _13510_);
  nand (_13517_, _13516_, _05535_);
  nand (_13518_, _07403_, _04020_);
  nor (_13519_, _07595_, _03401_);
  or (_13520_, _07411_, _06163_);
  nor (_13521_, _07421_, _04020_);
  or (_13523_, _07423_, \oc8051_golden_model_1.ACC [1]);
  nand (_13524_, _07423_, \oc8051_golden_model_1.ACC [1]);
  and (_13525_, _13524_, _13523_);
  and (_13526_, _13525_, _07421_);
  or (_13527_, _13526_, _07410_);
  or (_13528_, _13527_, _13521_);
  and (_13529_, _13528_, _03401_);
  and (_13530_, _13529_, _13520_);
  or (_13531_, _13530_, _13519_);
  and (_13532_, _13531_, _07437_);
  and (_13534_, _07441_, xram_data_in_reg[1]);
  or (_13535_, _13534_, _03840_);
  or (_13536_, _13535_, _13532_);
  or (_13537_, _06163_, _05371_);
  and (_13538_, _13537_, _03006_);
  and (_13539_, _13538_, _13536_);
  nor (_13540_, _04731_, \oc8051_golden_model_1.ACC [1]);
  and (_13541_, _10574_, _04731_);
  nor (_13542_, _13541_, _13540_);
  and (_13543_, _13542_, _02948_);
  or (_13544_, _13543_, _07405_);
  or (_13545_, _13544_, _13539_);
  nor (_13546_, _07448_, \oc8051_golden_model_1.PSW [6]);
  and (_13547_, _13546_, \oc8051_golden_model_1.ACC [1]);
  nor (_13548_, _13546_, \oc8051_golden_model_1.ACC [1]);
  nor (_13549_, _13548_, _13547_);
  nand (_13550_, _13549_, _07405_);
  and (_13551_, _13550_, _02976_);
  and (_13552_, _13551_, _13545_);
  nor (_13553_, _05313_, _02543_);
  and (_13554_, _10569_, _05313_);
  nor (_13555_, _13554_, _13553_);
  nor (_13556_, _13555_, _02934_);
  nor (_13557_, _13516_, _07474_);
  or (_13558_, _13557_, _07403_);
  or (_13559_, _13558_, _13556_);
  or (_13560_, _13559_, _13552_);
  and (_13561_, _13560_, _13518_);
  or (_13562_, _13561_, _03873_);
  or (_13563_, _06163_, _07481_);
  and (_13564_, _13563_, _02992_);
  and (_13565_, _13564_, _13562_);
  nor (_13566_, _07595_, _02992_);
  or (_13567_, _13566_, _07485_);
  or (_13568_, _13567_, _13565_);
  nand (_13569_, _07485_, _06858_);
  and (_13570_, _13569_, _13568_);
  or (_13571_, _13570_, _02877_);
  and (_13572_, _10572_, _05313_);
  nor (_13573_, _13572_, _13553_);
  nand (_13574_, _13573_, _02877_);
  and (_13575_, _13574_, _06246_);
  and (_13576_, _13575_, _13571_);
  and (_13577_, _13554_, _10568_);
  nor (_13578_, _13577_, _13553_);
  nor (_13579_, _13578_, _06246_);
  or (_13580_, _13579_, _06252_);
  or (_13581_, _13580_, _13576_);
  and (_13582_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_13583_, _13582_, _07076_);
  nor (_13584_, _13583_, _06714_);
  or (_13585_, _13584_, _06258_);
  and (_13586_, _13585_, _13581_);
  or (_13587_, _13586_, _07400_);
  and (_13588_, _07784_, _03838_);
  nor (_13589_, _13588_, _07701_);
  and (_13590_, _13589_, _07211_);
  nor (_13591_, _13589_, _07211_);
  or (_13592_, _13591_, _13590_);
  and (_13593_, _13592_, _07507_);
  or (_13594_, _13593_, _09320_);
  and (_13595_, _13594_, _13587_);
  and (_13596_, _07784_, _06164_);
  nor (_13597_, _13596_, _07701_);
  and (_13598_, _13597_, _08050_);
  nor (_13599_, _13597_, _08050_);
  or (_13600_, _13599_, _13598_);
  and (_13601_, _13600_, _07397_);
  or (_13602_, _13601_, _02979_);
  or (_13603_, _13602_, _13595_);
  nand (_13604_, _07707_, _02979_);
  and (_13605_, _13604_, _07541_);
  and (_13606_, _13605_, _13603_);
  nor (_13607_, _07789_, _07541_);
  or (_13608_, _13607_, _07721_);
  or (_13609_, _13608_, _13606_);
  nand (_13610_, _03687_, _07721_);
  and (_13611_, _13610_, _02986_);
  and (_13612_, _13611_, _13609_);
  nor (_13613_, _10618_, _07806_);
  nor (_13614_, _13613_, _13553_);
  nor (_13615_, _13614_, _02986_);
  or (_13616_, _13615_, _05535_);
  or (_13617_, _13616_, _13612_);
  and (_13618_, _13617_, _13517_);
  or (_13619_, _13618_, _02841_);
  and (_13620_, _06163_, _04731_);
  nor (_13621_, _13620_, _13510_);
  nand (_13622_, _13621_, _02841_);
  and (_13623_, _13622_, _02839_);
  and (_13624_, _13623_, _13619_);
  and (_13625_, _10674_, _04731_);
  nor (_13626_, _13625_, _13510_);
  nor (_13627_, _13626_, _02839_);
  or (_13628_, _13627_, _06786_);
  or (_13629_, _13628_, _13624_);
  or (_13630_, _07042_, _06792_);
  and (_13631_, _13630_, _13629_);
  and (_13632_, _13631_, _02609_);
  nor (_13633_, _03687_, _02609_);
  or (_13634_, _13633_, _02834_);
  or (_13635_, _13634_, _13632_);
  and (_13636_, _04731_, _03720_);
  nor (_13637_, _13636_, _13540_);
  or (_13638_, _13637_, _07140_);
  and (_13639_, _13638_, _07831_);
  and (_13640_, _13639_, _13635_);
  nor (_13641_, _07831_, _03687_);
  or (_13642_, _13641_, _07843_);
  or (_13643_, _13642_, _13640_);
  or (_13644_, _13372_, _03517_);
  nor (_13645_, _13644_, _07843_);
  not (_13646_, _13644_);
  and (_13647_, _13646_, _07211_);
  or (_13648_, _13647_, _13645_);
  and (_13649_, _13648_, _13643_);
  and (_13650_, _02845_, _02523_);
  and (_13651_, _13644_, _07211_);
  or (_13652_, _13651_, _13650_);
  or (_13653_, _13652_, _13649_);
  not (_13654_, _13650_);
  or (_13655_, _13654_, _07211_);
  and (_13656_, _13655_, _07850_);
  and (_13657_, _13656_, _13653_);
  and (_13658_, _07849_, _08050_);
  or (_13659_, _13658_, _03146_);
  or (_13660_, _13659_, _13657_);
  or (_13661_, _10565_, _03147_);
  and (_13662_, _13661_, _07861_);
  and (_13663_, _13662_, _13660_);
  nor (_13664_, _07861_, _07783_);
  or (_13665_, _13664_, _03051_);
  or (_13666_, _13665_, _13663_);
  and (_13667_, _13666_, _13514_);
  or (_13668_, _13667_, _03148_);
  or (_13669_, _13510_, _07150_);
  and (_13670_, _13669_, _07875_);
  and (_13671_, _13670_, _13668_);
  and (_13672_, _07876_, _07209_);
  or (_13673_, _13672_, _03758_);
  or (_13674_, _13673_, _13671_);
  and (_13675_, _07888_, _07209_);
  or (_13676_, _13675_, _07881_);
  and (_13677_, _13676_, _13674_);
  and (_13678_, _07884_, _07209_);
  or (_13679_, _13678_, _07890_);
  or (_13680_, _13679_, _13677_);
  and (_13681_, _13680_, _13509_);
  or (_13682_, _13681_, _03135_);
  or (_13683_, _10563_, _03136_);
  and (_13684_, _13683_, _07312_);
  and (_13685_, _13684_, _13682_);
  and (_13686_, _07781_, _07311_);
  or (_13687_, _13686_, _13685_);
  and (_13688_, _13687_, _03023_);
  and (_13689_, _10688_, _04731_);
  nor (_13690_, _13689_, _13510_);
  nor (_13691_, _13690_, _03023_);
  or (_13692_, _13691_, _07309_);
  or (_13693_, _13692_, _13688_);
  and (_13694_, _13693_, _13508_);
  or (_13695_, _13694_, _07906_);
  nand (_13696_, _07906_, _07210_);
  and (_13697_, _13696_, _07913_);
  and (_13698_, _13697_, _13695_);
  nor (_13699_, _07210_, _07913_);
  or (_13700_, _13699_, _07915_);
  or (_13701_, _13700_, _13698_);
  nand (_13702_, _07915_, _08049_);
  and (_13703_, _13702_, _03142_);
  and (_13704_, _13703_, _13701_);
  nand (_13705_, _10564_, _13434_);
  and (_13706_, _13705_, _13433_);
  or (_13707_, _13706_, _13704_);
  and (_13708_, _13707_, _13507_);
  or (_13709_, _13708_, _03042_);
  nor (_13710_, _10687_, _07319_);
  or (_13711_, _13710_, _13510_);
  or (_13712_, _13711_, _03043_);
  and (_13713_, _13712_, _07234_);
  and (_13714_, _13713_, _13709_);
  and (_13715_, _07292_, _07287_);
  nor (_13716_, _13715_, _07293_);
  and (_13717_, _13716_, _07931_);
  or (_13718_, _13717_, _07229_);
  or (_13719_, _13718_, _13714_);
  and (_13720_, _07945_, _07384_);
  nor (_13721_, _13720_, _07946_);
  or (_13722_, _13721_, _07936_);
  and (_13723_, _13722_, _13719_);
  or (_13724_, _13723_, _03133_);
  and (_13725_, _07976_, _07974_);
  nor (_13726_, _13725_, _07977_);
  or (_13727_, _13726_, _03134_);
  and (_13728_, _13727_, _07997_);
  and (_13729_, _13728_, _13724_);
  and (_13730_, _08007_, _08005_);
  nor (_13731_, _13730_, _08008_);
  and (_13732_, _13731_, _07964_);
  or (_13733_, _13732_, _07995_);
  or (_13734_, _13733_, _13729_);
  nand (_13735_, _07995_, _02696_);
  and (_13736_, _13735_, _07189_);
  and (_13737_, _13736_, _13734_);
  or (_13738_, _07212_, _07211_);
  nor (_13739_, _07213_, _07189_);
  and (_13740_, _13739_, _13738_);
  or (_13741_, _13740_, _13737_);
  and (_13742_, _13741_, _08031_);
  or (_13743_, _08051_, _08050_);
  nor (_13744_, _08052_, _08031_);
  and (_13745_, _13744_, _13743_);
  or (_13746_, _13745_, _03359_);
  or (_13747_, _13746_, _13742_);
  and (_13748_, _08093_, _07700_);
  nor (_13749_, _13748_, _08094_);
  or (_13750_, _13749_, _03166_);
  and (_13751_, _13750_, _08117_);
  and (_13752_, _13751_, _13747_);
  and (_13753_, _07783_, _08133_);
  nor (_13754_, _13753_, _08134_);
  and (_13755_, _13754_, _08070_);
  or (_13756_, _13755_, _08115_);
  or (_13757_, _13756_, _13752_);
  and (_13758_, _13757_, _13506_);
  or (_13759_, _13758_, _03174_);
  or (_13760_, _13542_, _03179_);
  and (_13761_, _13760_, _08156_);
  and (_13762_, _13761_, _13759_);
  nor (_13763_, _08185_, _08161_);
  nor (_13764_, _13763_, _08156_);
  or (_13765_, _13764_, _08160_);
  or (_13766_, _13765_, _13762_);
  nand (_13767_, _08160_, _06964_);
  and (_13768_, _13767_, _03183_);
  and (_13769_, _13768_, _13766_);
  nor (_13770_, _13573_, _03183_);
  or (_13771_, _13770_, _02887_);
  or (_13772_, _13771_, _13769_);
  nor (_13773_, _13541_, _13510_);
  nand (_13774_, _13773_, _02887_);
  and (_13775_, _13774_, _08178_);
  and (_13776_, _13775_, _13772_);
  and (_13777_, _13763_, _08177_);
  or (_13778_, _13777_, _08184_);
  or (_13779_, _13778_, _13776_);
  nand (_13780_, _08184_, _06964_);
  and (_13781_, _13780_, _34655_);
  and (_13782_, _13781_, _13779_);
  or (_13783_, _13782_, _13505_);
  and (_35827_[1], _13783_, _35796_);
  nor (_13784_, _34655_, _06964_);
  nand (_13785_, _08115_, _02543_);
  and (_13786_, _08095_, _08090_);
  nor (_13787_, _13786_, _08096_);
  or (_13788_, _13787_, _03166_);
  and (_13789_, _13788_, _08117_);
  nand (_13790_, _07995_, _02543_);
  and (_13791_, _07978_, _07679_);
  nor (_13792_, _13791_, _07979_);
  or (_13793_, _13792_, _03134_);
  and (_13794_, _13793_, _07997_);
  nand (_13795_, _07206_, _07309_);
  nor (_13796_, _04731_, _06964_);
  and (_13797_, _10770_, _04731_);
  nor (_13798_, _13797_, _13796_);
  nand (_13799_, _13798_, _03051_);
  nand (_13800_, _13654_, _07842_);
  and (_13801_, _13800_, _07207_);
  nor (_13802_, _07831_, _03356_);
  nor (_13803_, _07319_, _04449_);
  nor (_13804_, _13803_, _13796_);
  nand (_13805_, _13804_, _05535_);
  nand (_13806_, _07403_, _04449_);
  nor (_13807_, _07577_, _03401_);
  or (_13808_, _07411_, _06167_);
  nor (_13809_, _07421_, _04449_);
  or (_13810_, _07423_, \oc8051_golden_model_1.ACC [2]);
  nand (_13811_, _07423_, \oc8051_golden_model_1.ACC [2]);
  and (_13812_, _13811_, _13810_);
  and (_13813_, _13812_, _07421_);
  or (_13814_, _13813_, _07410_);
  or (_13815_, _13814_, _13809_);
  and (_13816_, _13815_, _03401_);
  and (_13817_, _13816_, _13808_);
  or (_13818_, _13817_, _13807_);
  and (_13819_, _13818_, _07437_);
  and (_13820_, _07441_, xram_data_in_reg[2]);
  or (_13821_, _13820_, _03840_);
  or (_13822_, _13821_, _13819_);
  or (_13823_, _06167_, _05371_);
  and (_13824_, _13823_, _03006_);
  and (_13825_, _13824_, _13822_);
  nor (_13826_, _10788_, _07319_);
  nor (_13827_, _13826_, _13796_);
  nor (_13828_, _13827_, _03006_);
  or (_13829_, _13828_, _07405_);
  or (_13830_, _13829_, _13825_);
  nand (_13831_, _13546_, \oc8051_golden_model_1.ACC [2]);
  and (_13832_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_13833_, _13832_, _07447_);
  or (_13834_, _13833_, _13546_);
  and (_13835_, _13834_, _13831_);
  nand (_13836_, _13835_, _07405_);
  and (_13837_, _13836_, _02976_);
  and (_13838_, _13837_, _13830_);
  nor (_13839_, _05313_, _06964_);
  and (_13840_, _10792_, _05313_);
  nor (_13841_, _13840_, _13839_);
  nor (_13842_, _13841_, _02934_);
  nor (_13843_, _13804_, _07474_);
  or (_13844_, _13843_, _07403_);
  or (_13845_, _13844_, _13842_);
  or (_13846_, _13845_, _13838_);
  and (_13847_, _13846_, _13806_);
  or (_13848_, _13847_, _03873_);
  or (_13849_, _06167_, _07481_);
  and (_13850_, _13849_, _02992_);
  and (_13851_, _13850_, _13848_);
  nor (_13852_, _07577_, _02992_);
  or (_13853_, _13852_, _07485_);
  or (_13854_, _13853_, _13851_);
  nand (_13855_, _07485_, _06807_);
  and (_13856_, _13855_, _13854_);
  or (_13857_, _13856_, _02877_);
  and (_13858_, _10773_, _05313_);
  nor (_13859_, _13858_, _13839_);
  nand (_13860_, _13859_, _02877_);
  and (_13861_, _13860_, _06246_);
  and (_13862_, _13861_, _13857_);
  and (_13863_, _13840_, _10807_);
  nor (_13864_, _13863_, _13839_);
  nor (_13865_, _13864_, _06246_);
  or (_13866_, _13865_, _06252_);
  or (_13867_, _13866_, _13862_);
  nor (_13868_, _06716_, _06714_);
  nor (_13869_, _13868_, _06717_);
  or (_13870_, _13869_, _06258_);
  and (_13871_, _13870_, _13867_);
  or (_13872_, _13871_, _07400_);
  and (_13873_, _04020_, \oc8051_golden_model_1.ACC [1]);
  and (_13874_, _03838_, _02696_);
  nor (_13875_, _13874_, _07211_);
  nor (_13876_, _13875_, _13873_);
  nor (_13877_, _07207_, _13876_);
  and (_13878_, _07207_, _13876_);
  nor (_13879_, _13878_, _13877_);
  nor (_13880_, _13369_, _07211_);
  not (_13881_, _13880_);
  or (_13882_, _13881_, _13879_);
  and (_13883_, _13882_, \oc8051_golden_model_1.PSW [7]);
  nor (_13884_, _13879_, \oc8051_golden_model_1.PSW [7]);
  or (_13885_, _13884_, _13883_);
  nand (_13886_, _13881_, _13879_);
  and (_13887_, _13886_, _13885_);
  nor (_13888_, _13887_, _07397_);
  or (_13889_, _13888_, _09320_);
  and (_13890_, _13889_, _13872_);
  and (_13891_, _05900_, \oc8051_golden_model_1.ACC [1]);
  and (_13892_, _06164_, _02696_);
  nor (_13893_, _13892_, _08050_);
  nor (_13894_, _13893_, _13891_);
  nor (_13895_, _08046_, _13894_);
  and (_13896_, _08046_, _13894_);
  nor (_13897_, _13896_, _13895_);
  nor (_13898_, _13249_, _08050_);
  not (_13899_, _13898_);
  or (_13900_, _13899_, _13897_);
  and (_13901_, _13900_, \oc8051_golden_model_1.PSW [7]);
  nor (_13902_, _13897_, \oc8051_golden_model_1.PSW [7]);
  or (_13903_, _13902_, _13901_);
  nand (_13904_, _13899_, _13897_);
  and (_13905_, _13904_, _13903_);
  nor (_13906_, _13905_, _07507_);
  or (_13907_, _13906_, _02979_);
  or (_13908_, _13907_, _13890_);
  nor (_13909_, _09288_, _07698_);
  or (_13910_, _13909_, _07699_);
  and (_13911_, _08090_, _13910_);
  nor (_13912_, _08090_, _13910_);
  nor (_13913_, _13912_, _13911_);
  and (_13914_, _09291_, \oc8051_golden_model_1.PSW [7]);
  not (_13915_, _13914_);
  nor (_13916_, _13915_, _13913_);
  and (_13917_, _13915_, _13913_);
  nor (_13918_, _13917_, _13916_);
  nand (_13919_, _13918_, _02979_);
  and (_13920_, _13919_, _07541_);
  and (_13921_, _13920_, _13908_);
  and (_13922_, _02833_, _02696_);
  nor (_13923_, _09273_, _13922_);
  nor (_13924_, _13923_, _09821_);
  nor (_13925_, _08130_, _13924_);
  and (_13926_, _08130_, _13924_);
  nor (_13927_, _13926_, _13925_);
  not (_13928_, _09274_);
  or (_13929_, _13928_, _13927_);
  and (_13930_, _13929_, \oc8051_golden_model_1.PSW [7]);
  nor (_13931_, _13927_, \oc8051_golden_model_1.PSW [7]);
  or (_13932_, _13931_, _13930_);
  nand (_13933_, _13928_, _13927_);
  and (_13934_, _13933_, _13932_);
  nor (_13935_, _13934_, _07541_);
  or (_13936_, _13935_, _07721_);
  or (_13937_, _13936_, _13921_);
  nand (_13938_, _03356_, _07721_);
  and (_13939_, _13938_, _02986_);
  and (_13940_, _13939_, _13937_);
  nor (_13941_, _10825_, _07806_);
  nor (_13942_, _13941_, _13839_);
  nor (_13943_, _13942_, _02986_);
  or (_13944_, _13943_, _05535_);
  or (_13945_, _13944_, _13940_);
  and (_13946_, _13945_, _13805_);
  or (_13947_, _13946_, _02841_);
  and (_13948_, _06167_, _04731_);
  nor (_13949_, _13948_, _13796_);
  nand (_13950_, _13949_, _02841_);
  and (_13951_, _13950_, _02839_);
  and (_13952_, _13951_, _13947_);
  nor (_13953_, _10881_, _07319_);
  nor (_13954_, _13953_, _13796_);
  nor (_13955_, _13954_, _02839_);
  or (_13956_, _13955_, _06786_);
  or (_13957_, _13956_, _13952_);
  or (_13958_, _06978_, _06792_);
  and (_13959_, _13958_, _13957_);
  and (_13960_, _13959_, _02609_);
  nor (_13961_, _03356_, _02609_);
  or (_13962_, _13961_, _02834_);
  or (_13963_, _13962_, _13960_);
  and (_13964_, _04731_, _05693_);
  nor (_13965_, _13964_, _13796_);
  nand (_13966_, _13965_, _02834_);
  and (_13967_, _13966_, _07831_);
  and (_13968_, _13967_, _13963_);
  or (_13969_, _13968_, _13802_);
  and (_13970_, _13969_, _07842_);
  or (_13971_, _13970_, _13644_);
  or (_13972_, _13646_, _07207_);
  and (_13973_, _13972_, _13654_);
  and (_13974_, _13973_, _13971_);
  or (_13975_, _13974_, _13801_);
  and (_13976_, _13975_, _13383_);
  and (_13977_, _13382_, _08046_);
  or (_13978_, _13977_, _13976_);
  and (_13979_, _13978_, _13261_);
  and (_13980_, _08046_, _03521_);
  or (_13981_, _13980_, _03146_);
  or (_13982_, _13981_, _13979_);
  or (_13983_, _10766_, _03147_);
  and (_13984_, _13983_, _07861_);
  and (_13985_, _13984_, _13982_);
  and (_13986_, _07860_, _08130_);
  or (_13987_, _13986_, _03051_);
  or (_13988_, _13987_, _13985_);
  and (_13989_, _13988_, _13799_);
  or (_13990_, _13989_, _03148_);
  nor (_13991_, _02856_, _03528_);
  nor (_13992_, _13796_, _07150_);
  nor (_13993_, _13992_, _13991_);
  and (_13994_, _13993_, _13990_);
  nor (_13995_, _03019_, _03528_);
  nor (_13996_, _13991_, _13995_);
  not (_13997_, _13996_);
  or (_13998_, _13995_, _07205_);
  and (_13999_, _13998_, _13997_);
  or (_14000_, _13999_, _13994_);
  not (_14001_, _07205_);
  nand (_14002_, _13995_, _14001_);
  and (_14003_, _14002_, _03533_);
  and (_14004_, _14003_, _14000_);
  and (_14005_, _07205_, _03532_);
  or (_14006_, _14005_, _07890_);
  or (_14007_, _14006_, _14004_);
  or (_14008_, _07891_, _08044_);
  and (_14009_, _14008_, _03136_);
  and (_14010_, _14009_, _14007_);
  or (_14011_, _10764_, _07311_);
  and (_14012_, _14011_, _09456_);
  or (_14013_, _14012_, _14010_);
  or (_14014_, _08128_, _07312_);
  and (_14015_, _14014_, _03023_);
  and (_14016_, _14015_, _14013_);
  or (_14017_, _13965_, _10765_);
  nor (_14018_, _14017_, _03023_);
  or (_14019_, _14018_, _07309_);
  or (_14020_, _14019_, _14016_);
  and (_14021_, _14020_, _13795_);
  or (_14022_, _14021_, _07906_);
  nand (_14023_, _07906_, _07206_);
  and (_14024_, _14023_, _07913_);
  and (_14025_, _14024_, _14022_);
  nor (_14026_, _07206_, _07913_);
  or (_14027_, _14026_, _07915_);
  or (_14028_, _14027_, _14025_);
  nand (_14029_, _07915_, _08045_);
  and (_14030_, _14029_, _03142_);
  and (_14031_, _14030_, _14028_);
  nor (_14032_, _10765_, _03142_);
  or (_14033_, _14032_, _07921_);
  or (_14034_, _14033_, _14031_);
  nand (_14035_, _07921_, _08129_);
  and (_14036_, _14035_, _14034_);
  or (_14037_, _14036_, _03042_);
  nor (_14038_, _10768_, _07319_);
  nor (_14039_, _14038_, _13796_);
  nand (_14040_, _14039_, _03042_);
  and (_14041_, _14040_, _07234_);
  and (_14042_, _14041_, _14037_);
  and (_14043_, _07294_, _07280_);
  nor (_14044_, _14043_, _07295_);
  and (_14045_, _14044_, _07931_);
  or (_14046_, _14045_, _07229_);
  or (_14047_, _14046_, _14042_);
  and (_14048_, _07947_, _07366_);
  nor (_14049_, _14048_, _07948_);
  or (_14050_, _14049_, _07936_);
  and (_14051_, _14050_, _14047_);
  or (_14052_, _14051_, _03133_);
  and (_14053_, _14052_, _13794_);
  and (_14054_, _08009_, _07761_);
  nor (_14055_, _14054_, _08010_);
  and (_14056_, _14055_, _07964_);
  or (_14057_, _14056_, _07995_);
  or (_14058_, _14057_, _14053_);
  and (_14059_, _14058_, _13790_);
  or (_14060_, _14059_, _10153_);
  and (_14061_, _07214_, _07208_);
  nor (_14062_, _14061_, _07215_);
  or (_14063_, _14062_, _07189_);
  and (_14064_, _14063_, _08031_);
  and (_14065_, _14064_, _14060_);
  and (_14066_, _08053_, _08047_);
  nor (_14067_, _14066_, _08054_);
  and (_14068_, _14067_, _07185_);
  or (_14069_, _14068_, _03359_);
  or (_14070_, _14069_, _14065_);
  and (_14071_, _14070_, _13789_);
  and (_14072_, _08135_, _08131_);
  nor (_14073_, _14072_, _08136_);
  and (_14074_, _14073_, _08070_);
  or (_14075_, _14074_, _08115_);
  or (_14076_, _14075_, _14071_);
  and (_14077_, _14076_, _13785_);
  or (_14078_, _14077_, _03174_);
  nand (_14079_, _13827_, _03174_);
  and (_14080_, _14079_, _08156_);
  and (_14081_, _14080_, _14078_);
  and (_14082_, _07447_, _02696_);
  nor (_14083_, _08161_, _06964_);
  or (_14084_, _14083_, _14082_);
  and (_14085_, _14084_, _08155_);
  or (_14086_, _14085_, _08160_);
  or (_14087_, _14086_, _14081_);
  nand (_14088_, _08160_, _02625_);
  and (_14089_, _14088_, _03183_);
  and (_14090_, _14089_, _14087_);
  nor (_14091_, _13859_, _03183_);
  or (_14092_, _14091_, _02887_);
  or (_14093_, _14092_, _14090_);
  and (_14094_, _10941_, _04731_);
  nor (_14095_, _14094_, _13796_);
  nand (_14096_, _14095_, _02887_);
  and (_14097_, _14096_, _08178_);
  and (_14098_, _14097_, _14093_);
  and (_14099_, _08185_, \oc8051_golden_model_1.ACC [2]);
  nor (_14100_, _08185_, \oc8051_golden_model_1.ACC [2]);
  nor (_14101_, _14100_, _14099_);
  nor (_14102_, _14101_, _08184_);
  nor (_14103_, _14102_, _09755_);
  or (_14104_, _14103_, _14098_);
  nand (_14105_, _08184_, _02625_);
  and (_14106_, _14105_, _34655_);
  and (_14107_, _14106_, _14104_);
  or (_14108_, _14107_, _13784_);
  and (_35827_[2], _14108_, _35796_);
  nor (_14109_, _34655_, _02625_);
  and (_14110_, _07995_, \oc8051_golden_model_1.ACC [2]);
  and (_14111_, _07296_, _07274_);
  nor (_14112_, _14111_, _07297_);
  or (_14113_, _14112_, _07234_);
  or (_14114_, _07891_, _08042_);
  nor (_14115_, _04731_, _02625_);
  and (_14116_, _10968_, _04731_);
  nor (_14117_, _14116_, _14115_);
  nand (_14118_, _14117_, _03051_);
  and (_14119_, _07830_, _02794_);
  nor (_14120_, _07319_, _04275_);
  nor (_14121_, _14120_, _14115_);
  nand (_14122_, _14121_, _05535_);
  nor (_14123_, _05313_, _02625_);
  and (_14124_, _10976_, _05313_);
  and (_14125_, _14124_, _10975_);
  nor (_14126_, _14125_, _14123_);
  nor (_14127_, _14126_, _06246_);
  nand (_14128_, _07403_, _04275_);
  nor (_14129_, _07566_, _03401_);
  or (_14130_, _07411_, _06166_);
  nor (_14131_, _07421_, _04275_);
  or (_14132_, _07423_, \oc8051_golden_model_1.ACC [3]);
  nand (_14133_, _07423_, \oc8051_golden_model_1.ACC [3]);
  and (_14134_, _14133_, _14132_);
  and (_14135_, _14134_, _07421_);
  or (_14136_, _14135_, _07410_);
  or (_14137_, _14136_, _14131_);
  and (_14138_, _14137_, _03401_);
  and (_14139_, _14138_, _14130_);
  or (_14140_, _14139_, _14129_);
  and (_14141_, _14140_, _07437_);
  and (_14142_, _07441_, xram_data_in_reg[3]);
  or (_14143_, _14142_, _03840_);
  or (_14144_, _14143_, _14141_);
  or (_14145_, _06166_, _05371_);
  and (_14146_, _14145_, _03006_);
  and (_14147_, _14146_, _14144_);
  nor (_14148_, _10983_, _07319_);
  nor (_14149_, _14148_, _14115_);
  nor (_14150_, _14149_, _03006_);
  or (_14151_, _14150_, _07405_);
  or (_14152_, _14151_, _14147_);
  not (_14153_, \oc8051_golden_model_1.PSW [6]);
  nor (_14154_, _07447_, _14153_);
  nor (_14155_, _14154_, \oc8051_golden_model_1.ACC [3]);
  nor (_14156_, _14155_, _07448_);
  not (_14157_, _14156_);
  nand (_14158_, _14157_, _07405_);
  and (_14159_, _14158_, _02976_);
  and (_14160_, _14159_, _14152_);
  nor (_14161_, _14124_, _14123_);
  nor (_14162_, _14161_, _02934_);
  nor (_14163_, _14121_, _07474_);
  or (_14164_, _14163_, _07403_);
  or (_14165_, _14164_, _14162_);
  or (_14166_, _14165_, _14160_);
  and (_14167_, _14166_, _14128_);
  or (_14168_, _14167_, _03873_);
  or (_14169_, _06166_, _07481_);
  and (_14170_, _14169_, _02992_);
  and (_14171_, _14170_, _14168_);
  nor (_14172_, _07566_, _02992_);
  or (_14173_, _14172_, _07485_);
  or (_14174_, _14173_, _14171_);
  nand (_14175_, _07485_, _05364_);
  and (_14176_, _14175_, _14174_);
  or (_14177_, _14176_, _02877_);
  and (_14178_, _10979_, _05313_);
  nor (_14179_, _14178_, _14123_);
  nand (_14180_, _14179_, _02877_);
  and (_14181_, _14180_, _06246_);
  and (_14182_, _14181_, _14177_);
  or (_14183_, _14182_, _14127_);
  and (_14184_, _14183_, _06258_);
  nor (_14185_, _06719_, _06717_);
  nor (_14186_, _14185_, _06720_);
  and (_14187_, _14186_, _06252_);
  or (_14188_, _14187_, _07400_);
  or (_14189_, _14188_, _14184_);
  and (_14190_, _04449_, \oc8051_golden_model_1.ACC [2]);
  nor (_14191_, _13877_, _14190_);
  nor (_14192_, _07203_, _07204_);
  nor (_14193_, _14192_, _14191_);
  and (_14194_, _14192_, _14191_);
  nor (_14195_, _14194_, _14193_);
  and (_14196_, _14195_, \oc8051_golden_model_1.PSW [7]);
  nor (_14197_, _14195_, \oc8051_golden_model_1.PSW [7]);
  nor (_14198_, _14197_, _14196_);
  and (_14199_, _14198_, _13883_);
  nor (_14200_, _14198_, _13883_);
  or (_14201_, _14200_, _14199_);
  nand (_14202_, _14201_, _07400_);
  and (_14203_, _14202_, _14189_);
  or (_14204_, _14203_, _07397_);
  and (_14205_, _06036_, \oc8051_golden_model_1.ACC [2]);
  nor (_14206_, _13895_, _14205_);
  nor (_14207_, _08042_, _08043_);
  nor (_14208_, _14207_, _14206_);
  and (_14209_, _14207_, _14206_);
  nor (_14210_, _14209_, _14208_);
  and (_14211_, _14210_, \oc8051_golden_model_1.PSW [7]);
  nor (_14212_, _14210_, \oc8051_golden_model_1.PSW [7]);
  nor (_14213_, _14212_, _14211_);
  and (_14214_, _14213_, _13901_);
  nor (_14215_, _14213_, _13901_);
  or (_14216_, _14215_, _14214_);
  nand (_14217_, _14216_, _07397_);
  and (_14218_, _14217_, _02991_);
  and (_14219_, _14218_, _14204_);
  and (_14220_, _09292_, \oc8051_golden_model_1.PSW [7]);
  nor (_14221_, _13911_, _08088_);
  not (_14222_, _09286_);
  and (_14223_, _14222_, _14221_);
  nor (_14224_, _14222_, _14221_);
  nor (_14225_, _14224_, _14223_);
  not (_14226_, _13916_);
  and (_14227_, _14226_, _14225_);
  nor (_14228_, _14227_, _14220_);
  nand (_14229_, _14228_, _07541_);
  and (_14230_, _14229_, _09325_);
  or (_14231_, _14230_, _14219_);
  and (_14232_, _03356_, \oc8051_golden_model_1.ACC [2]);
  nor (_14233_, _13925_, _14232_);
  nor (_14234_, _09269_, _14233_);
  and (_14235_, _09269_, _14233_);
  nor (_14236_, _14235_, _14234_);
  and (_14237_, _14236_, \oc8051_golden_model_1.PSW [7]);
  nor (_14238_, _14236_, \oc8051_golden_model_1.PSW [7]);
  nor (_14239_, _14238_, _14237_);
  and (_14240_, _14239_, _13930_);
  nor (_14241_, _14239_, _13930_);
  nor (_14242_, _14241_, _14240_);
  or (_14243_, _14242_, _07541_);
  and (_14244_, _14243_, _14231_);
  or (_14245_, _14244_, _07721_);
  or (_14246_, _02794_, _02571_);
  and (_14247_, _14246_, _02986_);
  and (_14248_, _14247_, _14245_);
  nor (_14249_, _10973_, _07806_);
  nor (_14250_, _14249_, _14123_);
  nor (_14251_, _14250_, _02986_);
  or (_14252_, _14251_, _05535_);
  or (_14253_, _14252_, _14248_);
  and (_14254_, _14253_, _14122_);
  or (_14255_, _14254_, _02841_);
  and (_14256_, _06166_, _04731_);
  nor (_14257_, _14256_, _14115_);
  nand (_14258_, _14257_, _02841_);
  and (_14259_, _14258_, _02839_);
  and (_14260_, _14259_, _14255_);
  nor (_14261_, _11076_, _07319_);
  nor (_14262_, _14261_, _14115_);
  nor (_14263_, _14262_, _02839_);
  or (_14264_, _14263_, _06786_);
  or (_14265_, _14264_, _14260_);
  or (_14266_, _06925_, _06792_);
  and (_14267_, _14266_, _14265_);
  and (_14268_, _14267_, _02609_);
  and (_14269_, _02794_, _02542_);
  or (_14270_, _14269_, _02834_);
  or (_14271_, _14270_, _14268_);
  and (_14272_, _04731_, _05654_);
  nor (_14273_, _14272_, _14115_);
  nand (_14274_, _14273_, _02834_);
  and (_14275_, _14274_, _07831_);
  and (_14276_, _14275_, _14271_);
  or (_14277_, _14276_, _14119_);
  and (_14278_, _14277_, _07845_);
  and (_14279_, _07846_, _14192_);
  or (_14280_, _14279_, _14278_);
  and (_14281_, _14280_, _07850_);
  and (_14282_, _07849_, _14207_);
  or (_14283_, _14282_, _03146_);
  or (_14284_, _14283_, _14281_);
  or (_14285_, _10964_, _03147_);
  and (_14286_, _14285_, _07861_);
  and (_14287_, _14286_, _14284_);
  and (_14288_, _07860_, _09269_);
  or (_14289_, _14288_, _03051_);
  or (_14290_, _14289_, _14287_);
  and (_14291_, _14290_, _14118_);
  or (_14292_, _14291_, _03148_);
  or (_14293_, _14115_, _07150_);
  and (_14294_, _14293_, _07882_);
  and (_14295_, _14294_, _14292_);
  and (_14296_, _07883_, _07203_);
  or (_14297_, _14296_, _07890_);
  or (_14298_, _14297_, _14295_);
  and (_14299_, _14298_, _14114_);
  or (_14300_, _14299_, _03135_);
  or (_14301_, _10963_, _03136_);
  and (_14302_, _14301_, _07312_);
  and (_14303_, _14302_, _14300_);
  and (_14304_, _08126_, _07311_);
  or (_14305_, _14304_, _14303_);
  and (_14306_, _14305_, _03023_);
  or (_14307_, _14273_, _10962_);
  nor (_14308_, _14307_, _03023_);
  or (_14309_, _14308_, _09468_);
  or (_14310_, _14309_, _14306_);
  nand (_14311_, _07915_, _08043_);
  not (_14312_, _08814_);
  nand (_14313_, _14312_, _07204_);
  and (_14314_, _14313_, _03142_);
  and (_14315_, _14314_, _14311_);
  and (_14316_, _14315_, _14310_);
  nand (_14317_, _10962_, _13434_);
  and (_14318_, _14317_, _13433_);
  or (_14319_, _14318_, _14316_);
  nand (_14320_, _07921_, _08127_);
  and (_14321_, _14320_, _03043_);
  and (_14322_, _14321_, _14319_);
  nor (_14323_, _10967_, _07319_);
  nor (_14324_, _14323_, _14115_);
  nor (_14325_, _14324_, _03043_);
  or (_14326_, _14325_, _07931_);
  or (_14327_, _14326_, _14322_);
  and (_14328_, _14327_, _14113_);
  or (_14329_, _14328_, _07229_);
  and (_14330_, _07949_, _07361_);
  nor (_14331_, _14330_, _07950_);
  or (_14332_, _14331_, _07936_);
  and (_14333_, _14332_, _03134_);
  and (_14334_, _14333_, _14329_);
  and (_14335_, _07980_, _07674_);
  nor (_14336_, _14335_, _07981_);
  or (_14337_, _14336_, _07964_);
  and (_14338_, _14337_, _07966_);
  or (_14339_, _14338_, _14334_);
  and (_14340_, _08011_, _07756_);
  nor (_14341_, _14340_, _08012_);
  or (_14342_, _14341_, _07997_);
  and (_14343_, _14342_, _07996_);
  and (_14344_, _14343_, _14339_);
  or (_14345_, _14344_, _14110_);
  and (_14346_, _14345_, _07189_);
  nor (_14347_, _07216_, _14192_);
  and (_14348_, _07216_, _14192_);
  nor (_14349_, _14348_, _14347_);
  nor (_14350_, _14349_, _07189_);
  or (_14351_, _14350_, _07185_);
  or (_14352_, _14351_, _14346_);
  nor (_14353_, _08055_, _14207_);
  and (_14354_, _08055_, _14207_);
  nor (_14355_, _14354_, _14353_);
  nand (_14356_, _14355_, _07185_);
  and (_14357_, _14356_, _03166_);
  and (_14358_, _14357_, _14352_);
  and (_14359_, _08097_, _14222_);
  nor (_14360_, _08097_, _14222_);
  nor (_14361_, _14360_, _14359_);
  nand (_14362_, _14361_, _04138_);
  and (_14363_, _14362_, _08112_);
  or (_14364_, _14363_, _14358_);
  nor (_14365_, _08137_, _09269_);
  and (_14366_, _08137_, _09269_);
  nor (_14367_, _14366_, _14365_);
  nand (_14368_, _14367_, _08070_);
  and (_14369_, _14368_, _08116_);
  and (_14370_, _14369_, _14364_);
  and (_14371_, _08115_, \oc8051_golden_model_1.ACC [2]);
  or (_14372_, _14371_, _03174_);
  or (_14373_, _14372_, _14370_);
  nand (_14374_, _14149_, _03174_);
  and (_14375_, _14374_, _08156_);
  and (_14376_, _14375_, _14373_);
  nor (_14377_, _14082_, _02625_);
  or (_14378_, _14377_, _08162_);
  and (_14379_, _14378_, _08155_);
  or (_14380_, _14379_, _08160_);
  or (_14381_, _14380_, _14376_);
  nand (_14382_, _08160_, _06864_);
  and (_14383_, _14382_, _03183_);
  and (_14384_, _14383_, _14381_);
  nor (_14385_, _14179_, _03183_);
  or (_14386_, _14385_, _02887_);
  or (_14387_, _14386_, _14384_);
  and (_14388_, _11136_, _04731_);
  nor (_14389_, _14388_, _14115_);
  nand (_14390_, _14389_, _02887_);
  and (_14391_, _14390_, _08178_);
  and (_14392_, _14391_, _14387_);
  or (_14393_, _14099_, \oc8051_golden_model_1.ACC [3]);
  and (_14394_, _14393_, _08186_);
  and (_14395_, _14394_, _08177_);
  or (_14396_, _14395_, _08184_);
  or (_14397_, _14396_, _14392_);
  nand (_14398_, _08184_, _06864_);
  and (_14399_, _14398_, _34655_);
  and (_14400_, _14399_, _14397_);
  or (_14401_, _14400_, _14109_);
  and (_35827_[3], _14401_, _35796_);
  nor (_14402_, _34655_, _06864_);
  nand (_14403_, _07995_, _02625_);
  nand (_14404_, _07201_, _07309_);
  nor (_14405_, _04731_, _06864_);
  and (_14406_, _11158_, _04731_);
  nor (_14407_, _14406_, _14405_);
  nand (_14408_, _14407_, _03051_);
  and (_14409_, _13800_, _07202_);
  nor (_14410_, _07831_, _03647_);
  nor (_14411_, _05192_, _07319_);
  nor (_14412_, _14411_, _14405_);
  nand (_14413_, _14412_, _05535_);
  nor (_14414_, _14221_, _09284_);
  or (_14415_, _14414_, _09285_);
  and (_14416_, _08085_, _14415_);
  nor (_14417_, _08085_, _14415_);
  nor (_14418_, _14417_, _14416_);
  not (_14419_, _14220_);
  nor (_14420_, _14419_, _14418_);
  and (_14421_, _14419_, _14418_);
  nor (_14422_, _14421_, _14420_);
  nand (_14423_, _14422_, _02979_);
  and (_14424_, _14423_, _07541_);
  nor (_14425_, _11184_, _07319_);
  nor (_14426_, _14425_, _14405_);
  nand (_14427_, _14426_, _02948_);
  nor (_14428_, _07638_, _03401_);
  or (_14429_, _07411_, _06171_);
  nor (_14430_, _07421_, _05192_);
  or (_14431_, _07423_, \oc8051_golden_model_1.ACC [4]);
  nand (_14432_, _07423_, \oc8051_golden_model_1.ACC [4]);
  and (_14433_, _14432_, _14431_);
  and (_14434_, _14433_, _07421_);
  or (_14435_, _14434_, _07410_);
  or (_14436_, _14435_, _14430_);
  and (_14437_, _14436_, _03401_);
  and (_14438_, _14437_, _14429_);
  or (_14439_, _14438_, _14428_);
  and (_14440_, _14439_, _07437_);
  and (_14441_, _07441_, xram_data_in_reg[4]);
  or (_14442_, _14441_, _02948_);
  or (_14443_, _14442_, _14440_);
  and (_14444_, _14443_, _14427_);
  or (_14445_, _14444_, _07405_);
  nor (_14446_, _07448_, \oc8051_golden_model_1.ACC [4]);
  nor (_14447_, _14446_, _07454_);
  not (_14448_, _14447_);
  nand (_14449_, _14448_, _07405_);
  and (_14450_, _14449_, _02976_);
  and (_14451_, _14450_, _14445_);
  nor (_14452_, _05313_, _06864_);
  and (_14453_, _11167_, _05313_);
  nor (_14454_, _14453_, _14452_);
  nor (_14455_, _14454_, _02934_);
  nor (_14456_, _14412_, _07474_);
  or (_14457_, _14456_, _07403_);
  or (_14458_, _14457_, _14455_);
  or (_14459_, _14458_, _14451_);
  nand (_14460_, _07403_, _05192_);
  and (_14461_, _14460_, _14459_);
  or (_14462_, _14461_, _03873_);
  or (_14463_, _06171_, _07481_);
  and (_14464_, _14463_, _02992_);
  and (_14465_, _14464_, _14462_);
  nor (_14466_, _07638_, _02992_);
  or (_14467_, _14466_, _07485_);
  or (_14468_, _14467_, _14465_);
  nand (_14469_, _07485_, _02696_);
  and (_14470_, _14469_, _14468_);
  or (_14471_, _14470_, _02877_);
  and (_14472_, _11165_, _05313_);
  nor (_14473_, _14472_, _14452_);
  nand (_14474_, _14473_, _02877_);
  and (_14475_, _14474_, _06246_);
  and (_14476_, _14475_, _14471_);
  and (_14477_, _14453_, _11201_);
  nor (_14478_, _14477_, _14452_);
  nor (_14479_, _14478_, _06246_);
  or (_14480_, _14479_, _06252_);
  or (_14481_, _14480_, _14476_);
  nor (_14482_, _06722_, _06720_);
  nor (_14483_, _14482_, _06723_);
  or (_14484_, _14483_, _06258_);
  and (_14485_, _14484_, _14481_);
  or (_14486_, _14485_, _07400_);
  or (_14487_, _14199_, _14196_);
  nor (_14488_, _04275_, \oc8051_golden_model_1.ACC [3]);
  nand (_14489_, _04275_, \oc8051_golden_model_1.ACC [3]);
  and (_14490_, _14489_, _14191_);
  or (_14491_, _14490_, _14488_);
  nor (_14492_, _07202_, _14491_);
  and (_14493_, _07202_, _14491_);
  nor (_14494_, _14493_, _14492_);
  and (_14495_, _14494_, \oc8051_golden_model_1.PSW [7]);
  nor (_14496_, _14494_, \oc8051_golden_model_1.PSW [7]);
  nor (_14497_, _14496_, _14495_);
  and (_14498_, _14497_, _14487_);
  nor (_14499_, _14497_, _14487_);
  nor (_14500_, _14499_, _14498_);
  and (_14501_, _14500_, _07507_);
  or (_14502_, _14501_, _09320_);
  and (_14503_, _14502_, _14486_);
  or (_14504_, _14214_, _14211_);
  and (_14505_, _06166_, _02625_);
  or (_14506_, _06166_, _02625_);
  and (_14507_, _14506_, _14206_);
  or (_14508_, _14507_, _14505_);
  nor (_14509_, _08041_, _14508_);
  and (_14510_, _08041_, _14508_);
  nor (_14511_, _14510_, _14509_);
  and (_14512_, _14511_, \oc8051_golden_model_1.PSW [7]);
  nor (_14513_, _14511_, \oc8051_golden_model_1.PSW [7]);
  nor (_14514_, _14513_, _14512_);
  and (_14515_, _14514_, _14504_);
  nor (_14516_, _14514_, _14504_);
  nor (_14517_, _14516_, _14515_);
  and (_14518_, _14517_, _07397_);
  or (_14519_, _14518_, _02979_);
  or (_14520_, _14519_, _14503_);
  and (_14521_, _14520_, _14424_);
  or (_14522_, _14240_, _14237_);
  nor (_14523_, _14233_, _09827_);
  nor (_14524_, _14523_, _09826_);
  nor (_14525_, _08125_, _14524_);
  and (_14526_, _08125_, _14524_);
  nor (_14527_, _14526_, _14525_);
  and (_14528_, _14527_, \oc8051_golden_model_1.PSW [7]);
  nor (_14529_, _14527_, \oc8051_golden_model_1.PSW [7]);
  nor (_14530_, _14529_, _14528_);
  and (_14531_, _14530_, _14522_);
  nor (_14532_, _14530_, _14522_);
  nor (_14533_, _14532_, _14531_);
  and (_14534_, _14533_, _07540_);
  or (_14535_, _14534_, _07721_);
  or (_14536_, _14535_, _14521_);
  nand (_14537_, _03647_, _07721_);
  and (_14538_, _14537_, _02986_);
  and (_14539_, _14538_, _14536_);
  nor (_14540_, _11163_, _07806_);
  nor (_14541_, _14540_, _14452_);
  nor (_14542_, _14541_, _02986_);
  or (_14543_, _14542_, _05535_);
  or (_14544_, _14543_, _14539_);
  and (_14545_, _14544_, _14413_);
  or (_14546_, _14545_, _02841_);
  and (_14547_, _06171_, _04731_);
  nor (_14548_, _14547_, _14405_);
  nand (_14549_, _14548_, _02841_);
  and (_14550_, _14549_, _02839_);
  and (_14551_, _14550_, _14546_);
  nor (_14552_, _11271_, _07319_);
  nor (_14553_, _14552_, _14405_);
  nor (_14554_, _14553_, _02839_);
  or (_14555_, _14554_, _06786_);
  or (_14556_, _14555_, _14551_);
  or (_14557_, _06872_, _06792_);
  and (_14558_, _14557_, _14556_);
  and (_14559_, _14558_, _02609_);
  nor (_14560_, _03647_, _02609_);
  or (_14561_, _14560_, _02834_);
  or (_14562_, _14561_, _14559_);
  and (_14563_, _05618_, _04731_);
  nor (_14564_, _14563_, _14405_);
  nand (_14565_, _14564_, _02834_);
  and (_14566_, _14565_, _07831_);
  and (_14567_, _14566_, _14562_);
  or (_14568_, _14567_, _14410_);
  and (_14569_, _14568_, _07842_);
  or (_14570_, _14569_, _13644_);
  or (_14571_, _13646_, _07202_);
  and (_14572_, _14571_, _13654_);
  and (_14573_, _14572_, _14570_);
  or (_14574_, _14573_, _14409_);
  and (_14575_, _14574_, _13383_);
  and (_14576_, _13382_, _08041_);
  or (_14577_, _14576_, _14575_);
  and (_14578_, _14577_, _13261_);
  and (_14579_, _08041_, _03521_);
  or (_14580_, _14579_, _03146_);
  or (_14581_, _14580_, _14578_);
  or (_14582_, _11154_, _03147_);
  and (_14583_, _14582_, _07861_);
  and (_14584_, _14583_, _14581_);
  and (_14585_, _07860_, _08125_);
  or (_14586_, _14585_, _03051_);
  or (_14587_, _14586_, _14584_);
  and (_14588_, _14587_, _14408_);
  or (_14589_, _14588_, _03148_);
  or (_14590_, _14405_, _07150_);
  and (_14591_, _14590_, _13996_);
  and (_14592_, _14591_, _14589_);
  and (_14593_, _13997_, _07200_);
  or (_14594_, _14593_, _03532_);
  or (_14595_, _14594_, _14592_);
  or (_14596_, _07200_, _03533_);
  and (_14597_, _14596_, _07891_);
  and (_14598_, _14597_, _14595_);
  and (_14599_, _07890_, _08039_);
  or (_14600_, _14599_, _03135_);
  or (_14601_, _14600_, _14598_);
  or (_14602_, _11153_, _03136_);
  and (_14603_, _14602_, _07312_);
  and (_14604_, _14603_, _14601_);
  and (_14605_, _08123_, _07311_);
  or (_14606_, _14605_, _14604_);
  and (_14607_, _14606_, _03023_);
  or (_14608_, _14564_, _11152_);
  nor (_14609_, _14608_, _03023_);
  or (_14610_, _14609_, _07309_);
  or (_14611_, _14610_, _14607_);
  and (_14612_, _14611_, _14404_);
  or (_14613_, _14612_, _07906_);
  nand (_14614_, _07906_, _07201_);
  and (_14615_, _14614_, _07913_);
  and (_14616_, _14615_, _14613_);
  nor (_14617_, _07201_, _07913_);
  or (_14618_, _14617_, _07915_);
  or (_14619_, _14618_, _14616_);
  nand (_14620_, _07915_, _08040_);
  and (_14621_, _14620_, _03142_);
  and (_14622_, _14621_, _14619_);
  nor (_14623_, _11152_, _03142_);
  or (_14624_, _14623_, _07921_);
  or (_14625_, _14624_, _14622_);
  nand (_14626_, _07921_, _08124_);
  and (_14627_, _14626_, _14625_);
  or (_14628_, _14627_, _03042_);
  nor (_14629_, _11157_, _07319_);
  nor (_14630_, _14629_, _14405_);
  nand (_14631_, _14630_, _03042_);
  and (_14632_, _14631_, _07234_);
  and (_14633_, _14632_, _14628_);
  and (_14634_, _07298_, _07265_);
  nor (_14635_, _14634_, _07299_);
  and (_14636_, _14635_, _07931_);
  or (_14637_, _14636_, _14633_);
  and (_14638_, _14637_, _07936_);
  and (_14639_, _07951_, _07352_);
  nor (_14640_, _14639_, _07952_);
  and (_14641_, _14640_, _07229_);
  or (_14642_, _14641_, _03133_);
  or (_14643_, _14642_, _14638_);
  and (_14644_, _07982_, _07667_);
  nor (_14645_, _14644_, _07983_);
  or (_14646_, _14645_, _03134_);
  and (_14647_, _14646_, _07997_);
  and (_14648_, _14647_, _14643_);
  and (_14649_, _08013_, _07749_);
  nor (_14650_, _14649_, _08014_);
  and (_14651_, _14650_, _07964_);
  or (_14652_, _14651_, _07995_);
  or (_14653_, _14652_, _14648_);
  and (_14654_, _14653_, _14403_);
  or (_14655_, _14654_, _10153_);
  nor (_14656_, _07218_, _07202_);
  nor (_14657_, _14656_, _07219_);
  or (_14658_, _14657_, _07189_);
  and (_14659_, _14658_, _08031_);
  and (_14660_, _14659_, _14655_);
  nor (_14661_, _08057_, _08041_);
  nor (_14662_, _14661_, _08058_);
  and (_14663_, _14662_, _07185_);
  or (_14664_, _14663_, _08112_);
  or (_14665_, _14664_, _14660_);
  nor (_14666_, _08101_, _08086_);
  nor (_14667_, _14666_, _08102_);
  or (_14668_, _14667_, _10168_);
  nor (_14669_, _08139_, _08125_);
  nor (_14670_, _14669_, _08140_);
  or (_14671_, _14670_, _08117_);
  and (_14672_, _14671_, _08116_);
  and (_14673_, _14672_, _14668_);
  and (_14674_, _14673_, _14665_);
  and (_14675_, _08115_, \oc8051_golden_model_1.ACC [3]);
  or (_14676_, _14675_, _03174_);
  or (_14677_, _14676_, _14674_);
  nand (_14678_, _14426_, _03174_);
  and (_14679_, _14678_, _08156_);
  and (_14680_, _14679_, _14677_);
  and (_14681_, _08162_, _06864_);
  nor (_14682_, _08162_, _06864_);
  nor (_14683_, _14682_, _14681_);
  not (_14684_, _14683_);
  nor (_14685_, _14684_, _08160_);
  nor (_14686_, _14685_, _09732_);
  or (_14687_, _14686_, _14680_);
  nand (_14688_, _08160_, _06858_);
  and (_14689_, _14688_, _03183_);
  and (_14690_, _14689_, _14687_);
  nor (_14691_, _14473_, _03183_);
  or (_14692_, _14691_, _02887_);
  or (_14693_, _14692_, _14690_);
  and (_14694_, _11338_, _04731_);
  nor (_14695_, _14694_, _14405_);
  nand (_14696_, _14695_, _02887_);
  and (_14697_, _14696_, _08178_);
  and (_14698_, _14697_, _14693_);
  and (_14699_, _08186_, _06864_);
  nor (_14700_, _14699_, _08187_);
  and (_14701_, _14700_, _08177_);
  or (_14702_, _14701_, _08184_);
  or (_14703_, _14702_, _14698_);
  nand (_14704_, _08184_, _06858_);
  and (_14705_, _14704_, _34655_);
  and (_14706_, _14705_, _14703_);
  or (_14707_, _14706_, _14402_);
  and (_35827_[4], _14707_, _35796_);
  nor (_14708_, _34655_, _06858_);
  and (_14709_, _07220_, _07199_);
  nor (_14710_, _14709_, _07221_);
  or (_14711_, _14710_, _07189_);
  and (_14712_, _07300_, _07257_);
  nor (_14713_, _14712_, _07301_);
  or (_14714_, _14713_, _07234_);
  nor (_14715_, _07416_, _03543_);
  and (_14716_, _07883_, _07196_);
  nor (_14717_, _04731_, _06858_);
  and (_14718_, _11482_, _04731_);
  nor (_14719_, _14718_, _14717_);
  nand (_14720_, _14719_, _03051_);
  or (_14721_, _08037_, _13261_);
  nor (_14722_, _07831_, _03220_);
  nor (_14723_, _04894_, _07319_);
  nor (_14724_, _14723_, _14717_);
  nand (_14725_, _14724_, _05535_);
  and (_14726_, _03647_, \oc8051_golden_model_1.ACC [4]);
  nor (_14727_, _14525_, _14726_);
  nor (_14728_, _09265_, _14727_);
  and (_14729_, _09265_, _14727_);
  nor (_14730_, _14729_, _14728_);
  and (_14731_, _14730_, \oc8051_golden_model_1.PSW [7]);
  nor (_14732_, _14730_, \oc8051_golden_model_1.PSW [7]);
  nor (_14733_, _14732_, _14731_);
  nor (_14734_, _14531_, _14528_);
  not (_14735_, _14734_);
  and (_14736_, _14735_, _14733_);
  nor (_14737_, _14735_, _14733_);
  nor (_14738_, _14737_, _14736_);
  or (_14739_, _14738_, _07541_);
  nor (_14740_, _05313_, _06858_);
  and (_14741_, _11365_, _05313_);
  and (_14742_, _14741_, _11397_);
  nor (_14743_, _14742_, _14740_);
  nor (_14744_, _14743_, _06246_);
  nor (_14745_, _11380_, _07319_);
  nor (_14746_, _14745_, _14717_);
  nand (_14747_, _14746_, _02948_);
  nor (_14748_, _07621_, _03401_);
  or (_14749_, _07411_, _06170_);
  nor (_14750_, _07421_, _04894_);
  or (_14751_, _07423_, \oc8051_golden_model_1.ACC [5]);
  nand (_14752_, _07423_, \oc8051_golden_model_1.ACC [5]);
  and (_14753_, _14752_, _14751_);
  and (_14754_, _14753_, _07421_);
  or (_14755_, _14754_, _07410_);
  or (_14756_, _14755_, _14750_);
  and (_14757_, _14756_, _03401_);
  and (_14758_, _14757_, _14749_);
  or (_14759_, _14758_, _14748_);
  and (_14760_, _14759_, _07437_);
  and (_14761_, _07441_, xram_data_in_reg[5]);
  or (_14762_, _14761_, _02948_);
  or (_14763_, _14762_, _14760_);
  and (_14764_, _14763_, _14747_);
  or (_14765_, _14764_, _07405_);
  and (_14766_, _09862_, _07456_);
  nor (_14767_, _09862_, _07456_);
  nor (_14768_, _14767_, _14766_);
  nand (_14769_, _14768_, _07405_);
  and (_14770_, _14769_, _02976_);
  and (_14771_, _14770_, _14765_);
  nor (_14772_, _14741_, _14740_);
  nor (_14773_, _14772_, _02934_);
  nor (_14774_, _14724_, _07474_);
  or (_14775_, _14774_, _07403_);
  or (_14776_, _14775_, _14773_);
  or (_14777_, _14776_, _14771_);
  nand (_14778_, _07403_, _04894_);
  and (_14779_, _14778_, _14777_);
  or (_14780_, _14779_, _03873_);
  or (_14781_, _06170_, _07481_);
  and (_14782_, _14781_, _02992_);
  and (_14783_, _14782_, _14780_);
  nor (_14784_, _07621_, _02992_);
  or (_14785_, _14784_, _07485_);
  or (_14786_, _14785_, _14783_);
  nand (_14787_, _07485_, _02543_);
  and (_14788_, _14787_, _14786_);
  or (_14789_, _14788_, _02877_);
  and (_14790_, _11363_, _05313_);
  nor (_14791_, _14790_, _14740_);
  nand (_14792_, _14791_, _02877_);
  and (_14793_, _14792_, _06246_);
  and (_14794_, _14793_, _14789_);
  or (_14795_, _14794_, _14744_);
  and (_14796_, _14795_, _06258_);
  nor (_14797_, _06725_, _06723_);
  nor (_14798_, _14797_, _06726_);
  and (_14799_, _14798_, _06252_);
  or (_14800_, _14799_, _07400_);
  or (_14801_, _14800_, _14796_);
  and (_14802_, _05192_, \oc8051_golden_model_1.ACC [4]);
  nor (_14803_, _14492_, _14802_);
  nor (_14804_, _07198_, _14803_);
  and (_14805_, _07198_, _14803_);
  nor (_14806_, _14805_, _14804_);
  and (_14807_, _14806_, \oc8051_golden_model_1.PSW [7]);
  nor (_14808_, _14806_, \oc8051_golden_model_1.PSW [7]);
  nor (_14809_, _14808_, _14807_);
  nor (_14810_, _14498_, _14495_);
  not (_14811_, _14810_);
  and (_14812_, _14811_, _14809_);
  nor (_14813_, _14811_, _14809_);
  nor (_14814_, _14813_, _14812_);
  or (_14815_, _14814_, _07399_);
  and (_14816_, _14815_, _14801_);
  or (_14817_, _14816_, _07397_);
  and (_14818_, _06128_, \oc8051_golden_model_1.ACC [4]);
  nor (_14819_, _14509_, _14818_);
  nor (_14820_, _08037_, _14819_);
  and (_14821_, _08037_, _14819_);
  nor (_14822_, _14821_, _14820_);
  and (_14823_, _14822_, \oc8051_golden_model_1.PSW [7]);
  nor (_14824_, _14822_, \oc8051_golden_model_1.PSW [7]);
  nor (_14825_, _14824_, _14823_);
  nor (_14826_, _14515_, _14512_);
  not (_14827_, _14826_);
  and (_14828_, _14827_, _14825_);
  nor (_14829_, _14827_, _14825_);
  nor (_14830_, _14829_, _14828_);
  or (_14831_, _14830_, _07507_);
  and (_14832_, _14831_, _02991_);
  and (_14833_, _14832_, _14817_);
  nor (_14834_, _14416_, _08083_);
  nor (_14835_, _08081_, _14834_);
  and (_14836_, _08081_, _14834_);
  or (_14837_, _14836_, _14835_);
  not (_14838_, _14420_);
  nor (_14839_, _14838_, _14837_);
  and (_14840_, _14838_, _14837_);
  nor (_14841_, _14840_, _14839_);
  nand (_14842_, _14841_, _07541_);
  and (_14843_, _14842_, _09325_);
  or (_14844_, _14843_, _14833_);
  and (_14845_, _14844_, _14739_);
  or (_14846_, _14845_, _07721_);
  nand (_14847_, _03220_, _07721_);
  and (_14848_, _14847_, _02986_);
  and (_14849_, _14848_, _14846_);
  nor (_14850_, _11361_, _07806_);
  nor (_14851_, _14850_, _14740_);
  nor (_14852_, _14851_, _02986_);
  or (_14853_, _14852_, _05535_);
  or (_14854_, _14853_, _14849_);
  and (_14855_, _14854_, _14725_);
  or (_14856_, _14855_, _02841_);
  and (_14857_, _06170_, _04731_);
  nor (_14858_, _14857_, _14717_);
  nand (_14859_, _14858_, _02841_);
  and (_14860_, _14859_, _02839_);
  and (_14861_, _14860_, _14856_);
  nor (_14862_, _11467_, _07319_);
  nor (_14863_, _14862_, _14717_);
  nor (_14864_, _14863_, _02839_);
  or (_14865_, _14864_, _06786_);
  or (_14866_, _14865_, _14861_);
  or (_14867_, _06840_, _06792_);
  and (_14868_, _14867_, _14866_);
  and (_14869_, _14868_, _02609_);
  nor (_14870_, _03220_, _02609_);
  or (_14871_, _14870_, _02834_);
  or (_14872_, _14871_, _14869_);
  and (_14873_, _05671_, _04731_);
  nor (_14874_, _14873_, _14717_);
  nand (_14875_, _14874_, _02834_);
  and (_14876_, _14875_, _07831_);
  and (_14877_, _14876_, _14872_);
  nor (_14878_, _14877_, _14722_);
  or (_14879_, _14878_, _07843_);
  nand (_14880_, _07843_, _07198_);
  and (_14881_, _14880_, _14879_);
  nor (_14882_, _14881_, _13644_);
  and (_14883_, _13644_, _07198_);
  or (_14884_, _14883_, _13650_);
  or (_14885_, _14884_, _14882_);
  or (_14886_, _13654_, _07198_);
  and (_14887_, _14886_, _13383_);
  and (_14888_, _14887_, _14885_);
  or (_14889_, _08037_, _03521_);
  and (_14890_, _14889_, _07849_);
  or (_14891_, _14890_, _14888_);
  and (_14892_, _14891_, _14721_);
  or (_14893_, _14892_, _03146_);
  or (_14894_, _11356_, _03147_);
  and (_14895_, _14894_, _07861_);
  and (_14896_, _14895_, _14893_);
  and (_14897_, _07860_, _09265_);
  or (_14898_, _14897_, _03051_);
  or (_14899_, _14898_, _14896_);
  and (_14900_, _14899_, _14720_);
  or (_14901_, _14900_, _03148_);
  or (_14902_, _14717_, _07150_);
  and (_14903_, _14902_, _07882_);
  and (_14904_, _14903_, _14901_);
  or (_14905_, _14904_, _14716_);
  and (_14906_, _14905_, _07891_);
  and (_14907_, _07890_, _08035_);
  or (_14908_, _14907_, _03135_);
  or (_14909_, _14908_, _14906_);
  or (_14910_, _11354_, _03136_);
  and (_14911_, _14910_, _07312_);
  and (_14912_, _14911_, _14909_);
  and (_14913_, _08121_, _07311_);
  or (_14914_, _14913_, _14912_);
  and (_14915_, _14914_, _03023_);
  or (_14916_, _14874_, _11355_);
  nor (_14917_, _14916_, _03023_);
  or (_14918_, _14917_, _03751_);
  or (_14919_, _14918_, _14915_);
  nand (_14920_, _07197_, _03751_);
  nand (_14921_, _14920_, _14919_);
  nor (_14922_, _14921_, _14715_);
  not (_14923_, _07197_);
  and (_14924_, _14715_, _14923_);
  or (_14925_, _14924_, _07906_);
  or (_14926_, _14925_, _14922_);
  nand (_14927_, _07906_, _07197_);
  and (_14928_, _14927_, _07913_);
  and (_14929_, _14928_, _14926_);
  nor (_14930_, _07197_, _07913_);
  or (_14931_, _14930_, _07915_);
  or (_14932_, _14931_, _14929_);
  nand (_14933_, _07915_, _08036_);
  and (_14934_, _14933_, _03142_);
  and (_14935_, _14934_, _14932_);
  nor (_14936_, _11355_, _03142_);
  or (_14937_, _14936_, _07921_);
  or (_14938_, _14937_, _14935_);
  nand (_14939_, _07921_, _08122_);
  and (_14940_, _14939_, _03043_);
  and (_14941_, _14940_, _14938_);
  nor (_14942_, _11480_, _07319_);
  nor (_14943_, _14942_, _14717_);
  nor (_14944_, _14943_, _03043_);
  or (_14945_, _14944_, _07931_);
  or (_14946_, _14945_, _14941_);
  and (_14947_, _14946_, _14714_);
  or (_14948_, _14947_, _07229_);
  and (_14949_, _07953_, _07350_);
  nor (_14950_, _14949_, _07954_);
  or (_14951_, _14950_, _07936_);
  and (_14952_, _14951_, _03134_);
  and (_14953_, _14952_, _14948_);
  and (_14954_, _07984_, _07665_);
  nor (_14955_, _14954_, _07985_);
  and (_14956_, _14955_, _03133_);
  or (_14957_, _14956_, _07964_);
  or (_14958_, _14957_, _14953_);
  and (_14959_, _08015_, _07747_);
  nor (_14960_, _14959_, _08016_);
  or (_14961_, _14960_, _07997_);
  and (_14962_, _14961_, _07996_);
  and (_14963_, _14962_, _14958_);
  nand (_14964_, _07995_, \oc8051_golden_model_1.ACC [4]);
  nand (_14965_, _14964_, _07189_);
  or (_14966_, _14965_, _14963_);
  and (_14967_, _14966_, _14711_);
  or (_14968_, _14967_, _07185_);
  and (_14969_, _08059_, _08038_);
  nor (_14970_, _14969_, _08060_);
  or (_14971_, _14970_, _08031_);
  and (_14972_, _14971_, _03166_);
  and (_14973_, _14972_, _14968_);
  and (_14974_, _08103_, _08081_);
  nor (_14975_, _14974_, _08104_);
  and (_14976_, _14975_, _02892_);
  or (_14977_, _14976_, _08070_);
  or (_14978_, _14977_, _14973_);
  nor (_14979_, _08141_, _09265_);
  and (_14980_, _08141_, _09265_);
  or (_14981_, _14980_, _14979_);
  or (_14982_, _14981_, _08117_);
  and (_14983_, _14982_, _08116_);
  and (_14984_, _14983_, _14978_);
  and (_14985_, _08115_, \oc8051_golden_model_1.ACC [4]);
  or (_14986_, _14985_, _03174_);
  or (_14987_, _14986_, _14984_);
  nand (_14988_, _14746_, _03174_);
  and (_14989_, _14988_, _08156_);
  and (_14990_, _14989_, _14987_);
  nor (_14991_, _14681_, _06858_);
  or (_14992_, _14991_, _08163_);
  and (_14993_, _14992_, _08155_);
  or (_14994_, _14993_, _08160_);
  or (_14995_, _14994_, _14990_);
  nand (_14996_, _08160_, _06807_);
  and (_14997_, _14996_, _03183_);
  and (_14998_, _14997_, _14995_);
  nor (_14999_, _14791_, _03183_);
  or (_15000_, _14999_, _02887_);
  or (_15001_, _15000_, _14998_);
  and (_15002_, _11541_, _04731_);
  nor (_15003_, _15002_, _14717_);
  nand (_15004_, _15003_, _02887_);
  and (_15005_, _15004_, _08178_);
  and (_15006_, _15005_, _15001_);
  nor (_15007_, _08187_, \oc8051_golden_model_1.ACC [5]);
  nor (_15008_, _15007_, _08188_);
  and (_15009_, _15008_, _08177_);
  or (_15010_, _15009_, _08184_);
  or (_15011_, _15010_, _15006_);
  nand (_15012_, _08184_, _06807_);
  and (_15013_, _15012_, _34655_);
  and (_15014_, _15013_, _15011_);
  or (_15015_, _15014_, _14708_);
  and (_35827_[5], _15015_, _35796_);
  nor (_15016_, _34655_, _06807_);
  nor (_15017_, _04731_, _06807_);
  and (_15018_, _11560_, _04731_);
  nor (_15019_, _15018_, _15017_);
  nand (_15020_, _15019_, _03051_);
  nor (_15021_, _07831_, _02924_);
  nor (_15022_, _04790_, _07319_);
  nor (_15023_, _15022_, _15017_);
  nand (_15024_, _15023_, _05535_);
  nor (_15025_, _14834_, _08079_);
  or (_15026_, _15025_, _08080_);
  and (_15027_, _15026_, _08077_);
  nor (_15028_, _15026_, _08077_);
  nor (_15029_, _15028_, _15027_);
  not (_15030_, _14839_);
  nor (_15031_, _15030_, _15029_);
  and (_15032_, _15030_, _15029_);
  nor (_15033_, _15032_, _15031_);
  nand (_15034_, _15033_, _02979_);
  and (_15035_, _15034_, _07541_);
  or (_15036_, _06170_, _06858_);
  and (_15037_, _06170_, _06858_);
  or (_15038_, _14819_, _15037_);
  and (_15039_, _15038_, _15036_);
  nor (_15040_, _15039_, _08034_);
  and (_15041_, _15039_, _08034_);
  nor (_15042_, _15041_, _15040_);
  nor (_15043_, _14828_, _14823_);
  and (_15044_, _15043_, \oc8051_golden_model_1.PSW [7]);
  nor (_15045_, _15044_, _15042_);
  and (_15046_, _15044_, _15042_);
  nor (_15047_, _15046_, _15045_);
  or (_15048_, _15047_, _07507_);
  nand (_15049_, _04894_, \oc8051_golden_model_1.ACC [5]);
  nor (_15050_, _04894_, \oc8051_golden_model_1.ACC [5]);
  or (_15051_, _14803_, _15050_);
  and (_15052_, _15051_, _15049_);
  nor (_15053_, _15052_, _07195_);
  and (_15054_, _15052_, _07195_);
  nor (_15055_, _15054_, _15053_);
  nor (_15056_, _14812_, _14807_);
  and (_15057_, _15056_, \oc8051_golden_model_1.PSW [7]);
  nor (_15058_, _15057_, _15055_);
  and (_15059_, _15057_, _15055_);
  nor (_15060_, _15059_, _15058_);
  or (_15061_, _15060_, _07399_);
  nor (_15062_, _05313_, _06807_);
  and (_15063_, _11564_, _05313_);
  and (_15064_, _15063_, _11596_);
  nor (_15065_, _15064_, _15062_);
  nor (_15066_, _15065_, _06246_);
  nand (_15067_, _07403_, _04790_);
  nor (_15068_, _11567_, _07319_);
  nor (_15069_, _15068_, _15017_);
  nand (_15070_, _15069_, _02948_);
  nor (_15071_, _07552_, _03401_);
  or (_15072_, _07411_, _06162_);
  nor (_15073_, _07421_, _04790_);
  or (_15074_, _07423_, \oc8051_golden_model_1.ACC [6]);
  nand (_15075_, _07423_, \oc8051_golden_model_1.ACC [6]);
  and (_15076_, _15075_, _15074_);
  and (_15077_, _15076_, _07421_);
  or (_15078_, _15077_, _07410_);
  or (_15079_, _15078_, _15073_);
  and (_15080_, _15079_, _03401_);
  and (_15081_, _15080_, _15072_);
  or (_15082_, _15081_, _15071_);
  and (_15083_, _15082_, _07437_);
  and (_15084_, _07441_, xram_data_in_reg[6]);
  or (_15085_, _15084_, _02948_);
  or (_15086_, _15085_, _15083_);
  and (_15087_, _15086_, _15070_);
  or (_15088_, _15087_, _07405_);
  not (_15089_, _07458_);
  nor (_15090_, _14767_, _15089_);
  and (_15091_, _09861_, _07459_);
  nor (_15092_, _15091_, _15090_);
  nand (_15093_, _15092_, _07405_);
  and (_15094_, _15093_, _02976_);
  and (_15095_, _15094_, _15088_);
  nor (_15096_, _15063_, _15062_);
  nor (_15097_, _15096_, _02934_);
  nor (_15098_, _15023_, _07474_);
  or (_15099_, _15098_, _07403_);
  or (_15100_, _15099_, _15097_);
  or (_15101_, _15100_, _15095_);
  and (_15102_, _15101_, _15067_);
  or (_15103_, _15102_, _03873_);
  or (_15104_, _06162_, _07481_);
  and (_15105_, _15104_, _02992_);
  and (_15106_, _15105_, _15103_);
  nor (_15107_, _07552_, _02992_);
  or (_15108_, _15107_, _07485_);
  or (_15109_, _15108_, _15106_);
  nand (_15110_, _07485_, _06964_);
  and (_15111_, _15110_, _15109_);
  or (_15112_, _15111_, _02877_);
  and (_15113_, _11562_, _05313_);
  nor (_15114_, _15113_, _15062_);
  nand (_15115_, _15114_, _02877_);
  and (_15116_, _15115_, _06246_);
  and (_15117_, _15116_, _15112_);
  or (_15118_, _15117_, _15066_);
  and (_15119_, _15118_, _06258_);
  nor (_15120_, _06728_, _06726_);
  nor (_15121_, _15120_, _06729_);
  and (_15122_, _15121_, _06252_);
  or (_15123_, _15122_, _09326_);
  or (_15124_, _15123_, _15119_);
  and (_15125_, _15124_, _15061_);
  and (_15126_, _15125_, _15048_);
  or (_15127_, _15126_, _02979_);
  and (_15128_, _15127_, _15035_);
  nor (_15129_, _14727_, _09834_);
  nor (_15130_, _15129_, _09833_);
  nor (_15131_, _15130_, _08120_);
  and (_15132_, _15130_, _08120_);
  nor (_15133_, _15132_, _15131_);
  nor (_15134_, _14736_, _14731_);
  and (_15135_, _15134_, \oc8051_golden_model_1.PSW [7]);
  nor (_15136_, _15135_, _15133_);
  and (_15137_, _15135_, _15133_);
  nor (_15138_, _15137_, _15136_);
  and (_15139_, _15138_, _07540_);
  or (_15140_, _15139_, _07721_);
  or (_15141_, _15140_, _15128_);
  nand (_15142_, _02924_, _07721_);
  and (_15143_, _15142_, _02986_);
  and (_15144_, _15143_, _15141_);
  nor (_15145_, _11614_, _07806_);
  nor (_15146_, _15145_, _15062_);
  nor (_15147_, _15146_, _02986_);
  or (_15148_, _15147_, _05535_);
  or (_15149_, _15148_, _15144_);
  and (_15150_, _15149_, _15024_);
  or (_15151_, _15150_, _02841_);
  and (_15152_, _06162_, _04731_);
  nor (_15153_, _15152_, _15017_);
  nand (_15154_, _15153_, _02841_);
  and (_15155_, _15154_, _02839_);
  and (_15156_, _15155_, _15151_);
  nor (_15157_, _11671_, _07319_);
  nor (_15158_, _15157_, _15017_);
  nor (_15159_, _15158_, _02839_);
  or (_15160_, _15159_, _06786_);
  or (_15161_, _15160_, _15156_);
  not (_15162_, _06808_);
  and (_15163_, _06813_, _15162_);
  or (_15164_, _15163_, _06792_);
  and (_15165_, _15164_, _15161_);
  and (_15166_, _15165_, _02609_);
  nor (_15167_, _02924_, _02609_);
  or (_15168_, _15167_, _02834_);
  or (_15169_, _15168_, _15166_);
  and (_15170_, _11678_, _04731_);
  nor (_15171_, _15170_, _15017_);
  nand (_15172_, _15171_, _02834_);
  and (_15173_, _15172_, _07831_);
  and (_15174_, _15173_, _15169_);
  or (_15175_, _15174_, _15021_);
  and (_15176_, _15175_, _07845_);
  and (_15177_, _07846_, _07195_);
  or (_15178_, _15177_, _15176_);
  and (_15179_, _15178_, _13383_);
  and (_15180_, _13382_, _08034_);
  or (_15181_, _15180_, _15179_);
  and (_15182_, _15181_, _13261_);
  and (_15183_, _08034_, _03521_);
  or (_15184_, _15183_, _03146_);
  or (_15185_, _15184_, _15182_);
  or (_15186_, _11556_, _03147_);
  and (_15187_, _15186_, _07861_);
  and (_15188_, _15187_, _15185_);
  and (_15189_, _07860_, _08120_);
  or (_15190_, _15189_, _03051_);
  or (_15191_, _15190_, _15188_);
  and (_15192_, _15191_, _15020_);
  or (_15193_, _15192_, _03148_);
  or (_15194_, _15017_, _07150_);
  and (_15195_, _15194_, _07882_);
  and (_15196_, _15195_, _15193_);
  and (_15197_, _07883_, _07193_);
  or (_15198_, _15197_, _07890_);
  or (_15199_, _15198_, _15196_);
  or (_15200_, _07891_, _08032_);
  and (_15201_, _15200_, _03136_);
  and (_15202_, _15201_, _15199_);
  and (_15203_, _11554_, _03135_);
  or (_15204_, _15203_, _07311_);
  or (_15205_, _15204_, _15202_);
  or (_15206_, _08118_, _07312_);
  and (_15207_, _15206_, _03023_);
  and (_15208_, _15207_, _15205_);
  or (_15209_, _15171_, _11555_);
  nor (_15210_, _15209_, _03023_);
  or (_15211_, _15210_, _13415_);
  or (_15212_, _15211_, _15208_);
  or (_15213_, _07194_, _03757_);
  nand (_15214_, _15213_, _13416_);
  and (_15215_, _15214_, _13422_);
  and (_15216_, _15215_, _15212_);
  nor (_15217_, _13421_, _03757_);
  nor (_15218_, _15217_, _07194_);
  or (_15219_, _15218_, _07915_);
  or (_15220_, _15219_, _15216_);
  nand (_15221_, _07915_, _08033_);
  and (_15222_, _15221_, _03142_);
  and (_15223_, _15222_, _15220_);
  nor (_15224_, _11555_, _03142_);
  or (_15225_, _15224_, _07921_);
  or (_15226_, _15225_, _15223_);
  nand (_15227_, _07921_, _08119_);
  nand (_15228_, _15227_, _15226_);
  and (_15229_, _15228_, _03043_);
  nor (_15230_, _11558_, _07319_);
  nor (_15231_, _15230_, _15017_);
  and (_15232_, _15231_, _03042_);
  or (_15233_, _15232_, _07931_);
  nor (_15234_, _15233_, _15229_);
  and (_15235_, _07302_, _07250_);
  nor (_15236_, _15235_, _07303_);
  or (_15237_, _15236_, _07229_);
  and (_15238_, _15237_, _09487_);
  or (_15239_, _15238_, _15234_);
  and (_15240_, _07955_, _07938_);
  nor (_15241_, _15240_, _07956_);
  or (_15242_, _15241_, _07936_);
  and (_15243_, _15242_, _03134_);
  and (_15244_, _15243_, _15239_);
  and (_15245_, _07986_, _07968_);
  nor (_15246_, _15245_, _07987_);
  and (_15247_, _15246_, _03133_);
  or (_15248_, _15247_, _07964_);
  or (_15250_, _15248_, _15244_);
  and (_15251_, _08017_, _07999_);
  nor (_15252_, _15251_, _08018_);
  or (_15253_, _15252_, _07997_);
  and (_15254_, _15253_, _15250_);
  or (_15255_, _15254_, _07995_);
  nand (_15256_, _07995_, _06858_);
  and (_15257_, _15256_, _07189_);
  and (_15258_, _15257_, _15255_);
  nor (_15259_, _07222_, _07195_);
  nor (_15261_, _15259_, _07223_);
  and (_15262_, _15261_, _10153_);
  or (_15263_, _15262_, _15258_);
  and (_15264_, _15263_, _08031_);
  nor (_15265_, _08061_, _08034_);
  nor (_15266_, _15265_, _08062_);
  and (_15267_, _15266_, _07185_);
  or (_15268_, _15267_, _08112_);
  or (_15269_, _15268_, _15264_);
  and (_15270_, _08105_, _08077_);
  nor (_15272_, _15270_, _08106_);
  or (_15273_, _15272_, _10168_);
  nor (_15274_, _08143_, _08120_);
  nor (_15275_, _15274_, _08144_);
  or (_15276_, _15275_, _08117_);
  and (_15277_, _15276_, _08116_);
  and (_15278_, _15277_, _15273_);
  and (_15279_, _15278_, _15269_);
  and (_15280_, _08115_, \oc8051_golden_model_1.ACC [5]);
  or (_15281_, _15280_, _03174_);
  or (_15283_, _15281_, _15279_);
  nand (_15284_, _15069_, _03174_);
  and (_15285_, _15284_, _08156_);
  and (_15286_, _15285_, _15283_);
  nor (_15287_, _08163_, _06807_);
  or (_15288_, _15287_, _08164_);
  nor (_15289_, _15288_, _08160_);
  nor (_15290_, _15289_, _09732_);
  or (_15291_, _15290_, _15286_);
  nand (_15292_, _08160_, _05364_);
  and (_15294_, _15292_, _03183_);
  and (_15295_, _15294_, _15291_);
  nor (_15296_, _15114_, _03183_);
  or (_15297_, _15296_, _02887_);
  or (_15298_, _15297_, _15295_);
  and (_15299_, _11744_, _04731_);
  nor (_15300_, _15299_, _15017_);
  nand (_15301_, _15300_, _02887_);
  and (_15302_, _15301_, _08178_);
  and (_15303_, _15302_, _15298_);
  nor (_15305_, _08188_, \oc8051_golden_model_1.ACC [6]);
  nor (_15306_, _15305_, _08189_);
  and (_15307_, _15306_, _08177_);
  or (_15308_, _15307_, _08184_);
  or (_15309_, _15308_, _15303_);
  nand (_15310_, _08184_, _05364_);
  and (_15311_, _15310_, _34655_);
  and (_15312_, _15311_, _15309_);
  or (_15313_, _15312_, _15016_);
  and (_35827_[6], _15313_, _35796_);
  not (_15315_, \oc8051_golden_model_1.DPL [0]);
  nor (_15316_, _34655_, _15315_);
  nor (_15317_, _05085_, _08203_);
  nor (_15318_, _04643_, _15315_);
  and (_15319_, _04643_, _05660_);
  or (_15320_, _15319_, _15318_);
  nand (_15321_, _15320_, _03022_);
  nor (_15322_, _15321_, _15317_);
  and (_15323_, _04643_, \oc8051_golden_model_1.ACC [0]);
  or (_15324_, _15323_, _15318_);
  or (_15326_, _15324_, _02992_);
  or (_15327_, _15318_, _15317_);
  or (_15328_, _15327_, _03006_);
  and (_15329_, _15324_, _03845_);
  nor (_15330_, _03845_, _15315_);
  or (_15331_, _15330_, _02948_);
  or (_15332_, _15331_, _15329_);
  and (_15333_, _15332_, _07474_);
  and (_15334_, _15333_, _15328_);
  and (_15335_, _04643_, _03838_);
  or (_15337_, _15335_, _15318_);
  and (_15338_, _15337_, _02946_);
  or (_15339_, _15338_, _02880_);
  or (_15340_, _15339_, _15334_);
  and (_15341_, _15340_, _15326_);
  or (_15342_, _15341_, _08226_);
  and (_15343_, _08226_, \oc8051_golden_model_1.DPL [0]);
  nor (_15344_, _15343_, _03046_);
  and (_15345_, _15344_, _15342_);
  nor (_15346_, _03505_, _08211_);
  or (_15348_, _15346_, _05535_);
  or (_15349_, _15348_, _15345_);
  or (_15350_, _15337_, _02859_);
  and (_15351_, _15350_, _15349_);
  or (_15352_, _15351_, _02841_);
  and (_15353_, _06164_, _04643_);
  or (_15354_, _15318_, _02842_);
  or (_15355_, _15354_, _15353_);
  and (_15356_, _15355_, _15352_);
  and (_15357_, _15356_, _02839_);
  nor (_15359_, _10475_, _08203_);
  or (_15360_, _15359_, _15318_);
  and (_15361_, _15360_, _02567_);
  or (_15362_, _15361_, _02834_);
  or (_15363_, _15362_, _15357_);
  or (_15364_, _15320_, _07140_);
  and (_15365_, _15364_, _07139_);
  and (_15366_, _15365_, _15363_);
  and (_15367_, _10372_, _04643_);
  or (_15368_, _15318_, _03148_);
  nor (_15370_, _15368_, _15367_);
  nor (_15371_, _15370_, _03149_);
  or (_15372_, _15371_, _15366_);
  and (_15373_, _10369_, _04643_);
  or (_15374_, _15318_, _07150_);
  or (_15375_, _15374_, _15373_);
  and (_15376_, _15375_, _03023_);
  and (_15377_, _15376_, _15372_);
  or (_15378_, _15377_, _15322_);
  and (_15379_, _15378_, _06213_);
  or (_15381_, _15318_, _05085_);
  and (_15382_, _15324_, _03137_);
  and (_15383_, _15382_, _15381_);
  or (_15384_, _15383_, _03042_);
  or (_15385_, _15384_, _15379_);
  nor (_15386_, _10365_, _08203_);
  or (_15387_, _15318_, _03043_);
  or (_15388_, _15387_, _15386_);
  and (_15389_, _15388_, _07161_);
  and (_15390_, _15389_, _15385_);
  nor (_15392_, _10367_, _08203_);
  or (_15393_, _15392_, _15318_);
  and (_15394_, _15393_, _03143_);
  or (_15395_, _15394_, _03361_);
  or (_15396_, _15395_, _15390_);
  or (_15397_, _15327_, _03360_);
  and (_15398_, _15397_, _34655_);
  and (_15399_, _15398_, _15396_);
  or (_15400_, _15399_, _15316_);
  and (_35830_[0], _15400_, _35796_);
  not (_15402_, \oc8051_golden_model_1.DPL [1]);
  nor (_15403_, _34655_, _15402_);
  nor (_15404_, _04643_, _15402_);
  nor (_15405_, _08203_, _04020_);
  or (_15406_, _15405_, _15404_);
  or (_15407_, _15406_, _07474_);
  or (_15408_, _04643_, \oc8051_golden_model_1.DPL [1]);
  and (_15409_, _10574_, _04643_);
  not (_15410_, _15409_);
  and (_15411_, _15410_, _15408_);
  and (_15413_, _15411_, _02948_);
  nand (_15414_, _04643_, _02543_);
  and (_15415_, _15414_, _15408_);
  and (_15416_, _15415_, _03845_);
  nor (_15417_, _03845_, _15402_);
  or (_15418_, _15417_, _15416_);
  and (_15419_, _15418_, _03006_);
  or (_15420_, _15419_, _02946_);
  or (_15421_, _15420_, _15413_);
  and (_15422_, _15421_, _15407_);
  or (_15423_, _15422_, _02880_);
  or (_15424_, _15415_, _02992_);
  and (_15425_, _15424_, _08227_);
  and (_15426_, _15425_, _15423_);
  nor (_15427_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_15428_, _15427_, _08231_);
  and (_15429_, _15428_, _08226_);
  or (_15430_, _15429_, _15426_);
  and (_15431_, _15430_, _08211_);
  nor (_15432_, _03720_, _08211_);
  or (_15434_, _15432_, _05535_);
  or (_15435_, _15434_, _15431_);
  or (_15436_, _15406_, _02859_);
  and (_15437_, _15436_, _15435_);
  or (_15438_, _15437_, _02841_);
  and (_15439_, _06163_, _04643_);
  or (_15440_, _15404_, _02842_);
  or (_15441_, _15440_, _15439_);
  and (_15442_, _15441_, _02839_);
  and (_15443_, _15442_, _15438_);
  and (_15445_, _10674_, _04643_);
  or (_15446_, _15445_, _15404_);
  and (_15447_, _15446_, _02567_);
  or (_15448_, _15447_, _15443_);
  and (_15449_, _15448_, _03052_);
  or (_15450_, _10689_, _08203_);
  and (_15451_, _15408_, _03051_);
  and (_15452_, _15451_, _15450_);
  nand (_15453_, _04643_, _03720_);
  and (_15454_, _15408_, _02834_);
  and (_15456_, _15454_, _15453_);
  or (_15457_, _15456_, _15452_);
  or (_15458_, _15457_, _15449_);
  and (_15459_, _15458_, _07150_);
  or (_15460_, _10565_, _08203_);
  and (_15461_, _15408_, _03148_);
  and (_15462_, _15461_, _15460_);
  or (_15463_, _15462_, _15459_);
  and (_15464_, _15463_, _03138_);
  or (_15465_, _15404_, _05038_);
  and (_15467_, _15415_, _03137_);
  and (_15468_, _15467_, _15465_);
  or (_15469_, _10688_, _08203_);
  and (_15470_, _15408_, _03022_);
  and (_15471_, _15470_, _15469_);
  or (_15472_, _15471_, _15468_);
  or (_15473_, _15472_, _15464_);
  and (_15474_, _15473_, _03144_);
  or (_15475_, _15414_, _05038_);
  and (_15476_, _15408_, _03143_);
  and (_15478_, _15476_, _15475_);
  or (_15479_, _15478_, _03174_);
  or (_15480_, _15453_, _05038_);
  and (_15481_, _15408_, _03042_);
  and (_15482_, _15481_, _15480_);
  or (_15483_, _15482_, _15479_);
  or (_15484_, _15483_, _15474_);
  or (_15485_, _15411_, _03179_);
  and (_15486_, _15485_, _15484_);
  or (_15487_, _15486_, _02887_);
  or (_15489_, _15404_, _02888_);
  or (_15490_, _15489_, _15409_);
  and (_15491_, _15490_, _34655_);
  and (_15492_, _15491_, _15487_);
  or (_15493_, _15492_, _15403_);
  and (_35830_[1], _15493_, _35796_);
  not (_15494_, \oc8051_golden_model_1.DPL [2]);
  nor (_15495_, _34655_, _15494_);
  nor (_15496_, _04643_, _15494_);
  nor (_15497_, _10765_, _08203_);
  or (_15499_, _15497_, _15496_);
  and (_15500_, _15499_, _03143_);
  and (_15501_, _10766_, _04643_);
  or (_15502_, _15501_, _15496_);
  and (_15503_, _15502_, _03148_);
  nor (_15504_, _08203_, _04449_);
  or (_15505_, _15504_, _15496_);
  or (_15506_, _15505_, _07474_);
  nor (_15507_, _10788_, _08203_);
  or (_15508_, _15507_, _15496_);
  and (_15510_, _15508_, _02948_);
  nor (_15511_, _03845_, _15494_);
  and (_15512_, _04643_, \oc8051_golden_model_1.ACC [2]);
  or (_15513_, _15512_, _15496_);
  and (_15514_, _15513_, _03845_);
  or (_15515_, _15514_, _15511_);
  and (_15516_, _15515_, _03006_);
  or (_15517_, _15516_, _02946_);
  or (_15518_, _15517_, _15510_);
  and (_15519_, _15518_, _15506_);
  or (_15521_, _15519_, _02880_);
  or (_15522_, _15513_, _02992_);
  and (_15523_, _15522_, _08227_);
  and (_15524_, _15523_, _15521_);
  nor (_15525_, _08231_, \oc8051_golden_model_1.DPL [2]);
  nor (_15526_, _15525_, _08232_);
  and (_15527_, _15526_, _08226_);
  or (_15528_, _15527_, _15524_);
  and (_15529_, _15528_, _08211_);
  nor (_15530_, _03262_, _08211_);
  or (_15532_, _15530_, _05535_);
  or (_15533_, _15532_, _15529_);
  or (_15534_, _15505_, _02859_);
  and (_15535_, _15534_, _15533_);
  or (_15536_, _15535_, _02841_);
  and (_15537_, _06167_, _04643_);
  or (_15538_, _15496_, _02842_);
  or (_15539_, _15538_, _15537_);
  and (_15540_, _15539_, _02839_);
  and (_15541_, _15540_, _15536_);
  nor (_15543_, _10881_, _08203_);
  or (_15544_, _15543_, _15496_);
  and (_15545_, _15544_, _02567_);
  or (_15546_, _15545_, _08207_);
  or (_15547_, _15546_, _15541_);
  and (_15548_, _10770_, _04643_);
  or (_15549_, _15496_, _07139_);
  or (_15550_, _15549_, _15548_);
  and (_15551_, _04643_, _05693_);
  or (_15552_, _15551_, _15496_);
  or (_15554_, _15552_, _07140_);
  and (_15555_, _15554_, _07150_);
  and (_15556_, _15555_, _15550_);
  and (_15557_, _15556_, _15547_);
  or (_15558_, _15557_, _15503_);
  and (_15559_, _15558_, _03138_);
  or (_15560_, _15496_, _05135_);
  and (_15561_, _15513_, _03137_);
  and (_15562_, _15552_, _03022_);
  or (_15563_, _15562_, _15561_);
  and (_15565_, _15563_, _15560_);
  or (_15566_, _15565_, _03042_);
  or (_15567_, _15566_, _15559_);
  nor (_15568_, _10768_, _08203_);
  or (_15569_, _15496_, _03043_);
  or (_15570_, _15569_, _15568_);
  and (_15571_, _15570_, _07161_);
  and (_15572_, _15571_, _15567_);
  or (_15573_, _15572_, _15500_);
  and (_15574_, _15573_, _03179_);
  and (_15576_, _15508_, _03174_);
  or (_15577_, _15576_, _02887_);
  or (_15578_, _15577_, _15574_);
  and (_15579_, _10941_, _04643_);
  or (_15580_, _15496_, _02888_);
  or (_15581_, _15580_, _15579_);
  and (_15582_, _15581_, _34655_);
  and (_15583_, _15582_, _15578_);
  or (_15584_, _15583_, _15495_);
  and (_35830_[2], _15584_, _35796_);
  or (_15586_, _34655_, \oc8051_golden_model_1.DPL [3]);
  and (_15587_, _15586_, _35796_);
  not (_15588_, \oc8051_golden_model_1.DPL [3]);
  nor (_15589_, _04643_, _15588_);
  and (_15590_, _10964_, _04643_);
  or (_15591_, _15590_, _15589_);
  and (_15592_, _15591_, _03148_);
  nor (_15593_, _10983_, _08203_);
  or (_15594_, _15593_, _15589_);
  or (_15595_, _15594_, _03006_);
  and (_15597_, _04643_, \oc8051_golden_model_1.ACC [3]);
  or (_15598_, _15597_, _15589_);
  and (_15599_, _15598_, _03845_);
  nor (_15600_, _03845_, _15588_);
  or (_15601_, _15600_, _02948_);
  or (_15602_, _15601_, _15599_);
  and (_15603_, _15602_, _07474_);
  and (_15604_, _15603_, _15595_);
  nor (_15605_, _08203_, _04275_);
  or (_15606_, _15605_, _15589_);
  and (_15608_, _15606_, _02946_);
  or (_15609_, _15608_, _02880_);
  or (_15610_, _15609_, _15604_);
  or (_15611_, _15598_, _02992_);
  and (_15612_, _15611_, _08227_);
  and (_15613_, _15612_, _15610_);
  nor (_15614_, _08232_, \oc8051_golden_model_1.DPL [3]);
  nor (_15615_, _15614_, _08233_);
  and (_15616_, _15615_, _08226_);
  or (_15617_, _15616_, _15613_);
  and (_15619_, _15617_, _08211_);
  nor (_15620_, _03128_, _08211_);
  or (_15621_, _15620_, _05535_);
  or (_15622_, _15621_, _15619_);
  or (_15623_, _15606_, _02859_);
  and (_15624_, _15623_, _15622_);
  or (_15625_, _15624_, _02841_);
  and (_15626_, _06166_, _04643_);
  or (_15627_, _15589_, _02842_);
  or (_15628_, _15627_, _15626_);
  and (_15630_, _15628_, _02839_);
  and (_15631_, _15630_, _15625_);
  nor (_15632_, _11076_, _08203_);
  or (_15633_, _15632_, _15589_);
  and (_15634_, _15633_, _02567_);
  or (_15635_, _15634_, _08207_);
  or (_15636_, _15635_, _15631_);
  and (_15637_, _10968_, _04643_);
  or (_15638_, _15589_, _07139_);
  or (_15639_, _15638_, _15637_);
  and (_15641_, _04643_, _05654_);
  or (_15642_, _15641_, _15589_);
  or (_15643_, _15642_, _07140_);
  and (_15644_, _15643_, _07150_);
  and (_15645_, _15644_, _15639_);
  and (_15646_, _15645_, _15636_);
  or (_15647_, _15646_, _15592_);
  and (_15648_, _15647_, _03138_);
  or (_15649_, _15589_, _04993_);
  and (_15650_, _15598_, _03137_);
  and (_15652_, _15642_, _03022_);
  or (_15653_, _15652_, _15650_);
  and (_15654_, _15653_, _15649_);
  or (_15655_, _15654_, _03042_);
  or (_15656_, _15655_, _15648_);
  nor (_15657_, _10967_, _08203_);
  or (_15658_, _15589_, _03043_);
  or (_15659_, _15658_, _15657_);
  and (_15660_, _15659_, _07161_);
  and (_15661_, _15660_, _15656_);
  nor (_15663_, _10962_, _08203_);
  or (_15664_, _15663_, _15589_);
  and (_15665_, _15664_, _03143_);
  or (_15666_, _15665_, _03174_);
  or (_15667_, _15666_, _15661_);
  or (_15668_, _15594_, _03179_);
  and (_15669_, _15668_, _02888_);
  and (_15670_, _15669_, _15667_);
  and (_15671_, _11136_, _04643_);
  or (_15672_, _15671_, _15589_);
  and (_15674_, _15672_, _02887_);
  or (_15675_, _15674_, _34659_);
  or (_15676_, _15675_, _15670_);
  and (_35830_[3], _15676_, _15587_);
  or (_15677_, _34655_, \oc8051_golden_model_1.DPL [4]);
  and (_15678_, _15677_, _35796_);
  not (_15679_, \oc8051_golden_model_1.DPL [4]);
  nor (_15680_, _04643_, _15679_);
  nor (_15681_, _05192_, _08203_);
  or (_15682_, _15681_, _15680_);
  or (_15684_, _15682_, _02859_);
  nor (_15685_, _11184_, _08203_);
  or (_15686_, _15685_, _15680_);
  or (_15687_, _15686_, _03006_);
  and (_15688_, _04643_, \oc8051_golden_model_1.ACC [4]);
  or (_15689_, _15688_, _15680_);
  and (_15690_, _15689_, _03845_);
  nor (_15691_, _03845_, _15679_);
  or (_15692_, _15691_, _02948_);
  or (_15693_, _15692_, _15690_);
  and (_15695_, _15693_, _07474_);
  and (_15696_, _15695_, _15687_);
  and (_15697_, _15682_, _02946_);
  or (_15698_, _15697_, _02880_);
  or (_15699_, _15698_, _15696_);
  or (_15700_, _15689_, _02992_);
  and (_15701_, _15700_, _08227_);
  and (_15702_, _15701_, _15699_);
  nor (_15703_, _08233_, \oc8051_golden_model_1.DPL [4]);
  nor (_15704_, _15703_, _08234_);
  and (_15706_, _15704_, _08226_);
  or (_15707_, _15706_, _15702_);
  and (_15708_, _15707_, _08211_);
  nor (_15709_, _05617_, _08211_);
  or (_15710_, _15709_, _05535_);
  or (_15711_, _15710_, _15708_);
  and (_15712_, _15711_, _15684_);
  or (_15713_, _15712_, _02841_);
  and (_15714_, _06171_, _04643_);
  or (_15715_, _15680_, _02842_);
  or (_15717_, _15715_, _15714_);
  and (_15718_, _15717_, _02839_);
  and (_15719_, _15718_, _15713_);
  nor (_15720_, _11271_, _08203_);
  or (_15721_, _15720_, _15680_);
  and (_15722_, _15721_, _02567_);
  or (_15723_, _15722_, _15719_);
  or (_15724_, _15723_, _08207_);
  and (_15725_, _11158_, _04643_);
  or (_15726_, _15680_, _07139_);
  or (_15728_, _15726_, _15725_);
  and (_15729_, _05618_, _04643_);
  or (_15730_, _15729_, _15680_);
  or (_15731_, _15730_, _07140_);
  and (_15732_, _15731_, _07150_);
  and (_15733_, _15732_, _15728_);
  and (_15734_, _15733_, _15724_);
  and (_15735_, _11154_, _04643_);
  or (_15736_, _15735_, _15680_);
  and (_15737_, _15736_, _03148_);
  or (_15739_, _15737_, _15734_);
  and (_15740_, _15739_, _03138_);
  or (_15741_, _15680_, _05240_);
  and (_15742_, _15689_, _03137_);
  and (_15743_, _15730_, _03022_);
  or (_15744_, _15743_, _15742_);
  and (_15745_, _15744_, _15741_);
  or (_15746_, _15745_, _03042_);
  or (_15747_, _15746_, _15740_);
  nor (_15748_, _11157_, _08203_);
  or (_15750_, _15680_, _03043_);
  or (_15751_, _15750_, _15748_);
  and (_15752_, _15751_, _07161_);
  and (_15753_, _15752_, _15747_);
  nor (_15754_, _11152_, _08203_);
  or (_15755_, _15754_, _15680_);
  and (_15756_, _15755_, _03143_);
  or (_15757_, _15756_, _03174_);
  or (_15758_, _15757_, _15753_);
  or (_15759_, _15686_, _03179_);
  and (_15761_, _15759_, _02888_);
  and (_15762_, _15761_, _15758_);
  and (_15763_, _11338_, _04643_);
  or (_15764_, _15763_, _15680_);
  and (_15765_, _15764_, _02887_);
  or (_15766_, _15765_, _34659_);
  or (_15767_, _15766_, _15762_);
  and (_35830_[4], _15767_, _15678_);
  or (_15768_, _34655_, \oc8051_golden_model_1.DPL [5]);
  and (_15769_, _15768_, _35796_);
  not (_15771_, \oc8051_golden_model_1.DPL [5]);
  nor (_15772_, _04643_, _15771_);
  nor (_15773_, _04894_, _08203_);
  or (_15774_, _15773_, _15772_);
  or (_15775_, _15774_, _02859_);
  nor (_15776_, _11380_, _08203_);
  or (_15777_, _15776_, _15772_);
  or (_15778_, _15777_, _03006_);
  and (_15779_, _04643_, \oc8051_golden_model_1.ACC [5]);
  or (_15780_, _15779_, _15772_);
  and (_15782_, _15780_, _03845_);
  nor (_15783_, _03845_, _15771_);
  or (_15784_, _15783_, _02948_);
  or (_15785_, _15784_, _15782_);
  and (_15786_, _15785_, _07474_);
  and (_15787_, _15786_, _15778_);
  and (_15788_, _15774_, _02946_);
  or (_15789_, _15788_, _02880_);
  or (_15790_, _15789_, _15787_);
  or (_15791_, _15780_, _02992_);
  and (_15793_, _15791_, _08227_);
  and (_15794_, _15793_, _15790_);
  nor (_15795_, _08234_, \oc8051_golden_model_1.DPL [5]);
  nor (_15796_, _15795_, _08235_);
  and (_15797_, _15796_, _08226_);
  or (_15798_, _15797_, _15794_);
  and (_15799_, _15798_, _08211_);
  nor (_15800_, _05649_, _08211_);
  or (_15801_, _15800_, _05535_);
  or (_15802_, _15801_, _15799_);
  and (_15804_, _15802_, _15775_);
  or (_15805_, _15804_, _02841_);
  and (_15806_, _06170_, _04643_);
  or (_15807_, _15772_, _02842_);
  or (_15808_, _15807_, _15806_);
  and (_15809_, _15808_, _02839_);
  and (_15810_, _15809_, _15805_);
  nor (_15811_, _11467_, _08203_);
  or (_15812_, _15811_, _15772_);
  and (_15813_, _15812_, _02567_);
  or (_15815_, _15813_, _15810_);
  or (_15816_, _15815_, _08207_);
  and (_15817_, _11482_, _04643_);
  or (_15818_, _15772_, _07139_);
  or (_15819_, _15818_, _15817_);
  and (_15820_, _05671_, _04643_);
  or (_15821_, _15820_, _15772_);
  or (_15822_, _15821_, _07140_);
  and (_15823_, _15822_, _07150_);
  and (_15824_, _15823_, _15819_);
  and (_15826_, _15824_, _15816_);
  and (_15827_, _11356_, _04643_);
  or (_15828_, _15827_, _15772_);
  and (_15829_, _15828_, _03148_);
  or (_15830_, _15829_, _15826_);
  and (_15831_, _15830_, _03138_);
  or (_15832_, _15772_, _04945_);
  and (_15833_, _15780_, _03137_);
  and (_15834_, _15821_, _03022_);
  or (_15835_, _15834_, _15833_);
  and (_15837_, _15835_, _15832_);
  or (_15838_, _15837_, _03042_);
  or (_15839_, _15838_, _15831_);
  nor (_15840_, _11480_, _08203_);
  or (_15841_, _15772_, _03043_);
  or (_15842_, _15841_, _15840_);
  and (_15843_, _15842_, _07161_);
  and (_15844_, _15843_, _15839_);
  nor (_15845_, _11355_, _08203_);
  or (_15846_, _15845_, _15772_);
  and (_15848_, _15846_, _03143_);
  or (_15849_, _15848_, _03174_);
  or (_15850_, _15849_, _15844_);
  or (_15851_, _15777_, _03179_);
  and (_15852_, _15851_, _02888_);
  and (_15853_, _15852_, _15850_);
  and (_15854_, _11541_, _04643_);
  or (_15855_, _15854_, _15772_);
  and (_15856_, _15855_, _02887_);
  or (_15857_, _15856_, _34659_);
  or (_15859_, _15857_, _15853_);
  and (_35830_[5], _15859_, _15769_);
  or (_15860_, _34655_, \oc8051_golden_model_1.DPL [6]);
  and (_15861_, _15860_, _35796_);
  not (_15862_, \oc8051_golden_model_1.DPL [6]);
  nor (_15863_, _04643_, _15862_);
  nor (_15864_, _04790_, _08203_);
  or (_15865_, _15864_, _15863_);
  or (_15866_, _15865_, _02859_);
  nor (_15867_, _11567_, _08203_);
  or (_15869_, _15867_, _15863_);
  or (_15870_, _15869_, _03006_);
  and (_15871_, _04643_, \oc8051_golden_model_1.ACC [6]);
  or (_15872_, _15871_, _15863_);
  and (_15873_, _15872_, _03845_);
  nor (_15874_, _03845_, _15862_);
  or (_15875_, _15874_, _02948_);
  or (_15876_, _15875_, _15873_);
  and (_15877_, _15876_, _07474_);
  and (_15878_, _15877_, _15870_);
  and (_15880_, _15865_, _02946_);
  or (_15881_, _15880_, _02880_);
  or (_15882_, _15881_, _15878_);
  or (_15883_, _15872_, _02992_);
  and (_15884_, _15883_, _08227_);
  and (_15885_, _15884_, _15882_);
  nor (_15886_, _08235_, \oc8051_golden_model_1.DPL [6]);
  nor (_15887_, _15886_, _08236_);
  and (_15888_, _15887_, _08226_);
  or (_15889_, _15888_, _15885_);
  and (_15891_, _15889_, _08211_);
  nor (_15892_, _05585_, _08211_);
  or (_15893_, _15892_, _05535_);
  or (_15894_, _15893_, _15891_);
  and (_15895_, _15894_, _15866_);
  or (_15896_, _15895_, _02841_);
  and (_15897_, _06162_, _04643_);
  or (_15898_, _15863_, _02842_);
  or (_15899_, _15898_, _15897_);
  and (_15900_, _15899_, _02839_);
  and (_15902_, _15900_, _15896_);
  nor (_15903_, _11671_, _08203_);
  or (_15904_, _15903_, _15863_);
  and (_15905_, _15904_, _02567_);
  or (_15906_, _15905_, _15902_);
  or (_15907_, _15906_, _08207_);
  and (_15908_, _11560_, _04643_);
  or (_15909_, _15863_, _07139_);
  or (_15910_, _15909_, _15908_);
  and (_15911_, _11678_, _04643_);
  or (_15913_, _15911_, _15863_);
  or (_15914_, _15913_, _07140_);
  and (_15915_, _15914_, _07150_);
  and (_15916_, _15915_, _15910_);
  and (_15917_, _15916_, _15907_);
  and (_15918_, _11556_, _04643_);
  or (_15919_, _15918_, _15863_);
  and (_15920_, _15919_, _03148_);
  or (_15921_, _15920_, _15917_);
  and (_15922_, _15921_, _03138_);
  or (_15924_, _15863_, _04838_);
  and (_15925_, _15872_, _03137_);
  and (_15926_, _15913_, _03022_);
  or (_15927_, _15926_, _15925_);
  and (_15928_, _15927_, _15924_);
  or (_15929_, _15928_, _03042_);
  or (_15930_, _15929_, _15922_);
  nor (_15931_, _11558_, _08203_);
  or (_15932_, _15863_, _03043_);
  or (_15933_, _15932_, _15931_);
  and (_15935_, _15933_, _07161_);
  and (_15936_, _15935_, _15930_);
  nor (_15937_, _11555_, _08203_);
  or (_15938_, _15937_, _15863_);
  and (_15939_, _15938_, _03143_);
  or (_15940_, _15939_, _03174_);
  or (_15941_, _15940_, _15936_);
  or (_15942_, _15869_, _03179_);
  and (_15943_, _15942_, _02888_);
  and (_15944_, _15943_, _15941_);
  and (_15946_, _11744_, _04643_);
  or (_15947_, _15946_, _15863_);
  and (_15948_, _15947_, _02887_);
  or (_15949_, _15948_, _34659_);
  or (_15950_, _15949_, _15944_);
  and (_35830_[6], _15950_, _15861_);
  nor (_15951_, _34655_, _09380_);
  nor (_15952_, _08298_, _09380_);
  and (_15953_, _04696_, _03838_);
  or (_15954_, _15953_, _15952_);
  or (_15956_, _15954_, _02859_);
  nor (_15957_, _08238_, \oc8051_golden_model_1.DPH [0]);
  nor (_15958_, _15957_, _08324_);
  and (_15959_, _15958_, _08226_);
  nor (_15960_, _05085_, _08300_);
  or (_15961_, _15960_, _15952_);
  or (_15962_, _15961_, _03006_);
  and (_15963_, _08298_, \oc8051_golden_model_1.ACC [0]);
  or (_15964_, _15963_, _15952_);
  and (_15965_, _15964_, _03845_);
  nor (_15967_, _03845_, _09380_);
  or (_15968_, _15967_, _02948_);
  or (_15969_, _15968_, _15965_);
  and (_15970_, _15969_, _07474_);
  and (_15971_, _15970_, _15962_);
  and (_15972_, _15954_, _02946_);
  or (_15973_, _15972_, _02880_);
  or (_15974_, _15973_, _15971_);
  or (_15975_, _15964_, _02992_);
  and (_15976_, _15975_, _08227_);
  and (_15978_, _15976_, _15974_);
  or (_15979_, _15978_, _15959_);
  and (_15980_, _15979_, _08211_);
  and (_15981_, _03046_, _02833_);
  or (_15982_, _15981_, _05535_);
  or (_15983_, _15982_, _15980_);
  and (_15984_, _15983_, _15956_);
  or (_15985_, _15984_, _02841_);
  or (_15986_, _15952_, _02842_);
  and (_15987_, _06164_, _08298_);
  or (_15989_, _15987_, _15986_);
  and (_15990_, _15989_, _15985_);
  and (_15991_, _15990_, _02839_);
  nor (_15992_, _10475_, _08300_);
  or (_15993_, _15992_, _15952_);
  and (_15994_, _15993_, _02567_);
  or (_15995_, _15994_, _02834_);
  or (_15996_, _15995_, _15991_);
  and (_15997_, _08298_, _05660_);
  or (_15998_, _15997_, _15952_);
  or (_16000_, _15998_, _07140_);
  and (_16001_, _16000_, _07139_);
  and (_16002_, _16001_, _15996_);
  nand (_16003_, _10372_, _04696_);
  nor (_16004_, _15952_, _03148_);
  and (_16005_, _16004_, _16003_);
  nor (_16006_, _16005_, _03149_);
  or (_16007_, _16006_, _16002_);
  and (_16008_, _10369_, _04696_);
  or (_16009_, _15952_, _07150_);
  or (_16011_, _16009_, _16008_);
  and (_16012_, _16011_, _03023_);
  and (_16013_, _16012_, _16007_);
  nand (_16014_, _15998_, _03022_);
  nor (_16015_, _16014_, _15960_);
  or (_16016_, _16015_, _16013_);
  and (_16017_, _16016_, _06213_);
  or (_16018_, _15952_, _05085_);
  and (_16019_, _15964_, _03137_);
  and (_16020_, _16019_, _16018_);
  or (_16022_, _16020_, _03042_);
  or (_16023_, _16022_, _16017_);
  nor (_16024_, _10365_, _08300_);
  or (_16025_, _15952_, _03043_);
  or (_16026_, _16025_, _16024_);
  and (_16027_, _16026_, _07161_);
  and (_16028_, _16027_, _16023_);
  nor (_16029_, _10367_, _08300_);
  or (_16030_, _16029_, _15952_);
  and (_16031_, _16030_, _03143_);
  or (_16033_, _16031_, _03361_);
  or (_16034_, _16033_, _16028_);
  or (_16035_, _15961_, _03360_);
  and (_16036_, _16035_, _34655_);
  and (_16037_, _16036_, _16034_);
  or (_16038_, _16037_, _15951_);
  and (_35829_[0], _16038_, _35796_);
  not (_16039_, \oc8051_golden_model_1.DPH [1]);
  nor (_16040_, _34655_, _16039_);
  or (_16041_, _10565_, _08300_);
  or (_16043_, _08298_, \oc8051_golden_model_1.DPH [1]);
  and (_16044_, _16043_, _03148_);
  and (_16045_, _16044_, _16041_);
  nor (_16046_, _08324_, \oc8051_golden_model_1.DPH [1]);
  nor (_16047_, _16046_, _08325_);
  and (_16048_, _16047_, _08226_);
  nand (_16049_, _10574_, _04696_);
  and (_16050_, _16049_, _16043_);
  or (_16051_, _16050_, _03006_);
  nand (_16052_, _04696_, _02543_);
  and (_16054_, _16052_, _16043_);
  and (_16055_, _16054_, _03845_);
  nor (_16056_, _03845_, _16039_);
  or (_16057_, _16056_, _02948_);
  or (_16058_, _16057_, _16055_);
  and (_16059_, _16058_, _07474_);
  and (_16060_, _16059_, _16051_);
  nor (_16061_, _08298_, _16039_);
  nor (_16062_, _08300_, _04020_);
  or (_16063_, _16062_, _16061_);
  and (_16065_, _16063_, _02946_);
  or (_16066_, _16065_, _02880_);
  or (_16067_, _16066_, _16060_);
  or (_16068_, _16054_, _02992_);
  and (_16069_, _16068_, _08227_);
  and (_16070_, _16069_, _16067_);
  or (_16071_, _16070_, _16048_);
  and (_16072_, _16071_, _08211_);
  nor (_16073_, _03687_, _08211_);
  or (_16074_, _16073_, _05535_);
  or (_16076_, _16074_, _16072_);
  or (_16077_, _16063_, _02859_);
  and (_16078_, _16077_, _16076_);
  or (_16079_, _16078_, _02841_);
  and (_16080_, _06163_, _08298_);
  or (_16081_, _16061_, _02842_);
  or (_16082_, _16081_, _16080_);
  and (_16083_, _16082_, _02839_);
  and (_16084_, _16083_, _16079_);
  and (_16085_, _16043_, _02567_);
  or (_16087_, _10674_, _08300_);
  and (_16088_, _16087_, _16085_);
  or (_16089_, _16088_, _16084_);
  and (_16090_, _16089_, _03052_);
  or (_16091_, _10689_, _08300_);
  and (_16092_, _16091_, _03051_);
  nand (_16093_, _04696_, _03720_);
  and (_16094_, _16093_, _02834_);
  or (_16095_, _16094_, _16092_);
  and (_16096_, _16095_, _16043_);
  or (_16098_, _16096_, _16090_);
  and (_16099_, _16098_, _07150_);
  or (_16100_, _16099_, _16045_);
  and (_16101_, _16100_, _03138_);
  or (_16102_, _16061_, _05038_);
  and (_16103_, _16054_, _03137_);
  and (_16104_, _16103_, _16102_);
  or (_16105_, _10688_, _08300_);
  and (_16106_, _16043_, _03022_);
  and (_16107_, _16106_, _16105_);
  or (_16109_, _16107_, _16104_);
  or (_16110_, _16109_, _16101_);
  and (_16111_, _16110_, _03144_);
  or (_16112_, _16052_, _05038_);
  and (_16113_, _16043_, _03143_);
  and (_16114_, _16113_, _16112_);
  or (_16115_, _16114_, _03174_);
  or (_16116_, _16093_, _05038_);
  and (_16117_, _16043_, _03042_);
  and (_16118_, _16117_, _16116_);
  or (_16120_, _16118_, _16115_);
  or (_16121_, _16120_, _16111_);
  or (_16122_, _16050_, _03179_);
  and (_16123_, _16122_, _16121_);
  or (_16124_, _16123_, _02887_);
  nor (_16125_, _16061_, _02888_);
  nand (_16126_, _16125_, _16049_);
  and (_16127_, _16126_, _34655_);
  and (_16128_, _16127_, _16124_);
  or (_16129_, _16128_, _16040_);
  and (_35829_[1], _16129_, _35796_);
  not (_16131_, \oc8051_golden_model_1.DPH [2]);
  nor (_16132_, _34655_, _16131_);
  nor (_16133_, _08298_, _16131_);
  nor (_16134_, _10765_, _08300_);
  or (_16135_, _16134_, _16133_);
  and (_16136_, _16135_, _03143_);
  and (_16137_, _10766_, _04696_);
  or (_16138_, _16137_, _16133_);
  and (_16139_, _16138_, _03148_);
  nor (_16141_, _08300_, _04449_);
  or (_16142_, _16141_, _16133_);
  or (_16143_, _16142_, _02859_);
  or (_16144_, _08325_, \oc8051_golden_model_1.DPH [2]);
  nor (_16145_, _08326_, _08227_);
  and (_16146_, _16145_, _16144_);
  nor (_16147_, _10788_, _08300_);
  or (_16148_, _16147_, _16133_);
  or (_16149_, _16148_, _03006_);
  and (_16150_, _08298_, \oc8051_golden_model_1.ACC [2]);
  or (_16152_, _16150_, _16133_);
  and (_16153_, _16152_, _03845_);
  nor (_16154_, _03845_, _16131_);
  or (_16155_, _16154_, _02948_);
  or (_16156_, _16155_, _16153_);
  and (_16157_, _16156_, _07474_);
  and (_16158_, _16157_, _16149_);
  and (_16159_, _16142_, _02946_);
  or (_16160_, _16159_, _02880_);
  or (_16161_, _16160_, _16158_);
  or (_16163_, _16152_, _02992_);
  and (_16164_, _16163_, _08227_);
  and (_16165_, _16164_, _16161_);
  or (_16166_, _16165_, _16146_);
  and (_16167_, _16166_, _08211_);
  nor (_16168_, _03356_, _08211_);
  or (_16169_, _16168_, _05535_);
  or (_16170_, _16169_, _16167_);
  and (_16171_, _16170_, _16143_);
  or (_16172_, _16171_, _02841_);
  or (_16174_, _16133_, _02842_);
  and (_16175_, _06167_, _08298_);
  or (_16176_, _16175_, _16174_);
  and (_16177_, _16176_, _16172_);
  or (_16178_, _16177_, _02567_);
  nor (_16179_, _10881_, _08300_);
  or (_16180_, _16133_, _02839_);
  or (_16181_, _16180_, _16179_);
  and (_16182_, _16181_, _16178_);
  or (_16183_, _16182_, _08207_);
  and (_16185_, _10770_, _04696_);
  or (_16186_, _16133_, _07139_);
  or (_16187_, _16186_, _16185_);
  and (_16188_, _08298_, _05693_);
  or (_16189_, _16188_, _16133_);
  or (_16190_, _16189_, _07140_);
  and (_16191_, _16190_, _07150_);
  and (_16192_, _16191_, _16187_);
  and (_16193_, _16192_, _16183_);
  or (_16194_, _16193_, _16139_);
  and (_16196_, _16194_, _03138_);
  or (_16197_, _16133_, _05135_);
  and (_16198_, _16152_, _03137_);
  and (_16199_, _16189_, _03022_);
  or (_16200_, _16199_, _16198_);
  and (_16201_, _16200_, _16197_);
  or (_16202_, _16201_, _03042_);
  or (_16203_, _16202_, _16196_);
  nor (_16204_, _10768_, _08300_);
  or (_16205_, _16133_, _03043_);
  or (_16207_, _16205_, _16204_);
  and (_16208_, _16207_, _07161_);
  and (_16209_, _16208_, _16203_);
  or (_16210_, _16209_, _16136_);
  and (_16211_, _16210_, _03179_);
  and (_16212_, _16148_, _03174_);
  or (_16213_, _16212_, _02887_);
  or (_16214_, _16213_, _16211_);
  and (_16215_, _10941_, _04696_);
  or (_16216_, _16133_, _02888_);
  or (_16218_, _16216_, _16215_);
  and (_16219_, _16218_, _34655_);
  and (_16220_, _16219_, _16214_);
  or (_16221_, _16220_, _16132_);
  and (_35829_[2], _16221_, _35796_);
  or (_16222_, _34655_, \oc8051_golden_model_1.DPH [3]);
  and (_16223_, _16222_, _35796_);
  not (_16224_, \oc8051_golden_model_1.DPH [3]);
  nor (_16225_, _08298_, _16224_);
  and (_16226_, _10964_, _04696_);
  or (_16228_, _16226_, _16225_);
  and (_16229_, _16228_, _03148_);
  or (_16230_, _08326_, \oc8051_golden_model_1.DPH [3]);
  nor (_16231_, _08327_, _08227_);
  and (_16232_, _16231_, _16230_);
  nor (_16233_, _10983_, _08300_);
  or (_16234_, _16233_, _16225_);
  or (_16235_, _16234_, _03006_);
  and (_16236_, _08298_, \oc8051_golden_model_1.ACC [3]);
  or (_16237_, _16236_, _16225_);
  and (_16239_, _16237_, _03845_);
  nor (_16240_, _03845_, _16224_);
  or (_16241_, _16240_, _02948_);
  or (_16242_, _16241_, _16239_);
  and (_16243_, _16242_, _07474_);
  and (_16244_, _16243_, _16235_);
  nor (_16245_, _08300_, _04275_);
  or (_16246_, _16245_, _16225_);
  and (_16247_, _16246_, _02946_);
  or (_16248_, _16247_, _02880_);
  or (_16250_, _16248_, _16244_);
  or (_16251_, _16237_, _02992_);
  and (_16252_, _16251_, _08227_);
  and (_16253_, _16252_, _16250_);
  or (_16254_, _16253_, _16232_);
  and (_16255_, _16254_, _08211_);
  and (_16256_, _03046_, _02794_);
  or (_16257_, _16256_, _05535_);
  or (_16258_, _16257_, _16255_);
  or (_16259_, _16246_, _02859_);
  and (_16261_, _16259_, _16258_);
  or (_16262_, _16261_, _02841_);
  and (_16263_, _06166_, _08298_);
  or (_16264_, _16225_, _02842_);
  or (_16265_, _16264_, _16263_);
  and (_16266_, _16265_, _02839_);
  and (_16267_, _16266_, _16262_);
  nor (_16268_, _11076_, _08300_);
  or (_16269_, _16268_, _16225_);
  and (_16270_, _16269_, _02567_);
  or (_16272_, _16270_, _08207_);
  or (_16273_, _16272_, _16267_);
  and (_16274_, _10968_, _04696_);
  or (_16275_, _16225_, _07139_);
  or (_16276_, _16275_, _16274_);
  and (_16277_, _08298_, _05654_);
  or (_16278_, _16277_, _16225_);
  or (_16279_, _16278_, _07140_);
  and (_16280_, _16279_, _07150_);
  and (_16281_, _16280_, _16276_);
  and (_16283_, _16281_, _16273_);
  or (_16284_, _16283_, _16229_);
  and (_16285_, _16284_, _03138_);
  or (_16286_, _16225_, _04993_);
  and (_16287_, _16237_, _03137_);
  and (_16288_, _16278_, _03022_);
  or (_16289_, _16288_, _16287_);
  and (_16290_, _16289_, _16286_);
  or (_16291_, _16290_, _03042_);
  or (_16292_, _16291_, _16285_);
  nor (_16294_, _10967_, _08300_);
  or (_16295_, _16225_, _03043_);
  or (_16296_, _16295_, _16294_);
  and (_16297_, _16296_, _07161_);
  and (_16298_, _16297_, _16292_);
  nor (_16299_, _10962_, _08300_);
  or (_16300_, _16299_, _16225_);
  and (_16301_, _16300_, _03143_);
  or (_16302_, _16301_, _03174_);
  or (_16303_, _16302_, _16298_);
  or (_16305_, _16234_, _03179_);
  and (_16306_, _16305_, _02888_);
  and (_16307_, _16306_, _16303_);
  and (_16308_, _11136_, _04696_);
  or (_16309_, _16308_, _16225_);
  and (_16310_, _16309_, _02887_);
  or (_16311_, _16310_, _34659_);
  or (_16312_, _16311_, _16307_);
  and (_35829_[3], _16312_, _16223_);
  or (_16313_, _34655_, \oc8051_golden_model_1.DPH [4]);
  and (_16315_, _16313_, _35796_);
  not (_16316_, \oc8051_golden_model_1.DPH [4]);
  nor (_16317_, _08298_, _16316_);
  nor (_16318_, _05192_, _08300_);
  or (_16319_, _16318_, _16317_);
  or (_16320_, _16319_, _02859_);
  nor (_16321_, _11184_, _08300_);
  or (_16322_, _16321_, _16317_);
  or (_16323_, _16322_, _03006_);
  and (_16324_, _08298_, \oc8051_golden_model_1.ACC [4]);
  or (_16326_, _16324_, _16317_);
  and (_16327_, _16326_, _03845_);
  nor (_16328_, _03845_, _16316_);
  or (_16329_, _16328_, _02948_);
  or (_16330_, _16329_, _16327_);
  and (_16331_, _16330_, _07474_);
  and (_16332_, _16331_, _16323_);
  and (_16333_, _16319_, _02946_);
  or (_16334_, _16333_, _02880_);
  or (_16335_, _16334_, _16332_);
  or (_16337_, _16326_, _02992_);
  and (_16338_, _16337_, _08227_);
  and (_16339_, _16338_, _16335_);
  or (_16340_, _08327_, \oc8051_golden_model_1.DPH [4]);
  nor (_16341_, _08328_, _08227_);
  and (_16342_, _16341_, _16340_);
  or (_16343_, _16342_, _16339_);
  and (_16344_, _16343_, _08211_);
  nor (_16345_, _03647_, _08211_);
  or (_16346_, _16345_, _05535_);
  or (_16348_, _16346_, _16344_);
  and (_16349_, _16348_, _16320_);
  or (_16350_, _16349_, _02841_);
  or (_16351_, _16317_, _02842_);
  and (_16352_, _06171_, _08298_);
  or (_16353_, _16352_, _16351_);
  and (_16354_, _16353_, _16350_);
  or (_16355_, _16354_, _02567_);
  nor (_16356_, _11271_, _08300_);
  or (_16357_, _16317_, _02839_);
  or (_16359_, _16357_, _16356_);
  and (_16360_, _16359_, _16355_);
  or (_16361_, _16360_, _08207_);
  and (_16362_, _11158_, _04696_);
  or (_16363_, _16317_, _07139_);
  or (_16364_, _16363_, _16362_);
  and (_16365_, _05618_, _08298_);
  or (_16366_, _16365_, _16317_);
  or (_16367_, _16366_, _07140_);
  and (_16368_, _16367_, _07150_);
  and (_16370_, _16368_, _16364_);
  and (_16371_, _16370_, _16361_);
  and (_16372_, _11154_, _04696_);
  or (_16373_, _16372_, _16317_);
  and (_16374_, _16373_, _03148_);
  or (_16375_, _16374_, _16371_);
  and (_16376_, _16375_, _03138_);
  or (_16377_, _16317_, _05240_);
  and (_16378_, _16326_, _03137_);
  and (_16379_, _16366_, _03022_);
  or (_16381_, _16379_, _16378_);
  and (_16382_, _16381_, _16377_);
  or (_16383_, _16382_, _03042_);
  or (_16384_, _16383_, _16376_);
  nor (_16385_, _11157_, _08300_);
  or (_16386_, _16317_, _03043_);
  or (_16387_, _16386_, _16385_);
  and (_16388_, _16387_, _07161_);
  and (_16389_, _16388_, _16384_);
  nor (_16390_, _11152_, _08300_);
  or (_16392_, _16390_, _16317_);
  and (_16393_, _16392_, _03143_);
  or (_16394_, _16393_, _03174_);
  or (_16395_, _16394_, _16389_);
  or (_16396_, _16322_, _03179_);
  and (_16397_, _16396_, _02888_);
  and (_16398_, _16397_, _16395_);
  and (_16399_, _11338_, _04696_);
  or (_16400_, _16399_, _16317_);
  and (_16401_, _16400_, _02887_);
  or (_16403_, _16401_, _34659_);
  or (_16404_, _16403_, _16398_);
  and (_35829_[4], _16404_, _16315_);
  or (_16405_, _34655_, \oc8051_golden_model_1.DPH [5]);
  and (_16406_, _16405_, _35796_);
  not (_16407_, \oc8051_golden_model_1.DPH [5]);
  nor (_16408_, _08298_, _16407_);
  nor (_16409_, _04894_, _08300_);
  or (_16410_, _16409_, _16408_);
  or (_16411_, _16410_, _02859_);
  nor (_16413_, _11380_, _08300_);
  or (_16414_, _16413_, _16408_);
  or (_16415_, _16414_, _03006_);
  and (_16416_, _08298_, \oc8051_golden_model_1.ACC [5]);
  or (_16417_, _16416_, _16408_);
  and (_16418_, _16417_, _03845_);
  nor (_16419_, _03845_, _16407_);
  or (_16420_, _16419_, _02948_);
  or (_16421_, _16420_, _16418_);
  and (_16422_, _16421_, _07474_);
  and (_16424_, _16422_, _16415_);
  and (_16425_, _16410_, _02946_);
  or (_16426_, _16425_, _02880_);
  or (_16427_, _16426_, _16424_);
  or (_16428_, _16417_, _02992_);
  and (_16429_, _16428_, _08227_);
  and (_16430_, _16429_, _16427_);
  or (_16431_, _08328_, \oc8051_golden_model_1.DPH [5]);
  nor (_16432_, _08329_, _08227_);
  and (_16433_, _16432_, _16431_);
  or (_16435_, _16433_, _16430_);
  and (_16436_, _16435_, _08211_);
  nor (_16437_, _03220_, _08211_);
  or (_16438_, _16437_, _05535_);
  or (_16439_, _16438_, _16436_);
  and (_16440_, _16439_, _16411_);
  or (_16441_, _16440_, _02841_);
  or (_16442_, _16408_, _02842_);
  and (_16443_, _06170_, _08298_);
  or (_16444_, _16443_, _16442_);
  and (_16447_, _16444_, _16441_);
  or (_16448_, _16447_, _02567_);
  nor (_16449_, _11467_, _08300_);
  or (_16450_, _16408_, _02839_);
  or (_16451_, _16450_, _16449_);
  and (_16452_, _16451_, _16448_);
  or (_16453_, _16452_, _08207_);
  and (_16454_, _11482_, _04696_);
  or (_16455_, _16408_, _07139_);
  or (_16456_, _16455_, _16454_);
  and (_16458_, _05671_, _08298_);
  or (_16459_, _16458_, _16408_);
  or (_16460_, _16459_, _07140_);
  and (_16461_, _16460_, _07150_);
  and (_16462_, _16461_, _16456_);
  and (_16463_, _16462_, _16453_);
  and (_16464_, _11356_, _04696_);
  or (_16465_, _16464_, _16408_);
  and (_16466_, _16465_, _03148_);
  or (_16467_, _16466_, _16463_);
  and (_16469_, _16467_, _03138_);
  or (_16470_, _16408_, _04945_);
  and (_16471_, _16417_, _03137_);
  and (_16472_, _16459_, _03022_);
  or (_16473_, _16472_, _16471_);
  and (_16474_, _16473_, _16470_);
  or (_16475_, _16474_, _03042_);
  or (_16476_, _16475_, _16469_);
  nor (_16477_, _11480_, _08300_);
  or (_16478_, _16408_, _03043_);
  or (_16480_, _16478_, _16477_);
  and (_16481_, _16480_, _07161_);
  and (_16482_, _16481_, _16476_);
  nor (_16483_, _11355_, _08300_);
  or (_16484_, _16483_, _16408_);
  and (_16485_, _16484_, _03143_);
  or (_16486_, _16485_, _03174_);
  or (_16487_, _16486_, _16482_);
  or (_16488_, _16414_, _03179_);
  and (_16489_, _16488_, _02888_);
  and (_16491_, _16489_, _16487_);
  and (_16492_, _11541_, _04696_);
  or (_16493_, _16492_, _16408_);
  and (_16494_, _16493_, _02887_);
  or (_16495_, _16494_, _34659_);
  or (_16496_, _16495_, _16491_);
  and (_35829_[5], _16496_, _16406_);
  or (_16497_, _34655_, \oc8051_golden_model_1.DPH [6]);
  and (_16498_, _16497_, _35796_);
  not (_16499_, \oc8051_golden_model_1.DPH [6]);
  nor (_16501_, _08298_, _16499_);
  nor (_16502_, _04790_, _08300_);
  or (_16503_, _16502_, _16501_);
  or (_16504_, _16503_, _02859_);
  nor (_16505_, _11567_, _08300_);
  or (_16506_, _16505_, _16501_);
  or (_16507_, _16506_, _03006_);
  and (_16508_, _08298_, \oc8051_golden_model_1.ACC [6]);
  or (_16509_, _16508_, _16501_);
  and (_16510_, _16509_, _03845_);
  nor (_16512_, _03845_, _16499_);
  or (_16513_, _16512_, _02948_);
  or (_16514_, _16513_, _16510_);
  and (_16515_, _16514_, _07474_);
  and (_16516_, _16515_, _16507_);
  and (_16517_, _16503_, _02946_);
  or (_16518_, _16517_, _02880_);
  or (_16519_, _16518_, _16516_);
  or (_16520_, _16509_, _02992_);
  and (_16521_, _16520_, _08227_);
  and (_16523_, _16521_, _16519_);
  or (_16524_, _08329_, \oc8051_golden_model_1.DPH [6]);
  nor (_16525_, _08330_, _08227_);
  and (_16526_, _16525_, _16524_);
  or (_16527_, _16526_, _16523_);
  and (_16528_, _16527_, _08211_);
  nor (_16529_, _08211_, _02924_);
  or (_16530_, _16529_, _05535_);
  or (_16531_, _16530_, _16528_);
  and (_16532_, _16531_, _16504_);
  or (_16534_, _16532_, _02841_);
  or (_16535_, _16501_, _02842_);
  and (_16536_, _06162_, _08298_);
  or (_16537_, _16536_, _16535_);
  and (_16538_, _16537_, _16534_);
  or (_16539_, _16538_, _02567_);
  nor (_16540_, _11671_, _08300_);
  or (_16541_, _16501_, _02839_);
  or (_16542_, _16541_, _16540_);
  and (_16543_, _16542_, _16539_);
  or (_16545_, _16543_, _08207_);
  and (_16546_, _11560_, _04696_);
  or (_16547_, _16501_, _07139_);
  or (_16548_, _16547_, _16546_);
  and (_16549_, _11678_, _08298_);
  or (_16550_, _16549_, _16501_);
  or (_16551_, _16550_, _07140_);
  and (_16552_, _16551_, _07150_);
  and (_16553_, _16552_, _16548_);
  and (_16554_, _16553_, _16545_);
  and (_16556_, _11556_, _04696_);
  or (_16557_, _16556_, _16501_);
  and (_16558_, _16557_, _03148_);
  or (_16559_, _16558_, _16554_);
  and (_16560_, _16559_, _03138_);
  or (_16561_, _16501_, _04838_);
  and (_16562_, _16509_, _03137_);
  and (_16563_, _16550_, _03022_);
  or (_16564_, _16563_, _16562_);
  and (_16565_, _16564_, _16561_);
  or (_16567_, _16565_, _03042_);
  or (_16568_, _16567_, _16560_);
  nor (_16569_, _11558_, _08300_);
  or (_16570_, _16501_, _03043_);
  or (_16571_, _16570_, _16569_);
  and (_16572_, _16571_, _07161_);
  and (_16573_, _16572_, _16568_);
  nor (_16574_, _11555_, _08300_);
  or (_16575_, _16574_, _16501_);
  and (_16576_, _16575_, _03143_);
  or (_16578_, _16576_, _03174_);
  or (_16579_, _16578_, _16573_);
  or (_16580_, _16506_, _03179_);
  and (_16581_, _16580_, _02888_);
  and (_16582_, _16581_, _16579_);
  and (_16583_, _11744_, _04696_);
  or (_16584_, _16583_, _16501_);
  and (_16585_, _16584_, _02887_);
  or (_16586_, _16585_, _34659_);
  or (_16587_, _16586_, _16582_);
  and (_35829_[6], _16587_, _16498_);
  and (_35831_[0], \oc8051_golden_model_1.IE [0], _35796_);
  and (_35831_[1], \oc8051_golden_model_1.IE [1], _35796_);
  and (_35831_[2], \oc8051_golden_model_1.IE [2], _35796_);
  and (_35831_[3], \oc8051_golden_model_1.IE [3], _35796_);
  and (_35831_[4], \oc8051_golden_model_1.IE [4], _35796_);
  and (_35831_[5], \oc8051_golden_model_1.IE [5], _35796_);
  and (_35831_[6], \oc8051_golden_model_1.IE [6], _35796_);
  and (_35832_[0], \oc8051_golden_model_1.IP [0], _35796_);
  and (_35832_[1], \oc8051_golden_model_1.IP [1], _35796_);
  and (_35832_[2], \oc8051_golden_model_1.IP [2], _35796_);
  and (_35832_[3], \oc8051_golden_model_1.IP [3], _35796_);
  and (_35832_[4], \oc8051_golden_model_1.IP [4], _35796_);
  and (_35832_[5], \oc8051_golden_model_1.IP [5], _35796_);
  and (_35832_[6], \oc8051_golden_model_1.IP [6], _35796_);
  not (_16590_, \oc8051_golden_model_1.P0 [0]);
  nor (_16591_, _34655_, _16590_);
  or (_16592_, _16591_, rst);
  nor (_16593_, _04654_, _16590_);
  and (_16594_, _10369_, _04654_);
  or (_16596_, _16594_, _16593_);
  and (_16597_, _16596_, _03148_);
  and (_16598_, _04654_, _03838_);
  or (_16599_, _16598_, _16593_);
  or (_16600_, _16599_, _02859_);
  nor (_16601_, _04635_, _16590_);
  and (_16602_, _10390_, _04635_);
  or (_16603_, _16602_, _16601_);
  and (_16604_, _16603_, _02884_);
  nor (_16605_, _05085_, _08393_);
  or (_16607_, _16605_, _16593_);
  or (_16608_, _16607_, _03006_);
  and (_16609_, _04654_, \oc8051_golden_model_1.ACC [0]);
  or (_16610_, _16609_, _16593_);
  and (_16611_, _16610_, _03845_);
  nor (_16612_, _03845_, _16590_);
  or (_16613_, _16612_, _02948_);
  or (_16614_, _16613_, _16611_);
  and (_16615_, _16614_, _02976_);
  and (_16616_, _16615_, _16608_);
  and (_16618_, _16599_, _02946_);
  or (_16619_, _16618_, _02880_);
  or (_16620_, _16619_, _16616_);
  or (_16621_, _16620_, _16604_);
  or (_16622_, _16610_, _02992_);
  and (_16623_, _16622_, _02987_);
  and (_16624_, _16623_, _16621_);
  and (_16625_, _16593_, _02877_);
  or (_16626_, _16625_, _02871_);
  or (_16627_, _16626_, _16624_);
  or (_16629_, _16607_, _06246_);
  and (_16630_, _16629_, _02986_);
  and (_16631_, _16630_, _16627_);
  or (_16632_, _10399_, _10376_);
  and (_16633_, _16632_, _04635_);
  or (_16634_, _16633_, _16601_);
  and (_16635_, _16634_, _02866_);
  or (_16636_, _16635_, _05535_);
  or (_16637_, _16636_, _16631_);
  and (_16638_, _16637_, _16600_);
  or (_16640_, _16638_, _02841_);
  and (_16641_, _06164_, _04654_);
  or (_16642_, _16593_, _02842_);
  or (_16643_, _16642_, _16641_);
  and (_16644_, _16643_, _02839_);
  and (_16645_, _16644_, _16640_);
  nor (_16646_, _10475_, _08393_);
  or (_16647_, _16646_, _16593_);
  and (_16648_, _16647_, _02567_);
  or (_16649_, _16648_, _08207_);
  or (_16651_, _16649_, _16645_);
  and (_16652_, _10372_, _04654_);
  or (_16653_, _16593_, _07139_);
  or (_16654_, _16653_, _16652_);
  and (_16655_, _04654_, _05660_);
  or (_16656_, _16655_, _16593_);
  or (_16657_, _16656_, _07140_);
  and (_16658_, _16657_, _07150_);
  and (_16659_, _16658_, _16654_);
  and (_16660_, _16659_, _16651_);
  or (_16662_, _16660_, _16597_);
  and (_16663_, _16662_, _03138_);
  nand (_16664_, _16656_, _03022_);
  nor (_16665_, _16664_, _16605_);
  or (_16666_, _16593_, _05085_);
  and (_16667_, _16610_, _03137_);
  and (_16668_, _16667_, _16666_);
  or (_16669_, _16668_, _03042_);
  or (_16670_, _16669_, _16665_);
  or (_16671_, _16670_, _16663_);
  nor (_16673_, _10365_, _08393_);
  or (_16674_, _16593_, _03043_);
  or (_16675_, _16674_, _16673_);
  and (_16676_, _16675_, _07161_);
  and (_16677_, _16676_, _16671_);
  nor (_16678_, _10367_, _08393_);
  or (_16679_, _16678_, _16593_);
  and (_16680_, _16679_, _03143_);
  or (_16681_, _16680_, _03174_);
  or (_16682_, _16681_, _16677_);
  or (_16684_, _16607_, _03179_);
  and (_16685_, _16684_, _03183_);
  and (_16686_, _16685_, _16682_);
  and (_16687_, _16593_, _02799_);
  or (_16688_, _16687_, _02887_);
  or (_16689_, _16688_, _16686_);
  or (_16690_, _16607_, _02888_);
  and (_16691_, _16690_, _34655_);
  and (_16692_, _16691_, _16689_);
  or (_35834_[0], _16692_, _16592_);
  not (_16694_, \oc8051_golden_model_1.P0 [1]);
  nor (_16695_, _34655_, _16694_);
  or (_16696_, _16695_, rst);
  or (_16697_, _10565_, _08393_);
  or (_16698_, _04654_, \oc8051_golden_model_1.P0 [1]);
  and (_16699_, _16698_, _03148_);
  and (_16700_, _16699_, _16697_);
  or (_16701_, _10617_, _10572_);
  and (_16702_, _16701_, _04635_);
  nor (_16703_, _04635_, _16694_);
  or (_16705_, _16703_, _02986_);
  or (_16706_, _16705_, _16702_);
  and (_16707_, _10574_, _04654_);
  not (_16708_, _16707_);
  and (_16709_, _16708_, _16698_);
  or (_16710_, _16709_, _03006_);
  nand (_16711_, _04654_, _02543_);
  and (_16712_, _16711_, _16698_);
  and (_16713_, _16712_, _03845_);
  nor (_16714_, _03845_, _16694_);
  or (_16716_, _16714_, _02948_);
  or (_16717_, _16716_, _16713_);
  and (_16718_, _16717_, _02976_);
  and (_16719_, _16718_, _16710_);
  nor (_16720_, _04654_, _16694_);
  nor (_16721_, _08393_, _04020_);
  or (_16722_, _16721_, _16720_);
  and (_16723_, _16722_, _02946_);
  and (_16724_, _10569_, _04635_);
  or (_16725_, _16724_, _16703_);
  and (_16727_, _16725_, _02884_);
  or (_16728_, _16727_, _16723_);
  or (_16729_, _16728_, _02880_);
  or (_16730_, _16729_, _16719_);
  or (_16731_, _16712_, _02992_);
  and (_16732_, _16731_, _16730_);
  or (_16733_, _16732_, _02877_);
  and (_16734_, _10572_, _04635_);
  or (_16735_, _16734_, _16703_);
  or (_16736_, _16735_, _02987_);
  and (_16738_, _16736_, _06246_);
  and (_16739_, _16738_, _16733_);
  and (_16740_, _16724_, _10568_);
  or (_16741_, _16740_, _16703_);
  and (_16742_, _16741_, _02871_);
  or (_16743_, _16742_, _02866_);
  or (_16744_, _16743_, _16739_);
  and (_16745_, _16744_, _16706_);
  or (_16746_, _16745_, _05535_);
  or (_16747_, _16722_, _02859_);
  and (_16749_, _16747_, _16746_);
  or (_16750_, _16749_, _02841_);
  and (_16751_, _06163_, _04654_);
  or (_16752_, _16720_, _02842_);
  or (_16753_, _16752_, _16751_);
  and (_16754_, _16753_, _02839_);
  and (_16755_, _16754_, _16750_);
  and (_16756_, _10674_, _04654_);
  or (_16757_, _16756_, _16720_);
  and (_16758_, _16757_, _02567_);
  or (_16760_, _16758_, _16755_);
  and (_16761_, _16760_, _03052_);
  or (_16762_, _10689_, _08393_);
  and (_16763_, _16762_, _03051_);
  nand (_16764_, _04654_, _03720_);
  and (_16765_, _16764_, _02834_);
  or (_16766_, _16765_, _16763_);
  and (_16767_, _16766_, _16698_);
  or (_16768_, _16767_, _16761_);
  and (_16769_, _16768_, _07150_);
  or (_16771_, _16769_, _16700_);
  and (_16772_, _16771_, _03138_);
  or (_16773_, _10688_, _08393_);
  and (_16774_, _16698_, _03022_);
  and (_16775_, _16774_, _16773_);
  or (_16776_, _16720_, _05038_);
  and (_16777_, _16712_, _03137_);
  and (_16778_, _16777_, _16776_);
  or (_16779_, _16778_, _16775_);
  or (_16780_, _16779_, _16772_);
  and (_16782_, _16780_, _03144_);
  or (_16783_, _16764_, _05038_);
  and (_16784_, _16698_, _03042_);
  and (_16785_, _16784_, _16783_);
  or (_16786_, _16711_, _05038_);
  and (_16787_, _16698_, _03143_);
  and (_16788_, _16787_, _16786_);
  or (_16789_, _16788_, _03174_);
  or (_16790_, _16789_, _16785_);
  or (_16791_, _16790_, _16782_);
  or (_16793_, _16709_, _03179_);
  and (_16794_, _16793_, _03183_);
  and (_16795_, _16794_, _16791_);
  and (_16796_, _16735_, _02799_);
  or (_16797_, _16796_, _02887_);
  or (_16798_, _16797_, _16795_);
  or (_16799_, _16720_, _02888_);
  or (_16800_, _16799_, _16707_);
  and (_16801_, _16800_, _34655_);
  and (_16802_, _16801_, _16798_);
  or (_35834_[1], _16802_, _16696_);
  not (_16804_, \oc8051_golden_model_1.P0 [2]);
  nor (_16805_, _34655_, _16804_);
  or (_16806_, _16805_, rst);
  nor (_16807_, _04654_, _16804_);
  nor (_16808_, _08393_, _04449_);
  or (_16809_, _16808_, _16807_);
  or (_16810_, _16809_, _02859_);
  and (_16811_, _04654_, \oc8051_golden_model_1.ACC [2]);
  or (_16812_, _16811_, _16807_);
  or (_16814_, _16812_, _02992_);
  nor (_16815_, _10788_, _08393_);
  or (_16816_, _16815_, _16807_);
  or (_16817_, _16816_, _03006_);
  and (_16818_, _16812_, _03845_);
  nor (_16819_, _03845_, _16804_);
  or (_16820_, _16819_, _02948_);
  or (_16821_, _16820_, _16818_);
  and (_16822_, _16821_, _02976_);
  and (_16823_, _16822_, _16817_);
  nor (_16825_, _04635_, _16804_);
  and (_16826_, _10792_, _04635_);
  or (_16827_, _16826_, _16825_);
  and (_16828_, _16827_, _02884_);
  and (_16829_, _16809_, _02946_);
  or (_16830_, _16829_, _02880_);
  or (_16831_, _16830_, _16828_);
  or (_16832_, _16831_, _16823_);
  and (_16833_, _16832_, _16814_);
  or (_16834_, _16833_, _02877_);
  and (_16836_, _10773_, _04635_);
  or (_16837_, _16836_, _16825_);
  or (_16838_, _16837_, _02987_);
  and (_16839_, _16838_, _06246_);
  and (_16840_, _16839_, _16834_);
  or (_16841_, _16825_, _10807_);
  and (_16842_, _16841_, _16827_);
  and (_16843_, _16842_, _02871_);
  or (_16844_, _16843_, _16840_);
  and (_16845_, _16844_, _02986_);
  or (_16847_, _10824_, _10773_);
  and (_16848_, _16847_, _04635_);
  or (_16849_, _16825_, _16848_);
  and (_16850_, _16849_, _02866_);
  or (_16851_, _16850_, _05535_);
  or (_16852_, _16851_, _16845_);
  and (_16853_, _16852_, _16810_);
  or (_16854_, _16853_, _02841_);
  and (_16855_, _06167_, _04654_);
  or (_16856_, _16807_, _02842_);
  or (_16858_, _16856_, _16855_);
  and (_16859_, _16858_, _02839_);
  and (_16860_, _16859_, _16854_);
  nor (_16861_, _10881_, _08393_);
  or (_16862_, _16861_, _16807_);
  and (_16863_, _16862_, _02567_);
  or (_16864_, _16863_, _16860_);
  or (_16865_, _16864_, _08207_);
  and (_16866_, _10770_, _04654_);
  or (_16867_, _16807_, _07139_);
  or (_16869_, _16867_, _16866_);
  and (_16870_, _04654_, _05693_);
  or (_16871_, _16870_, _16807_);
  or (_16872_, _16871_, _07140_);
  and (_16873_, _16872_, _07150_);
  and (_16874_, _16873_, _16869_);
  and (_16875_, _16874_, _16865_);
  and (_16876_, _10766_, _04654_);
  or (_16877_, _16876_, _16807_);
  and (_16878_, _16877_, _03148_);
  or (_16880_, _16878_, _16875_);
  and (_16881_, _16880_, _03138_);
  or (_16882_, _16807_, _05135_);
  and (_16883_, _16812_, _03137_);
  and (_16884_, _16871_, _03022_);
  or (_16885_, _16884_, _16883_);
  and (_16886_, _16885_, _16882_);
  or (_16887_, _16886_, _03042_);
  or (_16888_, _16887_, _16881_);
  nor (_16889_, _10768_, _08393_);
  or (_16891_, _16807_, _03043_);
  or (_16892_, _16891_, _16889_);
  and (_16893_, _16892_, _07161_);
  and (_16894_, _16893_, _16888_);
  nor (_16895_, _10765_, _08393_);
  or (_16896_, _16895_, _16807_);
  and (_16897_, _16896_, _03143_);
  or (_16898_, _16897_, _03174_);
  or (_16899_, _16898_, _16894_);
  or (_16900_, _16816_, _03179_);
  and (_16902_, _16900_, _03183_);
  and (_16903_, _16902_, _16899_);
  and (_16904_, _16837_, _02799_);
  or (_16905_, _16904_, _02887_);
  or (_16906_, _16905_, _16903_);
  and (_16907_, _10941_, _04654_);
  or (_16908_, _16807_, _02888_);
  or (_16909_, _16908_, _16907_);
  and (_16910_, _16909_, _34655_);
  and (_16911_, _16910_, _16906_);
  or (_35834_[2], _16911_, _16806_);
  not (_16913_, \oc8051_golden_model_1.P0 [3]);
  nor (_16914_, _34655_, _16913_);
  or (_16915_, _16914_, rst);
  nor (_16916_, _04654_, _16913_);
  nor (_16917_, _08393_, _04275_);
  or (_16918_, _16917_, _16916_);
  or (_16919_, _16918_, _02859_);
  or (_16920_, _10979_, _10971_);
  and (_16921_, _16920_, _04635_);
  nor (_16923_, _04635_, _16913_);
  or (_16924_, _16923_, _02986_);
  or (_16925_, _16924_, _16921_);
  nor (_16926_, _10983_, _08393_);
  or (_16927_, _16926_, _16916_);
  or (_16928_, _16927_, _03006_);
  and (_16929_, _04654_, \oc8051_golden_model_1.ACC [3]);
  or (_16930_, _16929_, _16916_);
  and (_16931_, _16930_, _03845_);
  nor (_16932_, _03845_, _16913_);
  or (_16934_, _16932_, _02948_);
  or (_16935_, _16934_, _16931_);
  and (_16936_, _16935_, _02976_);
  and (_16937_, _16936_, _16928_);
  and (_16938_, _16918_, _02946_);
  and (_16939_, _10976_, _04635_);
  or (_16940_, _16939_, _16923_);
  and (_16941_, _16940_, _02884_);
  or (_16942_, _16941_, _16938_);
  or (_16943_, _16942_, _02880_);
  or (_16945_, _16943_, _16937_);
  or (_16946_, _16930_, _02992_);
  and (_16947_, _16946_, _16945_);
  or (_16948_, _16947_, _02877_);
  and (_16949_, _10979_, _04635_);
  or (_16950_, _16949_, _16923_);
  or (_16951_, _16950_, _02987_);
  and (_16952_, _16951_, _06246_);
  and (_16953_, _16952_, _16948_);
  or (_16954_, _16923_, _10975_);
  and (_16956_, _16954_, _02871_);
  and (_16957_, _16956_, _16940_);
  or (_16958_, _16957_, _02866_);
  or (_16959_, _16958_, _16953_);
  and (_16960_, _16959_, _16925_);
  or (_16961_, _16960_, _05535_);
  and (_16962_, _16961_, _16919_);
  or (_16963_, _16962_, _02841_);
  and (_16964_, _06166_, _04654_);
  or (_16965_, _16916_, _02842_);
  or (_16967_, _16965_, _16964_);
  and (_16968_, _16967_, _02839_);
  and (_16969_, _16968_, _16963_);
  nor (_16970_, _11076_, _08393_);
  or (_16971_, _16916_, _16970_);
  and (_16972_, _16971_, _02567_);
  or (_16973_, _16972_, _16969_);
  or (_16974_, _16973_, _08207_);
  and (_16975_, _10968_, _04654_);
  or (_16976_, _16916_, _07139_);
  or (_16978_, _16976_, _16975_);
  and (_16979_, _04654_, _05654_);
  or (_16980_, _16979_, _16916_);
  or (_16981_, _16980_, _07140_);
  and (_16982_, _16981_, _07150_);
  and (_16983_, _16982_, _16978_);
  and (_16984_, _16983_, _16974_);
  and (_16985_, _10964_, _04654_);
  or (_16986_, _16985_, _16916_);
  and (_16987_, _16986_, _03148_);
  or (_16989_, _16987_, _16984_);
  and (_16990_, _16989_, _03138_);
  or (_16991_, _16916_, _04993_);
  and (_16992_, _16930_, _03137_);
  and (_16993_, _16980_, _03022_);
  or (_16994_, _16993_, _16992_);
  and (_16995_, _16994_, _16991_);
  or (_16996_, _16995_, _03042_);
  or (_16997_, _16996_, _16990_);
  nor (_16998_, _10967_, _08393_);
  or (_17000_, _16916_, _03043_);
  or (_17001_, _17000_, _16998_);
  and (_17002_, _17001_, _07161_);
  and (_17003_, _17002_, _16997_);
  nor (_17004_, _10962_, _08393_);
  or (_17005_, _17004_, _16916_);
  and (_17006_, _17005_, _03143_);
  or (_17007_, _17006_, _03174_);
  or (_17008_, _17007_, _17003_);
  or (_17009_, _16927_, _03179_);
  and (_17011_, _17009_, _03183_);
  and (_17012_, _17011_, _17008_);
  and (_17013_, _16950_, _02799_);
  or (_17014_, _17013_, _02887_);
  or (_17015_, _17014_, _17012_);
  and (_17016_, _11136_, _04654_);
  or (_17017_, _16916_, _02888_);
  or (_17018_, _17017_, _17016_);
  and (_17019_, _17018_, _34655_);
  and (_17020_, _17019_, _17015_);
  or (_35834_[3], _17020_, _16915_);
  not (_17022_, \oc8051_golden_model_1.P0 [4]);
  nor (_17023_, _34655_, _17022_);
  or (_17024_, _17023_, rst);
  nor (_17025_, _04654_, _17022_);
  nor (_17026_, _05192_, _08393_);
  or (_17027_, _17026_, _17025_);
  or (_17028_, _17027_, _02859_);
  nor (_17029_, _04635_, _17022_);
  and (_17030_, _11167_, _04635_);
  or (_17032_, _17030_, _17029_);
  or (_17033_, _17029_, _11201_);
  and (_17034_, _17033_, _02871_);
  and (_17035_, _17034_, _17032_);
  nor (_17036_, _11184_, _08393_);
  or (_17037_, _17036_, _17025_);
  or (_17038_, _17037_, _03006_);
  and (_17039_, _04654_, \oc8051_golden_model_1.ACC [4]);
  or (_17040_, _17039_, _17025_);
  and (_17041_, _17040_, _03845_);
  nor (_17043_, _03845_, _17022_);
  or (_17044_, _17043_, _02948_);
  or (_17045_, _17044_, _17041_);
  and (_17046_, _17045_, _02976_);
  and (_17047_, _17046_, _17038_);
  and (_17048_, _17027_, _02946_);
  and (_17049_, _17032_, _02884_);
  or (_17050_, _17049_, _17048_);
  or (_17051_, _17050_, _02880_);
  or (_17052_, _17051_, _17047_);
  or (_17054_, _17040_, _02992_);
  and (_17055_, _17054_, _17052_);
  or (_17056_, _17055_, _02877_);
  and (_17057_, _11165_, _04635_);
  or (_17058_, _17057_, _17029_);
  or (_17059_, _17058_, _02987_);
  and (_17060_, _17059_, _06246_);
  and (_17061_, _17060_, _17056_);
  or (_17062_, _17061_, _17035_);
  and (_17063_, _17062_, _02986_);
  or (_17065_, _11165_, _11162_);
  and (_17066_, _17065_, _04635_);
  or (_17067_, _17066_, _17029_);
  and (_17068_, _17067_, _02866_);
  or (_17069_, _17068_, _05535_);
  or (_17070_, _17069_, _17063_);
  and (_17071_, _17070_, _17028_);
  or (_17072_, _17071_, _02841_);
  and (_17073_, _06171_, _04654_);
  or (_17074_, _17025_, _02842_);
  or (_17076_, _17074_, _17073_);
  and (_17077_, _17076_, _02839_);
  and (_17078_, _17077_, _17072_);
  nor (_17079_, _11271_, _08393_);
  or (_17080_, _17079_, _17025_);
  and (_17081_, _17080_, _02567_);
  or (_17082_, _17081_, _17078_);
  or (_17083_, _17082_, _08207_);
  and (_17084_, _11158_, _04654_);
  or (_17085_, _17025_, _07139_);
  or (_17087_, _17085_, _17084_);
  and (_17088_, _05618_, _04654_);
  or (_17089_, _17088_, _17025_);
  or (_17090_, _17089_, _07140_);
  and (_17091_, _17090_, _07150_);
  and (_17092_, _17091_, _17087_);
  and (_17093_, _17092_, _17083_);
  and (_17094_, _11154_, _04654_);
  or (_17095_, _17094_, _17025_);
  and (_17096_, _17095_, _03148_);
  or (_17098_, _17096_, _17093_);
  and (_17099_, _17098_, _03138_);
  or (_17100_, _17025_, _05240_);
  and (_17101_, _17040_, _03137_);
  and (_17102_, _17089_, _03022_);
  or (_17103_, _17102_, _17101_);
  and (_17104_, _17103_, _17100_);
  or (_17105_, _17104_, _03042_);
  or (_17106_, _17105_, _17099_);
  nor (_17107_, _11157_, _08393_);
  or (_17109_, _17025_, _03043_);
  or (_17110_, _17109_, _17107_);
  and (_17111_, _17110_, _07161_);
  and (_17112_, _17111_, _17106_);
  nor (_17113_, _11152_, _08393_);
  or (_17114_, _17113_, _17025_);
  and (_17115_, _17114_, _03143_);
  or (_17116_, _17115_, _03174_);
  or (_17117_, _17116_, _17112_);
  or (_17118_, _17037_, _03179_);
  and (_17120_, _17118_, _03183_);
  and (_17121_, _17120_, _17117_);
  and (_17122_, _17058_, _02799_);
  or (_17123_, _17122_, _02887_);
  or (_17124_, _17123_, _17121_);
  and (_17125_, _11338_, _04654_);
  or (_17126_, _17025_, _02888_);
  or (_17127_, _17126_, _17125_);
  and (_17128_, _17127_, _34655_);
  and (_17129_, _17128_, _17124_);
  or (_35834_[4], _17129_, _17024_);
  not (_17131_, \oc8051_golden_model_1.P0 [5]);
  nor (_17132_, _34655_, _17131_);
  or (_17133_, _17132_, rst);
  nor (_17134_, _04654_, _17131_);
  nor (_17135_, _11380_, _08393_);
  or (_17136_, _17135_, _17134_);
  or (_17137_, _17136_, _03006_);
  and (_17138_, _04654_, \oc8051_golden_model_1.ACC [5]);
  or (_17139_, _17138_, _17134_);
  and (_17140_, _17139_, _03845_);
  nor (_17141_, _03845_, _17131_);
  or (_17142_, _17141_, _02948_);
  or (_17143_, _17142_, _17140_);
  and (_17144_, _17143_, _02976_);
  and (_17145_, _17144_, _17137_);
  nor (_17146_, _04894_, _08393_);
  or (_17147_, _17146_, _17134_);
  and (_17148_, _17147_, _02946_);
  nor (_17149_, _04635_, _17131_);
  and (_17152_, _11365_, _04635_);
  or (_17153_, _17152_, _17149_);
  and (_17154_, _17153_, _02884_);
  or (_17155_, _17154_, _17148_);
  or (_17156_, _17155_, _02880_);
  or (_17157_, _17156_, _17145_);
  or (_17158_, _17139_, _02992_);
  and (_17159_, _17158_, _17157_);
  or (_17160_, _17159_, _02877_);
  and (_17161_, _11363_, _04635_);
  or (_17162_, _17161_, _17149_);
  or (_17163_, _17162_, _02987_);
  and (_17164_, _17163_, _06246_);
  and (_17165_, _17164_, _17160_);
  and (_17166_, _11398_, _04635_);
  or (_17167_, _17166_, _17149_);
  and (_17168_, _17167_, _02871_);
  or (_17169_, _17168_, _17165_);
  and (_17170_, _17169_, _02986_);
  or (_17171_, _11363_, _11360_);
  and (_17174_, _17171_, _04635_);
  or (_17175_, _17174_, _17149_);
  and (_17176_, _17175_, _02866_);
  or (_17177_, _17176_, _05535_);
  or (_17178_, _17177_, _17170_);
  or (_17179_, _17147_, _02859_);
  and (_17180_, _17179_, _17178_);
  or (_17181_, _17180_, _02841_);
  and (_17182_, _06170_, _04654_);
  or (_17183_, _17134_, _02842_);
  or (_17185_, _17183_, _17182_);
  and (_17186_, _17185_, _02839_);
  and (_17187_, _17186_, _17181_);
  nor (_17188_, _11467_, _08393_);
  or (_17189_, _17188_, _17134_);
  and (_17190_, _17189_, _02567_);
  or (_17191_, _17190_, _08207_);
  or (_17192_, _17191_, _17187_);
  and (_17193_, _11482_, _04654_);
  or (_17194_, _17134_, _07139_);
  or (_17196_, _17194_, _17193_);
  and (_17197_, _05671_, _04654_);
  or (_17198_, _17197_, _17134_);
  or (_17199_, _17198_, _07140_);
  and (_17200_, _17199_, _07150_);
  and (_17201_, _17200_, _17196_);
  and (_17202_, _17201_, _17192_);
  and (_17203_, _11356_, _04654_);
  or (_17204_, _17203_, _17134_);
  and (_17205_, _17204_, _03148_);
  or (_17207_, _17205_, _17202_);
  and (_17208_, _17207_, _03138_);
  or (_17209_, _17134_, _04945_);
  and (_17210_, _17139_, _03137_);
  and (_17211_, _17198_, _03022_);
  or (_17212_, _17211_, _17210_);
  and (_17213_, _17212_, _17209_);
  or (_17214_, _17213_, _03042_);
  or (_17215_, _17214_, _17208_);
  nor (_17216_, _11480_, _08393_);
  or (_17218_, _17134_, _03043_);
  or (_17219_, _17218_, _17216_);
  and (_17220_, _17219_, _07161_);
  and (_17221_, _17220_, _17215_);
  nor (_17222_, _11355_, _08393_);
  or (_17223_, _17222_, _17134_);
  and (_17224_, _17223_, _03143_);
  or (_17225_, _17224_, _03174_);
  or (_17226_, _17225_, _17221_);
  or (_17227_, _17136_, _03179_);
  and (_17229_, _17227_, _03183_);
  and (_17230_, _17229_, _17226_);
  and (_17231_, _17162_, _02799_);
  or (_17232_, _17231_, _02887_);
  or (_17233_, _17232_, _17230_);
  and (_17234_, _11541_, _04654_);
  or (_17235_, _17134_, _02888_);
  or (_17236_, _17235_, _17234_);
  and (_17237_, _17236_, _34655_);
  and (_17238_, _17237_, _17233_);
  or (_35834_[5], _17238_, _17133_);
  not (_17240_, \oc8051_golden_model_1.P0 [6]);
  nor (_17241_, _34655_, _17240_);
  or (_17242_, _17241_, rst);
  nor (_17243_, _04635_, _17240_);
  and (_17244_, _11564_, _04635_);
  or (_17245_, _17244_, _17243_);
  or (_17246_, _17243_, _11596_);
  and (_17247_, _17246_, _02871_);
  and (_17248_, _17247_, _17245_);
  nor (_17250_, _04654_, _17240_);
  nor (_17251_, _11567_, _08393_);
  or (_17252_, _17251_, _17250_);
  or (_17253_, _17252_, _03006_);
  and (_17254_, _04654_, \oc8051_golden_model_1.ACC [6]);
  or (_17255_, _17254_, _17250_);
  and (_17256_, _17255_, _03845_);
  nor (_17257_, _03845_, _17240_);
  or (_17258_, _17257_, _02948_);
  or (_17259_, _17258_, _17256_);
  and (_17261_, _17259_, _02976_);
  and (_17262_, _17261_, _17253_);
  nor (_17263_, _04790_, _08393_);
  or (_17264_, _17263_, _17250_);
  and (_17265_, _17264_, _02946_);
  and (_17266_, _17245_, _02884_);
  or (_17267_, _17266_, _17265_);
  or (_17268_, _17267_, _02880_);
  or (_17269_, _17268_, _17262_);
  or (_17270_, _17255_, _02992_);
  and (_17272_, _17270_, _17269_);
  or (_17273_, _17272_, _02877_);
  and (_17274_, _11562_, _04635_);
  or (_17275_, _17274_, _17243_);
  or (_17276_, _17275_, _02987_);
  and (_17277_, _17276_, _06246_);
  and (_17278_, _17277_, _17273_);
  or (_17279_, _17278_, _17248_);
  and (_17280_, _17279_, _02986_);
  or (_17281_, _11613_, _11562_);
  and (_17283_, _17281_, _04635_);
  or (_17284_, _17283_, _17243_);
  and (_17285_, _17284_, _02866_);
  or (_17286_, _17285_, _05535_);
  or (_17287_, _17286_, _17280_);
  or (_17288_, _17264_, _02859_);
  and (_17289_, _17288_, _17287_);
  or (_17290_, _17289_, _02841_);
  and (_17291_, _06162_, _04654_);
  or (_17292_, _17250_, _02842_);
  or (_17294_, _17292_, _17291_);
  and (_17295_, _17294_, _02839_);
  and (_17296_, _17295_, _17290_);
  nor (_17297_, _11671_, _08393_);
  or (_17298_, _17297_, _17250_);
  and (_17299_, _17298_, _02567_);
  or (_17300_, _17299_, _08207_);
  or (_17301_, _17300_, _17296_);
  and (_17302_, _11560_, _04654_);
  or (_17303_, _17250_, _07139_);
  or (_17305_, _17303_, _17302_);
  and (_17306_, _11678_, _04654_);
  or (_17307_, _17306_, _17250_);
  or (_17308_, _17307_, _07140_);
  and (_17309_, _17308_, _07150_);
  and (_17310_, _17309_, _17305_);
  and (_17311_, _17310_, _17301_);
  and (_17312_, _11556_, _04654_);
  or (_17313_, _17312_, _17250_);
  and (_17314_, _17313_, _03148_);
  or (_17316_, _17314_, _17311_);
  and (_17317_, _17316_, _03138_);
  or (_17318_, _17250_, _04838_);
  and (_17319_, _17255_, _03137_);
  and (_17320_, _17307_, _03022_);
  or (_17321_, _17320_, _17319_);
  and (_17322_, _17321_, _17318_);
  or (_17323_, _17322_, _03042_);
  or (_17324_, _17323_, _17317_);
  nor (_17325_, _11558_, _08393_);
  or (_17327_, _17250_, _03043_);
  or (_17328_, _17327_, _17325_);
  and (_17329_, _17328_, _07161_);
  and (_17330_, _17329_, _17324_);
  nor (_17331_, _11555_, _08393_);
  or (_17332_, _17331_, _17250_);
  and (_17333_, _17332_, _03143_);
  or (_17334_, _17333_, _03174_);
  or (_17335_, _17334_, _17330_);
  or (_17336_, _17252_, _03179_);
  and (_17338_, _17336_, _03183_);
  and (_17339_, _17338_, _17335_);
  and (_17340_, _17275_, _02799_);
  or (_17341_, _17340_, _02887_);
  or (_17342_, _17341_, _17339_);
  and (_17343_, _11744_, _04654_);
  or (_17344_, _17250_, _02888_);
  or (_17345_, _17344_, _17343_);
  and (_17346_, _17345_, _34655_);
  and (_17347_, _17346_, _17342_);
  or (_35834_[6], _17347_, _17242_);
  not (_17349_, \oc8051_golden_model_1.P1 [0]);
  nor (_17350_, _34655_, _17349_);
  or (_17351_, _17350_, rst);
  nor (_17352_, _04660_, _17349_);
  and (_17353_, _10369_, _04660_);
  or (_17354_, _17353_, _17352_);
  and (_17355_, _17354_, _03148_);
  and (_17356_, _04660_, _03838_);
  or (_17357_, _17356_, _17352_);
  or (_17359_, _17357_, _02859_);
  nor (_17360_, _05332_, _17349_);
  and (_17361_, _10390_, _05332_);
  or (_17362_, _17361_, _17360_);
  and (_17363_, _17362_, _02884_);
  nor (_17364_, _05085_, _08493_);
  or (_17365_, _17364_, _17352_);
  or (_17366_, _17365_, _03006_);
  and (_17367_, _04660_, \oc8051_golden_model_1.ACC [0]);
  or (_17368_, _17367_, _17352_);
  and (_17370_, _17368_, _03845_);
  nor (_17371_, _03845_, _17349_);
  or (_17372_, _17371_, _02948_);
  or (_17373_, _17372_, _17370_);
  and (_17374_, _17373_, _02976_);
  and (_17375_, _17374_, _17366_);
  and (_17376_, _17357_, _02946_);
  or (_17377_, _17376_, _02880_);
  or (_17378_, _17377_, _17375_);
  or (_17379_, _17378_, _17363_);
  or (_17381_, _17368_, _02992_);
  and (_17382_, _17381_, _02987_);
  and (_17383_, _17382_, _17379_);
  and (_17384_, _17352_, _02877_);
  or (_17385_, _17384_, _02871_);
  or (_17386_, _17385_, _17383_);
  or (_17387_, _17365_, _06246_);
  and (_17388_, _17387_, _02986_);
  and (_17389_, _17388_, _17386_);
  and (_17390_, _16632_, _05332_);
  or (_17392_, _17390_, _17360_);
  and (_17393_, _17392_, _02866_);
  or (_17394_, _17393_, _05535_);
  or (_17395_, _17394_, _17389_);
  and (_17396_, _17395_, _17359_);
  or (_17397_, _17396_, _02841_);
  and (_17398_, _06164_, _04660_);
  or (_17399_, _17352_, _02842_);
  or (_17400_, _17399_, _17398_);
  and (_17401_, _17400_, _02839_);
  and (_17403_, _17401_, _17397_);
  nor (_17404_, _10475_, _08493_);
  or (_17405_, _17404_, _17352_);
  and (_17406_, _17405_, _02567_);
  or (_17407_, _17406_, _08207_);
  or (_17408_, _17407_, _17403_);
  and (_17409_, _10372_, _04660_);
  or (_17410_, _17352_, _07139_);
  or (_17411_, _17410_, _17409_);
  and (_17412_, _04660_, _05660_);
  or (_17414_, _17412_, _17352_);
  or (_17415_, _17414_, _07140_);
  and (_17416_, _17415_, _07150_);
  and (_17417_, _17416_, _17411_);
  and (_17418_, _17417_, _17408_);
  or (_17419_, _17418_, _17355_);
  and (_17420_, _17419_, _03138_);
  nand (_17421_, _17414_, _03022_);
  nor (_17422_, _17421_, _17364_);
  or (_17423_, _17352_, _05085_);
  and (_17425_, _17368_, _03137_);
  and (_17426_, _17425_, _17423_);
  or (_17427_, _17426_, _03042_);
  or (_17428_, _17427_, _17422_);
  or (_17429_, _17428_, _17420_);
  nor (_17430_, _10365_, _08493_);
  or (_17431_, _17352_, _03043_);
  or (_17432_, _17431_, _17430_);
  and (_17433_, _17432_, _07161_);
  and (_17434_, _17433_, _17429_);
  nor (_17436_, _10367_, _08493_);
  or (_17437_, _17436_, _17352_);
  and (_17438_, _17437_, _03143_);
  or (_17439_, _17438_, _03174_);
  or (_17440_, _17439_, _17434_);
  or (_17441_, _17365_, _03179_);
  and (_17442_, _17441_, _03183_);
  and (_17443_, _17442_, _17440_);
  and (_17444_, _17352_, _02799_);
  or (_17445_, _17444_, _02887_);
  or (_17447_, _17445_, _17443_);
  or (_17448_, _17365_, _02888_);
  and (_17449_, _17448_, _34655_);
  and (_17450_, _17449_, _17447_);
  or (_35836_[0], _17450_, _17351_);
  not (_17451_, \oc8051_golden_model_1.P1 [1]);
  nor (_17452_, _34655_, _17451_);
  or (_17453_, _17452_, rst);
  or (_17454_, _10565_, _08493_);
  or (_17455_, _04660_, \oc8051_golden_model_1.P1 [1]);
  and (_17457_, _17455_, _03148_);
  and (_17458_, _17457_, _17454_);
  and (_17459_, _16701_, _05332_);
  nor (_17460_, _05332_, _17451_);
  or (_17461_, _17460_, _02986_);
  or (_17462_, _17461_, _17459_);
  and (_17463_, _10574_, _04660_);
  not (_17464_, _17463_);
  and (_17465_, _17464_, _17455_);
  or (_17466_, _17465_, _03006_);
  nand (_17468_, _04660_, _02543_);
  and (_17469_, _17468_, _17455_);
  and (_17470_, _17469_, _03845_);
  nor (_17471_, _03845_, _17451_);
  or (_17472_, _17471_, _02948_);
  or (_17473_, _17472_, _17470_);
  and (_17474_, _17473_, _02976_);
  and (_17475_, _17474_, _17466_);
  nor (_17476_, _04660_, _17451_);
  nor (_17477_, _08493_, _04020_);
  or (_17479_, _17477_, _17476_);
  and (_17480_, _17479_, _02946_);
  and (_17481_, _10569_, _05332_);
  or (_17482_, _17481_, _17460_);
  and (_17483_, _17482_, _02884_);
  or (_17484_, _17483_, _17480_);
  or (_17485_, _17484_, _02880_);
  or (_17486_, _17485_, _17475_);
  or (_17487_, _17469_, _02992_);
  and (_17488_, _17487_, _17486_);
  or (_17490_, _17488_, _02877_);
  and (_17491_, _10572_, _05332_);
  or (_17492_, _17491_, _17460_);
  or (_17493_, _17492_, _02987_);
  and (_17494_, _17493_, _06246_);
  and (_17495_, _17494_, _17490_);
  and (_17496_, _17481_, _10568_);
  or (_17497_, _17496_, _17460_);
  and (_17498_, _17497_, _02871_);
  or (_17499_, _17498_, _02866_);
  or (_17501_, _17499_, _17495_);
  and (_17502_, _17501_, _17462_);
  or (_17503_, _17502_, _05535_);
  or (_17504_, _17479_, _02859_);
  and (_17505_, _17504_, _17503_);
  or (_17506_, _17505_, _02841_);
  and (_17507_, _06163_, _04660_);
  or (_17508_, _17476_, _02842_);
  or (_17509_, _17508_, _17507_);
  and (_17510_, _17509_, _02839_);
  and (_17512_, _17510_, _17506_);
  and (_17513_, _10674_, _04660_);
  or (_17514_, _17513_, _17476_);
  and (_17515_, _17514_, _02567_);
  or (_17516_, _17515_, _17512_);
  and (_17517_, _17516_, _03052_);
  or (_17518_, _10689_, _08493_);
  and (_17519_, _17518_, _03051_);
  nand (_17520_, _04660_, _03720_);
  and (_17521_, _17520_, _02834_);
  or (_17523_, _17521_, _17519_);
  and (_17524_, _17523_, _17455_);
  or (_17525_, _17524_, _17517_);
  and (_17526_, _17525_, _07150_);
  or (_17527_, _17526_, _17458_);
  and (_17528_, _17527_, _03138_);
  or (_17529_, _10688_, _08493_);
  and (_17530_, _17455_, _03022_);
  and (_17531_, _17530_, _17529_);
  or (_17532_, _17476_, _05038_);
  and (_17534_, _17469_, _03137_);
  and (_17535_, _17534_, _17532_);
  or (_17536_, _17535_, _17531_);
  or (_17537_, _17536_, _17528_);
  and (_17538_, _17537_, _03144_);
  or (_17539_, _17520_, _05038_);
  and (_17540_, _17455_, _03042_);
  and (_17541_, _17540_, _17539_);
  or (_17542_, _17468_, _05038_);
  and (_17543_, _17455_, _03143_);
  and (_17545_, _17543_, _17542_);
  or (_17546_, _17545_, _03174_);
  or (_17547_, _17546_, _17541_);
  or (_17548_, _17547_, _17538_);
  or (_17549_, _17465_, _03179_);
  and (_17550_, _17549_, _03183_);
  and (_17551_, _17550_, _17548_);
  and (_17552_, _17492_, _02799_);
  or (_17553_, _17552_, _02887_);
  or (_17554_, _17553_, _17551_);
  or (_17556_, _17476_, _02888_);
  or (_17557_, _17556_, _17463_);
  and (_17558_, _17557_, _34655_);
  and (_17559_, _17558_, _17554_);
  or (_35836_[1], _17559_, _17453_);
  not (_17560_, \oc8051_golden_model_1.P1 [2]);
  nor (_17561_, _34655_, _17560_);
  or (_17562_, _17561_, rst);
  nor (_17563_, _04660_, _17560_);
  nor (_17564_, _08493_, _04449_);
  or (_17566_, _17564_, _17563_);
  or (_17567_, _17566_, _02859_);
  nor (_17568_, _10788_, _08493_);
  or (_17569_, _17568_, _17563_);
  or (_17570_, _17569_, _03006_);
  and (_17571_, _04660_, \oc8051_golden_model_1.ACC [2]);
  or (_17572_, _17571_, _17563_);
  and (_17573_, _17572_, _03845_);
  nor (_17574_, _03845_, _17560_);
  or (_17575_, _17574_, _02948_);
  or (_17577_, _17575_, _17573_);
  and (_17578_, _17577_, _02976_);
  and (_17579_, _17578_, _17570_);
  and (_17580_, _17566_, _02946_);
  nor (_17581_, _05332_, _17560_);
  and (_17582_, _10792_, _05332_);
  or (_17583_, _17582_, _17581_);
  and (_17584_, _17583_, _02884_);
  or (_17585_, _17584_, _17580_);
  or (_17586_, _17585_, _02880_);
  or (_17588_, _17586_, _17579_);
  or (_17589_, _17572_, _02992_);
  and (_17590_, _17589_, _17588_);
  or (_17591_, _17590_, _02877_);
  and (_17592_, _10773_, _05332_);
  or (_17593_, _17592_, _17581_);
  or (_17594_, _17593_, _02987_);
  and (_17595_, _17594_, _06246_);
  and (_17596_, _17595_, _17591_);
  and (_17597_, _17582_, _10807_);
  or (_17599_, _17597_, _17581_);
  and (_17600_, _17599_, _02871_);
  or (_17601_, _17600_, _17596_);
  and (_17602_, _17601_, _02986_);
  and (_17603_, _16847_, _05332_);
  or (_17604_, _17581_, _17603_);
  and (_17605_, _17604_, _02866_);
  or (_17606_, _17605_, _05535_);
  or (_17607_, _17606_, _17602_);
  and (_17608_, _17607_, _17567_);
  or (_17610_, _17608_, _02841_);
  and (_17611_, _06167_, _04660_);
  or (_17612_, _17563_, _02842_);
  or (_17613_, _17612_, _17611_);
  and (_17614_, _17613_, _02839_);
  and (_17615_, _17614_, _17610_);
  nor (_17616_, _10881_, _08493_);
  or (_17617_, _17616_, _17563_);
  and (_17618_, _17617_, _02567_);
  or (_17619_, _17618_, _17615_);
  or (_17621_, _17619_, _08207_);
  and (_17622_, _10770_, _04660_);
  or (_17623_, _17563_, _07139_);
  or (_17624_, _17623_, _17622_);
  and (_17625_, _04660_, _05693_);
  or (_17626_, _17625_, _17563_);
  or (_17627_, _17626_, _07140_);
  and (_17628_, _17627_, _07150_);
  and (_17629_, _17628_, _17624_);
  and (_17630_, _17629_, _17621_);
  and (_17632_, _10766_, _04660_);
  or (_17633_, _17632_, _17563_);
  and (_17634_, _17633_, _03148_);
  or (_17635_, _17634_, _17630_);
  and (_17636_, _17635_, _03138_);
  or (_17637_, _17563_, _05135_);
  and (_17638_, _17572_, _03137_);
  and (_17639_, _17626_, _03022_);
  or (_17640_, _17639_, _17638_);
  and (_17641_, _17640_, _17637_);
  or (_17643_, _17641_, _03042_);
  or (_17644_, _17643_, _17636_);
  nor (_17645_, _10768_, _08493_);
  or (_17646_, _17563_, _03043_);
  or (_17647_, _17646_, _17645_);
  and (_17648_, _17647_, _07161_);
  and (_17649_, _17648_, _17644_);
  nor (_17650_, _10765_, _08493_);
  or (_17651_, _17650_, _17563_);
  and (_17652_, _17651_, _03143_);
  or (_17654_, _17652_, _03174_);
  or (_17655_, _17654_, _17649_);
  or (_17656_, _17569_, _03179_);
  and (_17657_, _17656_, _03183_);
  and (_17658_, _17657_, _17655_);
  and (_17659_, _17593_, _02799_);
  or (_17660_, _17659_, _02887_);
  or (_17661_, _17660_, _17658_);
  and (_17662_, _10941_, _04660_);
  or (_17663_, _17563_, _02888_);
  or (_17665_, _17663_, _17662_);
  and (_17666_, _17665_, _34655_);
  and (_17667_, _17666_, _17661_);
  or (_35836_[2], _17667_, _17562_);
  nor (_17668_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_17669_, _17668_, _04552_);
  and (_17670_, _08493_, \oc8051_golden_model_1.P1 [3]);
  nor (_17671_, _08493_, _04275_);
  or (_17672_, _17671_, _17670_);
  or (_17673_, _17672_, _02859_);
  and (_17675_, _16920_, _05332_);
  not (_17676_, _05332_);
  and (_17677_, _17676_, \oc8051_golden_model_1.P1 [3]);
  or (_17678_, _17677_, _02986_);
  or (_17679_, _17678_, _17675_);
  nor (_17680_, _10983_, _08493_);
  or (_17681_, _17680_, _17670_);
  or (_17682_, _17681_, _03006_);
  and (_17683_, _04660_, \oc8051_golden_model_1.ACC [3]);
  or (_17684_, _17683_, _17670_);
  and (_17686_, _17684_, _03845_);
  and (_17687_, _04194_, \oc8051_golden_model_1.P1 [3]);
  or (_17688_, _17687_, _02948_);
  or (_17689_, _17688_, _17686_);
  and (_17690_, _17689_, _02976_);
  and (_17691_, _17690_, _17682_);
  and (_17692_, _17672_, _02946_);
  and (_17693_, _10976_, _05332_);
  or (_17694_, _17693_, _17677_);
  and (_17695_, _17694_, _02884_);
  or (_17697_, _17695_, _17692_);
  or (_17698_, _17697_, _02880_);
  or (_17699_, _17698_, _17691_);
  or (_17700_, _17684_, _02992_);
  and (_17701_, _17700_, _17699_);
  or (_17702_, _17701_, _02877_);
  and (_17703_, _10979_, _05332_);
  or (_17704_, _17703_, _17677_);
  or (_17705_, _17704_, _02987_);
  and (_17706_, _17705_, _06246_);
  and (_17708_, _17706_, _17702_);
  or (_17709_, _17677_, _10975_);
  and (_17710_, _17709_, _02871_);
  and (_17711_, _17710_, _17694_);
  or (_17712_, _17711_, _02866_);
  or (_17713_, _17712_, _17708_);
  and (_17714_, _17713_, _17679_);
  or (_17715_, _17714_, _05535_);
  and (_17716_, _17715_, _17673_);
  or (_17717_, _17716_, _02841_);
  and (_17719_, _06166_, _04660_);
  or (_17720_, _17670_, _02842_);
  or (_17721_, _17720_, _17719_);
  and (_17722_, _17721_, _02839_);
  and (_17723_, _17722_, _17717_);
  nor (_17724_, _11076_, _08493_);
  or (_17725_, _17670_, _17724_);
  and (_17726_, _17725_, _02567_);
  or (_17727_, _17726_, _17723_);
  or (_17728_, _17727_, _08207_);
  and (_17730_, _10968_, _04660_);
  or (_17731_, _17670_, _07139_);
  or (_17732_, _17731_, _17730_);
  and (_17733_, _04660_, _05654_);
  or (_17734_, _17733_, _17670_);
  or (_17735_, _17734_, _07140_);
  and (_17736_, _17735_, _07150_);
  and (_17737_, _17736_, _17732_);
  and (_17738_, _17737_, _17728_);
  and (_17739_, _10964_, _04660_);
  or (_17741_, _17739_, _17670_);
  and (_17742_, _17741_, _03148_);
  or (_17743_, _17742_, _17738_);
  and (_17744_, _17743_, _03138_);
  or (_17745_, _17670_, _04993_);
  and (_17746_, _17684_, _03137_);
  and (_17747_, _17734_, _03022_);
  or (_17748_, _17747_, _17746_);
  and (_17749_, _17748_, _17745_);
  or (_17750_, _17749_, _03042_);
  or (_17752_, _17750_, _17744_);
  nor (_17753_, _10967_, _08493_);
  or (_17754_, _17670_, _03043_);
  or (_17755_, _17754_, _17753_);
  and (_17756_, _17755_, _07161_);
  and (_17757_, _17756_, _17752_);
  nor (_17758_, _10962_, _08493_);
  or (_17759_, _17758_, _17670_);
  and (_17760_, _17759_, _03143_);
  or (_17761_, _17760_, _03174_);
  or (_17763_, _17761_, _17757_);
  or (_17764_, _17681_, _03179_);
  and (_17765_, _17764_, _03183_);
  and (_17766_, _17765_, _17763_);
  and (_17767_, _17704_, _02799_);
  or (_17768_, _17767_, _02887_);
  or (_17769_, _17768_, _17766_);
  and (_17770_, _11136_, _04660_);
  or (_17771_, _17670_, _02888_);
  or (_17772_, _17771_, _17770_);
  and (_17774_, _17772_, _34655_);
  and (_17775_, _17774_, _17769_);
  or (_35836_[3], _17775_, _17669_);
  nor (_17776_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_17777_, _17776_, _04552_);
  and (_17778_, _08493_, \oc8051_golden_model_1.P1 [4]);
  nor (_17779_, _05192_, _08493_);
  or (_17780_, _17779_, _17778_);
  or (_17781_, _17780_, _02859_);
  and (_17782_, _17676_, \oc8051_golden_model_1.P1 [4]);
  and (_17784_, _11167_, _05332_);
  or (_17785_, _17784_, _17782_);
  or (_17786_, _17782_, _11201_);
  and (_17787_, _17786_, _02871_);
  and (_17788_, _17787_, _17785_);
  nor (_17789_, _11184_, _08493_);
  or (_17790_, _17789_, _17778_);
  or (_17791_, _17790_, _03006_);
  and (_17792_, _04660_, \oc8051_golden_model_1.ACC [4]);
  or (_17793_, _17792_, _17778_);
  and (_17795_, _17793_, _03845_);
  and (_17796_, _04194_, \oc8051_golden_model_1.P1 [4]);
  or (_17797_, _17796_, _02948_);
  or (_17798_, _17797_, _17795_);
  and (_17799_, _17798_, _02976_);
  and (_17800_, _17799_, _17791_);
  and (_17801_, _17780_, _02946_);
  and (_17802_, _17785_, _02884_);
  or (_17803_, _17802_, _17801_);
  or (_17804_, _17803_, _02880_);
  or (_17806_, _17804_, _17800_);
  or (_17807_, _17793_, _02992_);
  and (_17808_, _17807_, _17806_);
  or (_17809_, _17808_, _02877_);
  and (_17810_, _11165_, _05332_);
  or (_17811_, _17810_, _17782_);
  or (_17812_, _17811_, _02987_);
  and (_17813_, _17812_, _06246_);
  and (_17814_, _17813_, _17809_);
  or (_17815_, _17814_, _17788_);
  and (_17817_, _17815_, _02986_);
  and (_17818_, _17065_, _05332_);
  or (_17819_, _17818_, _17782_);
  and (_17820_, _17819_, _02866_);
  or (_17821_, _17820_, _05535_);
  or (_17822_, _17821_, _17817_);
  and (_17823_, _17822_, _17781_);
  or (_17824_, _17823_, _02841_);
  and (_17825_, _06171_, _04660_);
  or (_17826_, _17778_, _02842_);
  or (_17828_, _17826_, _17825_);
  and (_17829_, _17828_, _02839_);
  and (_17830_, _17829_, _17824_);
  nor (_17831_, _11271_, _08493_);
  or (_17832_, _17831_, _17778_);
  and (_17833_, _17832_, _02567_);
  or (_17834_, _17833_, _17830_);
  or (_17835_, _17834_, _08207_);
  and (_17836_, _11158_, _04660_);
  or (_17837_, _17778_, _07139_);
  or (_17839_, _17837_, _17836_);
  and (_17840_, _05618_, _04660_);
  or (_17841_, _17840_, _17778_);
  or (_17842_, _17841_, _07140_);
  and (_17843_, _17842_, _07150_);
  and (_17844_, _17843_, _17839_);
  and (_17845_, _17844_, _17835_);
  and (_17846_, _11154_, _04660_);
  or (_17847_, _17846_, _17778_);
  and (_17848_, _17847_, _03148_);
  or (_17850_, _17848_, _17845_);
  and (_17851_, _17850_, _03138_);
  or (_17852_, _17778_, _05240_);
  and (_17853_, _17793_, _03137_);
  and (_17854_, _17841_, _03022_);
  or (_17855_, _17854_, _17853_);
  and (_17856_, _17855_, _17852_);
  or (_17857_, _17856_, _03042_);
  or (_17858_, _17857_, _17851_);
  nor (_17859_, _11157_, _08493_);
  or (_17861_, _17778_, _03043_);
  or (_17862_, _17861_, _17859_);
  and (_17863_, _17862_, _07161_);
  and (_17864_, _17863_, _17858_);
  nor (_17865_, _11152_, _08493_);
  or (_17866_, _17865_, _17778_);
  and (_17867_, _17866_, _03143_);
  or (_17868_, _17867_, _03174_);
  or (_17869_, _17868_, _17864_);
  or (_17870_, _17790_, _03179_);
  and (_17872_, _17870_, _03183_);
  and (_17873_, _17872_, _17869_);
  and (_17874_, _17811_, _02799_);
  or (_17875_, _17874_, _02887_);
  or (_17876_, _17875_, _17873_);
  and (_17877_, _11338_, _04660_);
  or (_17878_, _17778_, _02888_);
  or (_17879_, _17878_, _17877_);
  and (_17880_, _17879_, _34655_);
  and (_17881_, _17880_, _17876_);
  or (_35836_[4], _17881_, _17777_);
  nor (_17883_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_17884_, _17883_, _04552_);
  and (_17885_, _08493_, \oc8051_golden_model_1.P1 [5]);
  nor (_17886_, _11380_, _08493_);
  or (_17887_, _17886_, _17885_);
  or (_17888_, _17887_, _03006_);
  and (_17889_, _04660_, \oc8051_golden_model_1.ACC [5]);
  or (_17890_, _17889_, _17885_);
  and (_17891_, _17890_, _03845_);
  and (_17893_, _04194_, \oc8051_golden_model_1.P1 [5]);
  or (_17894_, _17893_, _02948_);
  or (_17895_, _17894_, _17891_);
  and (_17896_, _17895_, _02976_);
  and (_17897_, _17896_, _17888_);
  nor (_17898_, _04894_, _08493_);
  or (_17899_, _17898_, _17885_);
  and (_17900_, _17899_, _02946_);
  and (_17901_, _17676_, \oc8051_golden_model_1.P1 [5]);
  and (_17902_, _11365_, _05332_);
  or (_17904_, _17902_, _17901_);
  and (_17905_, _17904_, _02884_);
  or (_17906_, _17905_, _17900_);
  or (_17907_, _17906_, _02880_);
  or (_17908_, _17907_, _17897_);
  or (_17909_, _17890_, _02992_);
  and (_17910_, _17909_, _17908_);
  or (_17911_, _17910_, _02877_);
  and (_17912_, _11363_, _05332_);
  or (_17913_, _17912_, _17901_);
  or (_17915_, _17913_, _02987_);
  and (_17916_, _17915_, _06246_);
  and (_17917_, _17916_, _17911_);
  and (_17918_, _11398_, _05332_);
  or (_17919_, _17918_, _17901_);
  and (_17920_, _17919_, _02871_);
  or (_17921_, _17920_, _17917_);
  and (_17922_, _17921_, _02986_);
  and (_17923_, _17171_, _05332_);
  or (_17924_, _17923_, _17901_);
  and (_17926_, _17924_, _02866_);
  or (_17927_, _17926_, _05535_);
  or (_17928_, _17927_, _17922_);
  or (_17929_, _17899_, _02859_);
  and (_17930_, _17929_, _17928_);
  or (_17931_, _17930_, _02841_);
  and (_17932_, _06170_, _04660_);
  or (_17933_, _17885_, _02842_);
  or (_17934_, _17933_, _17932_);
  and (_17935_, _17934_, _02839_);
  and (_17937_, _17935_, _17931_);
  nor (_17938_, _11467_, _08493_);
  or (_17939_, _17938_, _17885_);
  and (_17940_, _17939_, _02567_);
  or (_17941_, _17940_, _08207_);
  or (_17942_, _17941_, _17937_);
  and (_17943_, _11482_, _04660_);
  or (_17944_, _17885_, _07139_);
  or (_17945_, _17944_, _17943_);
  and (_17946_, _05671_, _04660_);
  or (_17948_, _17946_, _17885_);
  or (_17949_, _17948_, _07140_);
  and (_17950_, _17949_, _07150_);
  and (_17951_, _17950_, _17945_);
  and (_17952_, _17951_, _17942_);
  and (_17953_, _11356_, _04660_);
  or (_17954_, _17953_, _17885_);
  and (_17955_, _17954_, _03148_);
  or (_17956_, _17955_, _17952_);
  and (_17957_, _17956_, _03138_);
  or (_17959_, _17885_, _04945_);
  and (_17960_, _17890_, _03137_);
  and (_17961_, _17948_, _03022_);
  or (_17962_, _17961_, _17960_);
  and (_17963_, _17962_, _17959_);
  or (_17964_, _17963_, _03042_);
  or (_17965_, _17964_, _17957_);
  nor (_17966_, _11480_, _08493_);
  or (_17967_, _17885_, _03043_);
  or (_17968_, _17967_, _17966_);
  and (_17970_, _17968_, _07161_);
  and (_17971_, _17970_, _17965_);
  nor (_17972_, _11355_, _08493_);
  or (_17973_, _17972_, _17885_);
  and (_17974_, _17973_, _03143_);
  or (_17975_, _17974_, _03174_);
  or (_17976_, _17975_, _17971_);
  or (_17977_, _17887_, _03179_);
  and (_17978_, _17977_, _03183_);
  and (_17979_, _17978_, _17976_);
  and (_17981_, _17913_, _02799_);
  or (_17982_, _17981_, _02887_);
  or (_17983_, _17982_, _17979_);
  and (_17984_, _11541_, _04660_);
  or (_17985_, _17885_, _02888_);
  or (_17986_, _17985_, _17984_);
  and (_17987_, _17986_, _34655_);
  and (_17988_, _17987_, _17983_);
  or (_35836_[5], _17988_, _17884_);
  not (_17989_, \oc8051_golden_model_1.P1 [6]);
  nor (_17991_, _34655_, _17989_);
  or (_17992_, _17991_, rst);
  nor (_17993_, _05332_, _17989_);
  and (_17994_, _11564_, _05332_);
  or (_17995_, _17994_, _17993_);
  or (_17996_, _17993_, _11596_);
  and (_17997_, _17996_, _02871_);
  and (_17998_, _17997_, _17995_);
  nor (_17999_, _04660_, _17989_);
  nor (_18000_, _11567_, _08493_);
  or (_18002_, _18000_, _17999_);
  or (_18003_, _18002_, _03006_);
  and (_18004_, _04660_, \oc8051_golden_model_1.ACC [6]);
  or (_18005_, _18004_, _17999_);
  and (_18006_, _18005_, _03845_);
  nor (_18007_, _03845_, _17989_);
  or (_18008_, _18007_, _02948_);
  or (_18009_, _18008_, _18006_);
  and (_18010_, _18009_, _02976_);
  and (_18011_, _18010_, _18003_);
  nor (_18013_, _04790_, _08493_);
  or (_18014_, _18013_, _17999_);
  and (_18015_, _18014_, _02946_);
  and (_18016_, _17995_, _02884_);
  or (_18017_, _18016_, _18015_);
  or (_18018_, _18017_, _02880_);
  or (_18019_, _18018_, _18011_);
  or (_18020_, _18005_, _02992_);
  and (_18021_, _18020_, _18019_);
  or (_18022_, _18021_, _02877_);
  and (_18024_, _11562_, _05332_);
  or (_18025_, _18024_, _17993_);
  or (_18026_, _18025_, _02987_);
  and (_18027_, _18026_, _06246_);
  and (_18028_, _18027_, _18022_);
  or (_18029_, _18028_, _17998_);
  and (_18030_, _18029_, _02986_);
  and (_18031_, _17281_, _05332_);
  or (_18032_, _18031_, _17993_);
  and (_18033_, _18032_, _02866_);
  or (_18035_, _18033_, _05535_);
  or (_18036_, _18035_, _18030_);
  or (_18037_, _18014_, _02859_);
  and (_18038_, _18037_, _18036_);
  or (_18039_, _18038_, _02841_);
  and (_18040_, _06162_, _04660_);
  or (_18041_, _17999_, _02842_);
  or (_18042_, _18041_, _18040_);
  and (_18043_, _18042_, _02839_);
  and (_18044_, _18043_, _18039_);
  nor (_18046_, _11671_, _08493_);
  or (_18047_, _18046_, _17999_);
  and (_18048_, _18047_, _02567_);
  or (_18049_, _18048_, _08207_);
  or (_18050_, _18049_, _18044_);
  and (_18051_, _11560_, _04660_);
  or (_18052_, _17999_, _07139_);
  or (_18053_, _18052_, _18051_);
  and (_18054_, _11678_, _04660_);
  or (_18055_, _18054_, _17999_);
  or (_18057_, _18055_, _07140_);
  and (_18058_, _18057_, _07150_);
  and (_18059_, _18058_, _18053_);
  and (_18060_, _18059_, _18050_);
  and (_18061_, _11556_, _04660_);
  or (_18062_, _18061_, _17999_);
  and (_18063_, _18062_, _03148_);
  or (_18064_, _18063_, _18060_);
  and (_18065_, _18064_, _03138_);
  or (_18066_, _17999_, _04838_);
  and (_18068_, _18005_, _03137_);
  and (_18069_, _18055_, _03022_);
  or (_18070_, _18069_, _18068_);
  and (_18071_, _18070_, _18066_);
  or (_18072_, _18071_, _03042_);
  or (_18073_, _18072_, _18065_);
  nor (_18074_, _11558_, _08493_);
  or (_18075_, _17999_, _03043_);
  or (_18076_, _18075_, _18074_);
  and (_18077_, _18076_, _07161_);
  and (_18079_, _18077_, _18073_);
  nor (_18080_, _11555_, _08493_);
  or (_18081_, _18080_, _17999_);
  and (_18082_, _18081_, _03143_);
  or (_18083_, _18082_, _03174_);
  or (_18084_, _18083_, _18079_);
  or (_18085_, _18002_, _03179_);
  and (_18086_, _18085_, _03183_);
  and (_18087_, _18086_, _18084_);
  and (_18088_, _18025_, _02799_);
  or (_18090_, _18088_, _02887_);
  or (_18091_, _18090_, _18087_);
  and (_18092_, _11744_, _04660_);
  or (_18093_, _17999_, _02888_);
  or (_18094_, _18093_, _18092_);
  and (_18095_, _18094_, _34655_);
  and (_18096_, _18095_, _18091_);
  or (_35836_[6], _18096_, _17992_);
  not (_18097_, \oc8051_golden_model_1.P2 [0]);
  nor (_18098_, _34655_, _18097_);
  or (_18100_, _18098_, rst);
  nor (_18101_, _04666_, _18097_);
  and (_18102_, _10369_, _04666_);
  or (_18103_, _18102_, _18101_);
  and (_18104_, _18103_, _03148_);
  and (_18105_, _04666_, _03838_);
  or (_18106_, _18105_, _18101_);
  or (_18107_, _18106_, _02859_);
  nor (_18108_, _05335_, _18097_);
  and (_18109_, _10390_, _05335_);
  or (_18111_, _18109_, _18108_);
  and (_18112_, _18111_, _02884_);
  nor (_18113_, _05085_, _08592_);
  or (_18114_, _18113_, _18101_);
  or (_18115_, _18114_, _03006_);
  and (_18116_, _04666_, \oc8051_golden_model_1.ACC [0]);
  or (_18117_, _18116_, _18101_);
  and (_18118_, _18117_, _03845_);
  nor (_18119_, _03845_, _18097_);
  or (_18120_, _18119_, _02948_);
  or (_18122_, _18120_, _18118_);
  and (_18123_, _18122_, _02976_);
  and (_18124_, _18123_, _18115_);
  and (_18125_, _18106_, _02946_);
  or (_18126_, _18125_, _02880_);
  or (_18127_, _18126_, _18124_);
  or (_18128_, _18127_, _18112_);
  or (_18129_, _18117_, _02992_);
  and (_18130_, _18129_, _02987_);
  and (_18131_, _18130_, _18128_);
  and (_18133_, _18101_, _02877_);
  or (_18134_, _18133_, _02871_);
  or (_18135_, _18134_, _18131_);
  or (_18136_, _18114_, _06246_);
  and (_18137_, _18136_, _02986_);
  and (_18138_, _18137_, _18135_);
  and (_18139_, _16632_, _05335_);
  or (_18140_, _18139_, _18108_);
  and (_18141_, _18140_, _02866_);
  or (_18142_, _18141_, _05535_);
  or (_18144_, _18142_, _18138_);
  and (_18145_, _18144_, _18107_);
  or (_18146_, _18145_, _02841_);
  and (_18147_, _06164_, _04666_);
  or (_18148_, _18101_, _02842_);
  or (_18149_, _18148_, _18147_);
  and (_18150_, _18149_, _02839_);
  and (_18151_, _18150_, _18146_);
  nor (_18152_, _10475_, _08592_);
  or (_18153_, _18152_, _18101_);
  and (_18155_, _18153_, _02567_);
  or (_18156_, _18155_, _08207_);
  or (_18157_, _18156_, _18151_);
  and (_18158_, _10372_, _04666_);
  or (_18159_, _18101_, _07139_);
  or (_18160_, _18159_, _18158_);
  and (_18161_, _04666_, _05660_);
  or (_18162_, _18161_, _18101_);
  or (_18163_, _18162_, _07140_);
  and (_18164_, _18163_, _07150_);
  and (_18166_, _18164_, _18160_);
  and (_18167_, _18166_, _18157_);
  or (_18168_, _18167_, _18104_);
  and (_18169_, _18168_, _03138_);
  nand (_18170_, _18162_, _03022_);
  nor (_18171_, _18170_, _18113_);
  or (_18172_, _18101_, _05085_);
  and (_18173_, _18117_, _03137_);
  and (_18174_, _18173_, _18172_);
  or (_18175_, _18174_, _03042_);
  or (_18177_, _18175_, _18171_);
  or (_18178_, _18177_, _18169_);
  nor (_18179_, _10365_, _08592_);
  or (_18180_, _18101_, _03043_);
  or (_18181_, _18180_, _18179_);
  and (_18182_, _18181_, _07161_);
  and (_18183_, _18182_, _18178_);
  nor (_18184_, _10367_, _08592_);
  or (_18185_, _18184_, _18101_);
  and (_18186_, _18185_, _03143_);
  or (_18188_, _18186_, _03174_);
  or (_18189_, _18188_, _18183_);
  or (_18190_, _18114_, _03179_);
  and (_18191_, _18190_, _03183_);
  and (_18192_, _18191_, _18189_);
  and (_18193_, _18101_, _02799_);
  or (_18194_, _18193_, _02887_);
  or (_18195_, _18194_, _18192_);
  or (_18196_, _18114_, _02888_);
  and (_18197_, _18196_, _34655_);
  and (_18199_, _18197_, _18195_);
  or (_35838_[0], _18199_, _18100_);
  not (_18200_, \oc8051_golden_model_1.P2 [1]);
  nor (_18201_, _34655_, _18200_);
  or (_18202_, _18201_, rst);
  and (_18203_, _16701_, _05335_);
  nor (_18204_, _05335_, _18200_);
  or (_18205_, _18204_, _02986_);
  or (_18206_, _18205_, _18203_);
  or (_18207_, _04666_, \oc8051_golden_model_1.P2 [1]);
  and (_18209_, _10574_, _04666_);
  not (_18210_, _18209_);
  and (_18211_, _18210_, _18207_);
  or (_18212_, _18211_, _03006_);
  nand (_18213_, _04666_, _02543_);
  and (_18214_, _18213_, _18207_);
  and (_18215_, _18214_, _03845_);
  nor (_18216_, _03845_, _18200_);
  or (_18217_, _18216_, _02948_);
  or (_18218_, _18217_, _18215_);
  and (_18220_, _18218_, _02976_);
  and (_18221_, _18220_, _18212_);
  nor (_18222_, _04666_, _18200_);
  nor (_18223_, _08592_, _04020_);
  or (_18224_, _18223_, _18222_);
  and (_18225_, _18224_, _02946_);
  and (_18226_, _10569_, _05335_);
  or (_18227_, _18226_, _18204_);
  and (_18228_, _18227_, _02884_);
  or (_18229_, _18228_, _18225_);
  or (_18231_, _18229_, _02880_);
  or (_18232_, _18231_, _18221_);
  or (_18233_, _18214_, _02992_);
  and (_18234_, _18233_, _18232_);
  or (_18235_, _18234_, _02877_);
  and (_18236_, _10572_, _05335_);
  or (_18237_, _18236_, _18204_);
  or (_18238_, _18237_, _02987_);
  and (_18239_, _18238_, _06246_);
  and (_18240_, _18239_, _18235_);
  and (_18242_, _18226_, _10568_);
  or (_18243_, _18242_, _18204_);
  and (_18244_, _18243_, _02871_);
  or (_18245_, _18244_, _02866_);
  or (_18246_, _18245_, _18240_);
  and (_18247_, _18246_, _18206_);
  or (_18248_, _18247_, _05535_);
  or (_18249_, _18224_, _02859_);
  and (_18250_, _18249_, _18248_);
  or (_18251_, _18250_, _02841_);
  and (_18253_, _06163_, _04666_);
  or (_18254_, _18222_, _02842_);
  or (_18255_, _18254_, _18253_);
  and (_18256_, _18255_, _02839_);
  and (_18257_, _18256_, _18251_);
  and (_18258_, _10674_, _04666_);
  or (_18259_, _18258_, _18222_);
  and (_18260_, _18259_, _02567_);
  or (_18261_, _18260_, _18257_);
  and (_18262_, _18261_, _03052_);
  or (_18264_, _10689_, _08592_);
  and (_18265_, _18264_, _03051_);
  nand (_18266_, _04666_, _03720_);
  and (_18267_, _18266_, _02834_);
  or (_18268_, _18267_, _18265_);
  and (_18269_, _18268_, _18207_);
  or (_18270_, _18269_, _18262_);
  and (_18271_, _18270_, _07150_);
  or (_18272_, _10565_, _08592_);
  and (_18273_, _18207_, _03148_);
  and (_18275_, _18273_, _18272_);
  or (_18276_, _18275_, _18271_);
  and (_18277_, _18276_, _03138_);
  or (_18278_, _18222_, _05038_);
  and (_18279_, _18214_, _03137_);
  and (_18280_, _18279_, _18278_);
  or (_18281_, _10688_, _08592_);
  and (_18282_, _18207_, _03022_);
  and (_18283_, _18282_, _18281_);
  or (_18284_, _18283_, _18280_);
  or (_18286_, _18284_, _18277_);
  and (_18287_, _18286_, _03144_);
  or (_18288_, _18266_, _05038_);
  and (_18289_, _18207_, _03042_);
  and (_18290_, _18289_, _18288_);
  or (_18291_, _18213_, _05038_);
  and (_18292_, _18207_, _03143_);
  and (_18293_, _18292_, _18291_);
  or (_18294_, _18293_, _03174_);
  or (_18295_, _18294_, _18290_);
  or (_18297_, _18295_, _18287_);
  or (_18298_, _18211_, _03179_);
  and (_18299_, _18298_, _03183_);
  and (_18300_, _18299_, _18297_);
  and (_18301_, _18237_, _02799_);
  or (_18302_, _18301_, _02887_);
  or (_18303_, _18302_, _18300_);
  or (_18304_, _18222_, _02888_);
  or (_18305_, _18304_, _18209_);
  and (_18306_, _18305_, _34655_);
  and (_18308_, _18306_, _18303_);
  or (_35838_[1], _18308_, _18202_);
  not (_18309_, \oc8051_golden_model_1.P2 [2]);
  nor (_18310_, _34655_, _18309_);
  or (_18311_, _18310_, rst);
  nor (_18312_, _04666_, _18309_);
  nor (_18313_, _08592_, _04449_);
  or (_18314_, _18313_, _18312_);
  or (_18315_, _18314_, _02859_);
  nor (_18316_, _10788_, _08592_);
  or (_18318_, _18316_, _18312_);
  or (_18319_, _18318_, _03006_);
  and (_18320_, _04666_, \oc8051_golden_model_1.ACC [2]);
  or (_18321_, _18320_, _18312_);
  and (_18322_, _18321_, _03845_);
  nor (_18323_, _03845_, _18309_);
  or (_18324_, _18323_, _02948_);
  or (_18325_, _18324_, _18322_);
  and (_18326_, _18325_, _02976_);
  and (_18327_, _18326_, _18319_);
  and (_18329_, _18314_, _02946_);
  nor (_18330_, _05335_, _18309_);
  and (_18331_, _10792_, _05335_);
  or (_18332_, _18331_, _18330_);
  and (_18333_, _18332_, _02884_);
  or (_18334_, _18333_, _18329_);
  or (_18335_, _18334_, _02880_);
  or (_18336_, _18335_, _18327_);
  or (_18337_, _18321_, _02992_);
  and (_18338_, _18337_, _18336_);
  or (_18340_, _18338_, _02877_);
  and (_18341_, _10773_, _05335_);
  or (_18342_, _18341_, _18330_);
  or (_18343_, _18342_, _02987_);
  and (_18344_, _18343_, _06246_);
  and (_18345_, _18344_, _18340_);
  and (_18346_, _18331_, _10807_);
  or (_18347_, _18346_, _18330_);
  and (_18348_, _18347_, _02871_);
  or (_18349_, _18348_, _18345_);
  and (_18351_, _18349_, _02986_);
  and (_18352_, _16847_, _05335_);
  or (_18353_, _18330_, _18352_);
  and (_18354_, _18353_, _02866_);
  or (_18355_, _18354_, _05535_);
  or (_18356_, _18355_, _18351_);
  and (_18357_, _18356_, _18315_);
  or (_18358_, _18357_, _02841_);
  and (_18359_, _06167_, _04666_);
  or (_18360_, _18312_, _02842_);
  or (_18362_, _18360_, _18359_);
  and (_18363_, _18362_, _02839_);
  and (_18364_, _18363_, _18358_);
  nor (_18365_, _10881_, _08592_);
  or (_18366_, _18365_, _18312_);
  and (_18367_, _18366_, _02567_);
  or (_18368_, _18367_, _18364_);
  or (_18369_, _18368_, _08207_);
  and (_18370_, _10770_, _04666_);
  or (_18371_, _18312_, _07139_);
  or (_18373_, _18371_, _18370_);
  and (_18374_, _04666_, _05693_);
  or (_18375_, _18374_, _18312_);
  or (_18376_, _18375_, _07140_);
  and (_18377_, _18376_, _07150_);
  and (_18378_, _18377_, _18373_);
  and (_18379_, _18378_, _18369_);
  and (_18380_, _10766_, _04666_);
  or (_18381_, _18380_, _18312_);
  and (_18382_, _18381_, _03148_);
  or (_18384_, _18382_, _18379_);
  and (_18385_, _18384_, _03138_);
  or (_18386_, _18312_, _05135_);
  and (_18387_, _18321_, _03137_);
  and (_18388_, _18375_, _03022_);
  or (_18389_, _18388_, _18387_);
  and (_18390_, _18389_, _18386_);
  or (_18391_, _18390_, _03042_);
  or (_18392_, _18391_, _18385_);
  nor (_18393_, _10768_, _08592_);
  or (_18395_, _18312_, _03043_);
  or (_18396_, _18395_, _18393_);
  and (_18397_, _18396_, _07161_);
  and (_18398_, _18397_, _18392_);
  nor (_18399_, _10765_, _08592_);
  or (_18400_, _18399_, _18312_);
  and (_18401_, _18400_, _03143_);
  or (_18402_, _18401_, _03174_);
  or (_18403_, _18402_, _18398_);
  or (_18404_, _18318_, _03179_);
  and (_18406_, _18404_, _03183_);
  and (_18407_, _18406_, _18403_);
  and (_18408_, _18342_, _02799_);
  or (_18409_, _18408_, _02887_);
  or (_18410_, _18409_, _18407_);
  and (_18411_, _10941_, _04666_);
  or (_18412_, _18312_, _02888_);
  or (_18413_, _18412_, _18411_);
  and (_18414_, _18413_, _34655_);
  and (_18415_, _18414_, _18410_);
  or (_35838_[2], _18415_, _18311_);
  nor (_18417_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_18418_, _18417_, _04552_);
  and (_18419_, _08592_, \oc8051_golden_model_1.P2 [3]);
  nor (_18420_, _08592_, _04275_);
  or (_18421_, _18420_, _18419_);
  or (_18422_, _18421_, _02859_);
  and (_18423_, _16920_, _05335_);
  not (_18424_, _05335_);
  and (_18425_, _18424_, \oc8051_golden_model_1.P2 [3]);
  or (_18427_, _18425_, _02986_);
  or (_18428_, _18427_, _18423_);
  nor (_18429_, _10983_, _08592_);
  or (_18430_, _18429_, _18419_);
  or (_18431_, _18430_, _03006_);
  and (_18432_, _04666_, \oc8051_golden_model_1.ACC [3]);
  or (_18433_, _18432_, _18419_);
  and (_18434_, _18433_, _03845_);
  and (_18435_, _04194_, \oc8051_golden_model_1.P2 [3]);
  or (_18436_, _18435_, _02948_);
  or (_18438_, _18436_, _18434_);
  and (_18439_, _18438_, _02976_);
  and (_18440_, _18439_, _18431_);
  and (_18441_, _18421_, _02946_);
  and (_18442_, _10976_, _05335_);
  or (_18443_, _18442_, _18425_);
  and (_18444_, _18443_, _02884_);
  or (_18445_, _18444_, _18441_);
  or (_18446_, _18445_, _02880_);
  or (_18447_, _18446_, _18440_);
  or (_18449_, _18433_, _02992_);
  and (_18450_, _18449_, _18447_);
  or (_18451_, _18450_, _02877_);
  and (_18452_, _10979_, _05335_);
  or (_18453_, _18452_, _18425_);
  or (_18454_, _18453_, _02987_);
  and (_18455_, _18454_, _06246_);
  and (_18456_, _18455_, _18451_);
  or (_18457_, _18425_, _10975_);
  and (_18458_, _18457_, _02871_);
  and (_18460_, _18458_, _18443_);
  or (_18461_, _18460_, _02866_);
  or (_18462_, _18461_, _18456_);
  and (_18463_, _18462_, _18428_);
  or (_18464_, _18463_, _05535_);
  and (_18465_, _18464_, _18422_);
  or (_18466_, _18465_, _02841_);
  and (_18467_, _06166_, _04666_);
  or (_18468_, _18419_, _02842_);
  or (_18469_, _18468_, _18467_);
  and (_18471_, _18469_, _02839_);
  and (_18472_, _18471_, _18466_);
  nor (_18473_, _11076_, _08592_);
  or (_18474_, _18419_, _18473_);
  and (_18475_, _18474_, _02567_);
  or (_18476_, _18475_, _18472_);
  or (_18477_, _18476_, _08207_);
  and (_18478_, _10968_, _04666_);
  or (_18479_, _18419_, _07139_);
  or (_18480_, _18479_, _18478_);
  and (_18482_, _04666_, _05654_);
  or (_18483_, _18482_, _18419_);
  or (_18484_, _18483_, _07140_);
  and (_18485_, _18484_, _07150_);
  and (_18486_, _18485_, _18480_);
  and (_18487_, _18486_, _18477_);
  and (_18488_, _10964_, _04666_);
  or (_18489_, _18488_, _18419_);
  and (_18490_, _18489_, _03148_);
  or (_18491_, _18490_, _18487_);
  and (_18493_, _18491_, _03138_);
  or (_18494_, _18419_, _04993_);
  and (_18495_, _18433_, _03137_);
  and (_18496_, _18483_, _03022_);
  or (_18497_, _18496_, _18495_);
  and (_18498_, _18497_, _18494_);
  or (_18499_, _18498_, _03042_);
  or (_18500_, _18499_, _18493_);
  nor (_18501_, _10967_, _08592_);
  or (_18502_, _18419_, _03043_);
  or (_18504_, _18502_, _18501_);
  and (_18505_, _18504_, _07161_);
  and (_18506_, _18505_, _18500_);
  nor (_18507_, _10962_, _08592_);
  or (_18508_, _18507_, _18419_);
  and (_18509_, _18508_, _03143_);
  or (_18510_, _18509_, _03174_);
  or (_18511_, _18510_, _18506_);
  or (_18512_, _18430_, _03179_);
  and (_18513_, _18512_, _03183_);
  and (_18515_, _18513_, _18511_);
  and (_18516_, _18453_, _02799_);
  or (_18517_, _18516_, _02887_);
  or (_18518_, _18517_, _18515_);
  and (_18519_, _11136_, _04666_);
  or (_18520_, _18419_, _02888_);
  or (_18521_, _18520_, _18519_);
  and (_18522_, _18521_, _34655_);
  and (_18523_, _18522_, _18518_);
  or (_35838_[3], _18523_, _18418_);
  nor (_18525_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_18526_, _18525_, _04552_);
  and (_18527_, _08592_, \oc8051_golden_model_1.P2 [4]);
  nor (_18528_, _05192_, _08592_);
  or (_18529_, _18528_, _18527_);
  or (_18530_, _18529_, _02859_);
  nor (_18531_, _11184_, _08592_);
  or (_18532_, _18531_, _18527_);
  or (_18533_, _18532_, _03006_);
  and (_18534_, _04666_, \oc8051_golden_model_1.ACC [4]);
  or (_18536_, _18534_, _18527_);
  and (_18537_, _18536_, _03845_);
  and (_18538_, _04194_, \oc8051_golden_model_1.P2 [4]);
  or (_18539_, _18538_, _02948_);
  or (_18540_, _18539_, _18537_);
  and (_18541_, _18540_, _02976_);
  and (_18542_, _18541_, _18533_);
  and (_18543_, _18529_, _02946_);
  and (_18544_, _18424_, \oc8051_golden_model_1.P2 [4]);
  and (_18545_, _11167_, _05335_);
  or (_18547_, _18545_, _18544_);
  and (_18548_, _18547_, _02884_);
  or (_18549_, _18548_, _18543_);
  or (_18550_, _18549_, _02880_);
  or (_18551_, _18550_, _18542_);
  or (_18552_, _18536_, _02992_);
  and (_18553_, _18552_, _18551_);
  or (_18554_, _18553_, _02877_);
  and (_18555_, _11165_, _05335_);
  or (_18556_, _18555_, _18544_);
  or (_18558_, _18556_, _02987_);
  and (_18559_, _18558_, _06246_);
  and (_18560_, _18559_, _18554_);
  and (_18561_, _11202_, _05335_);
  or (_18562_, _18561_, _18544_);
  and (_18563_, _18562_, _02871_);
  or (_18564_, _18563_, _18560_);
  and (_18565_, _18564_, _02986_);
  and (_18566_, _17065_, _05335_);
  or (_18567_, _18566_, _18544_);
  and (_18569_, _18567_, _02866_);
  or (_18570_, _18569_, _05535_);
  or (_18571_, _18570_, _18565_);
  and (_18572_, _18571_, _18530_);
  or (_18573_, _18572_, _02841_);
  and (_18574_, _06171_, _04666_);
  or (_18575_, _18527_, _02842_);
  or (_18576_, _18575_, _18574_);
  and (_18577_, _18576_, _02839_);
  and (_18578_, _18577_, _18573_);
  nor (_18580_, _11271_, _08592_);
  or (_18581_, _18580_, _18527_);
  and (_18582_, _18581_, _02567_);
  or (_18583_, _18582_, _18578_);
  or (_18584_, _18583_, _08207_);
  and (_18585_, _11158_, _04666_);
  or (_18586_, _18527_, _07139_);
  or (_18587_, _18586_, _18585_);
  and (_18588_, _05618_, _04666_);
  or (_18589_, _18588_, _18527_);
  or (_18591_, _18589_, _07140_);
  and (_18592_, _18591_, _07150_);
  and (_18593_, _18592_, _18587_);
  and (_18594_, _18593_, _18584_);
  and (_18595_, _11154_, _04666_);
  or (_18596_, _18595_, _18527_);
  and (_18597_, _18596_, _03148_);
  or (_18598_, _18597_, _18594_);
  and (_18599_, _18598_, _03138_);
  or (_18600_, _18527_, _05240_);
  and (_18602_, _18536_, _03137_);
  and (_18603_, _18589_, _03022_);
  or (_18604_, _18603_, _18602_);
  and (_18605_, _18604_, _18600_);
  or (_18606_, _18605_, _03042_);
  or (_18607_, _18606_, _18599_);
  nor (_18608_, _11157_, _08592_);
  or (_18609_, _18527_, _03043_);
  or (_18610_, _18609_, _18608_);
  and (_18611_, _18610_, _07161_);
  and (_18613_, _18611_, _18607_);
  nor (_18614_, _11152_, _08592_);
  or (_18615_, _18614_, _18527_);
  and (_18616_, _18615_, _03143_);
  or (_18617_, _18616_, _03174_);
  or (_18618_, _18617_, _18613_);
  or (_18619_, _18532_, _03179_);
  and (_18620_, _18619_, _03183_);
  and (_18621_, _18620_, _18618_);
  and (_18622_, _18556_, _02799_);
  or (_18624_, _18622_, _02887_);
  or (_18625_, _18624_, _18621_);
  and (_18626_, _11338_, _04666_);
  or (_18627_, _18527_, _02888_);
  or (_18628_, _18627_, _18626_);
  and (_18629_, _18628_, _34655_);
  and (_18630_, _18629_, _18625_);
  or (_35838_[4], _18630_, _18526_);
  nor (_18631_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_18632_, _18631_, _04552_);
  and (_18634_, _18424_, \oc8051_golden_model_1.P2 [5]);
  and (_18635_, _11365_, _05335_);
  or (_18636_, _18635_, _18634_);
  or (_18637_, _18634_, _11397_);
  and (_18638_, _18637_, _02871_);
  and (_18639_, _18638_, _18636_);
  and (_18640_, _08592_, \oc8051_golden_model_1.P2 [5]);
  nor (_18641_, _11380_, _08592_);
  or (_18642_, _18641_, _18640_);
  or (_18643_, _18642_, _03006_);
  and (_18645_, _04666_, \oc8051_golden_model_1.ACC [5]);
  or (_18646_, _18645_, _18640_);
  and (_18647_, _18646_, _03845_);
  and (_18648_, _04194_, \oc8051_golden_model_1.P2 [5]);
  or (_18649_, _18648_, _02948_);
  or (_18650_, _18649_, _18647_);
  and (_18651_, _18650_, _02976_);
  and (_18652_, _18651_, _18643_);
  nor (_18653_, _04894_, _08592_);
  or (_18654_, _18653_, _18640_);
  and (_18656_, _18654_, _02946_);
  and (_18657_, _18636_, _02884_);
  or (_18658_, _18657_, _18656_);
  or (_18659_, _18658_, _02880_);
  or (_18660_, _18659_, _18652_);
  or (_18661_, _18646_, _02992_);
  and (_18662_, _18661_, _18660_);
  or (_18663_, _18662_, _02877_);
  and (_18664_, _11363_, _05335_);
  or (_18665_, _18664_, _18634_);
  or (_18667_, _18665_, _02987_);
  and (_18668_, _18667_, _06246_);
  and (_18669_, _18668_, _18663_);
  or (_18670_, _18669_, _18639_);
  and (_18671_, _18670_, _02986_);
  and (_18672_, _17171_, _05335_);
  or (_18673_, _18672_, _18634_);
  and (_18674_, _18673_, _02866_);
  or (_18675_, _18674_, _05535_);
  or (_18676_, _18675_, _18671_);
  or (_18678_, _18654_, _02859_);
  and (_18679_, _18678_, _18676_);
  or (_18680_, _18679_, _02841_);
  and (_18681_, _06170_, _04666_);
  or (_18682_, _18640_, _02842_);
  or (_18683_, _18682_, _18681_);
  and (_18684_, _18683_, _02839_);
  and (_18685_, _18684_, _18680_);
  nor (_18686_, _11467_, _08592_);
  or (_18687_, _18686_, _18640_);
  and (_18689_, _18687_, _02567_);
  or (_18690_, _18689_, _08207_);
  or (_18691_, _18690_, _18685_);
  and (_18692_, _11482_, _04666_);
  or (_18693_, _18640_, _07139_);
  or (_18694_, _18693_, _18692_);
  and (_18695_, _05671_, _04666_);
  or (_18696_, _18695_, _18640_);
  or (_18697_, _18696_, _07140_);
  and (_18698_, _18697_, _07150_);
  and (_18700_, _18698_, _18694_);
  and (_18701_, _18700_, _18691_);
  and (_18702_, _11356_, _04666_);
  or (_18703_, _18702_, _18640_);
  and (_18704_, _18703_, _03148_);
  or (_18705_, _18704_, _18701_);
  and (_18706_, _18705_, _03138_);
  or (_18707_, _18640_, _04945_);
  and (_18708_, _18646_, _03137_);
  and (_18709_, _18696_, _03022_);
  or (_18711_, _18709_, _18708_);
  and (_18712_, _18711_, _18707_);
  or (_18713_, _18712_, _03042_);
  or (_18714_, _18713_, _18706_);
  nor (_18715_, _11480_, _08592_);
  or (_18716_, _18640_, _03043_);
  or (_18717_, _18716_, _18715_);
  and (_18718_, _18717_, _07161_);
  and (_18719_, _18718_, _18714_);
  nor (_18720_, _11355_, _08592_);
  or (_18722_, _18720_, _18640_);
  and (_18723_, _18722_, _03143_);
  or (_18724_, _18723_, _03174_);
  or (_18725_, _18724_, _18719_);
  or (_18726_, _18642_, _03179_);
  and (_18727_, _18726_, _03183_);
  and (_18728_, _18727_, _18725_);
  and (_18729_, _18665_, _02799_);
  or (_18730_, _18729_, _02887_);
  or (_18731_, _18730_, _18728_);
  and (_18733_, _11541_, _04666_);
  or (_18734_, _18640_, _02888_);
  or (_18735_, _18734_, _18733_);
  and (_18736_, _18735_, _34655_);
  and (_18737_, _18736_, _18731_);
  or (_35838_[5], _18737_, _18632_);
  not (_18738_, \oc8051_golden_model_1.P2 [6]);
  nor (_18739_, _34655_, _18738_);
  or (_18740_, _18739_, rst);
  nor (_18741_, _05335_, _18738_);
  and (_18743_, _11564_, _05335_);
  or (_18744_, _18743_, _18741_);
  or (_18745_, _18741_, _11596_);
  and (_18746_, _18745_, _02871_);
  and (_18747_, _18746_, _18744_);
  nor (_18748_, _04666_, _18738_);
  nor (_18749_, _11567_, _08592_);
  or (_18750_, _18749_, _18748_);
  or (_18751_, _18750_, _03006_);
  and (_18752_, _04666_, \oc8051_golden_model_1.ACC [6]);
  or (_18754_, _18752_, _18748_);
  and (_18755_, _18754_, _03845_);
  nor (_18756_, _03845_, _18738_);
  or (_18757_, _18756_, _02948_);
  or (_18758_, _18757_, _18755_);
  and (_18759_, _18758_, _02976_);
  and (_18760_, _18759_, _18751_);
  nor (_18761_, _04790_, _08592_);
  or (_18762_, _18761_, _18748_);
  and (_18763_, _18762_, _02946_);
  and (_18765_, _18744_, _02884_);
  or (_18766_, _18765_, _18763_);
  or (_18767_, _18766_, _02880_);
  or (_18768_, _18767_, _18760_);
  or (_18769_, _18754_, _02992_);
  and (_18770_, _18769_, _18768_);
  or (_18771_, _18770_, _02877_);
  and (_18772_, _11562_, _05335_);
  or (_18773_, _18772_, _18741_);
  or (_18774_, _18773_, _02987_);
  and (_18776_, _18774_, _06246_);
  and (_18777_, _18776_, _18771_);
  or (_18778_, _18777_, _18747_);
  and (_18779_, _18778_, _02986_);
  and (_18780_, _17281_, _05335_);
  or (_18781_, _18780_, _18741_);
  and (_18782_, _18781_, _02866_);
  or (_18783_, _18782_, _05535_);
  or (_18784_, _18783_, _18779_);
  or (_18785_, _18762_, _02859_);
  and (_18787_, _18785_, _18784_);
  or (_18788_, _18787_, _02841_);
  and (_18789_, _06162_, _04666_);
  or (_18790_, _18748_, _02842_);
  or (_18791_, _18790_, _18789_);
  and (_18792_, _18791_, _02839_);
  and (_18793_, _18792_, _18788_);
  nor (_18794_, _11671_, _08592_);
  or (_18795_, _18794_, _18748_);
  and (_18796_, _18795_, _02567_);
  or (_18798_, _18796_, _08207_);
  or (_18799_, _18798_, _18793_);
  and (_18800_, _11560_, _04666_);
  or (_18801_, _18748_, _07139_);
  or (_18802_, _18801_, _18800_);
  and (_18803_, _11678_, _04666_);
  or (_18804_, _18803_, _18748_);
  or (_18805_, _18804_, _07140_);
  and (_18806_, _18805_, _07150_);
  and (_18807_, _18806_, _18802_);
  and (_18809_, _18807_, _18799_);
  and (_18810_, _11556_, _04666_);
  or (_18811_, _18810_, _18748_);
  and (_18812_, _18811_, _03148_);
  or (_18813_, _18812_, _18809_);
  and (_18814_, _18813_, _03138_);
  or (_18815_, _18748_, _04838_);
  and (_18816_, _18754_, _03137_);
  and (_18817_, _18804_, _03022_);
  or (_18818_, _18817_, _18816_);
  and (_18820_, _18818_, _18815_);
  or (_18821_, _18820_, _03042_);
  or (_18822_, _18821_, _18814_);
  nor (_18823_, _11558_, _08592_);
  or (_18824_, _18748_, _03043_);
  or (_18825_, _18824_, _18823_);
  and (_18826_, _18825_, _07161_);
  and (_18827_, _18826_, _18822_);
  nor (_18828_, _11555_, _08592_);
  or (_18829_, _18828_, _18748_);
  and (_18831_, _18829_, _03143_);
  or (_18832_, _18831_, _03174_);
  or (_18833_, _18832_, _18827_);
  or (_18834_, _18750_, _03179_);
  and (_18835_, _18834_, _03183_);
  and (_18836_, _18835_, _18833_);
  and (_18837_, _18773_, _02799_);
  or (_18838_, _18837_, _02887_);
  or (_18839_, _18838_, _18836_);
  and (_18840_, _11744_, _04666_);
  or (_18842_, _18748_, _02888_);
  or (_18843_, _18842_, _18840_);
  and (_18844_, _18843_, _34655_);
  and (_18845_, _18844_, _18839_);
  or (_35838_[6], _18845_, _18740_);
  not (_18846_, \oc8051_golden_model_1.P3 [0]);
  nor (_18847_, _34655_, _18846_);
  or (_18848_, _18847_, rst);
  nor (_18849_, _04670_, _18846_);
  and (_18850_, _10369_, _04670_);
  or (_18852_, _18850_, _18849_);
  and (_18853_, _18852_, _03148_);
  and (_18854_, _04670_, _03838_);
  or (_18855_, _18854_, _18849_);
  or (_18856_, _18855_, _02859_);
  nor (_18857_, _05337_, _18846_);
  and (_18858_, _10390_, _05337_);
  or (_18859_, _18858_, _18857_);
  and (_18860_, _18859_, _02884_);
  nor (_18861_, _05085_, _08691_);
  or (_18863_, _18861_, _18849_);
  or (_18864_, _18863_, _03006_);
  and (_18865_, _04670_, \oc8051_golden_model_1.ACC [0]);
  or (_18866_, _18865_, _18849_);
  and (_18867_, _18866_, _03845_);
  nor (_18868_, _03845_, _18846_);
  or (_18869_, _18868_, _02948_);
  or (_18870_, _18869_, _18867_);
  and (_18871_, _18870_, _02976_);
  and (_18872_, _18871_, _18864_);
  and (_18874_, _18855_, _02946_);
  or (_18875_, _18874_, _02880_);
  or (_18876_, _18875_, _18872_);
  or (_18877_, _18876_, _18860_);
  or (_18878_, _18866_, _02992_);
  and (_18879_, _18878_, _02987_);
  and (_18880_, _18879_, _18877_);
  and (_18881_, _18849_, _02877_);
  or (_18882_, _18881_, _02871_);
  or (_18883_, _18882_, _18880_);
  or (_18885_, _18863_, _06246_);
  and (_18886_, _18885_, _02986_);
  and (_18887_, _18886_, _18883_);
  and (_18888_, _16632_, _05337_);
  or (_18889_, _18888_, _18857_);
  and (_18890_, _18889_, _02866_);
  or (_18891_, _18890_, _05535_);
  or (_18892_, _18891_, _18887_);
  and (_18893_, _18892_, _18856_);
  or (_18894_, _18893_, _02841_);
  and (_18896_, _06164_, _04670_);
  or (_18897_, _18849_, _02842_);
  or (_18898_, _18897_, _18896_);
  and (_18899_, _18898_, _02839_);
  and (_18900_, _18899_, _18894_);
  nor (_18901_, _10475_, _08691_);
  or (_18902_, _18901_, _18849_);
  and (_18903_, _18902_, _02567_);
  or (_18904_, _18903_, _08207_);
  or (_18905_, _18904_, _18900_);
  and (_18907_, _10372_, _04670_);
  or (_18908_, _18849_, _07139_);
  or (_18909_, _18908_, _18907_);
  and (_18910_, _04670_, _05660_);
  or (_18911_, _18910_, _18849_);
  or (_18912_, _18911_, _07140_);
  and (_18913_, _18912_, _07150_);
  and (_18914_, _18913_, _18909_);
  and (_18915_, _18914_, _18905_);
  or (_18916_, _18915_, _18853_);
  and (_18918_, _18916_, _03138_);
  nand (_18919_, _18911_, _03022_);
  nor (_18920_, _18919_, _18861_);
  or (_18921_, _18849_, _05085_);
  and (_18922_, _18866_, _03137_);
  and (_18923_, _18922_, _18921_);
  or (_18924_, _18923_, _03042_);
  or (_18925_, _18924_, _18920_);
  or (_18926_, _18925_, _18918_);
  nor (_18927_, _10365_, _08691_);
  or (_18929_, _18849_, _03043_);
  or (_18930_, _18929_, _18927_);
  and (_18931_, _18930_, _07161_);
  and (_18932_, _18931_, _18926_);
  nor (_18933_, _10367_, _08691_);
  or (_18934_, _18933_, _18849_);
  and (_18935_, _18934_, _03143_);
  or (_18936_, _18935_, _03174_);
  or (_18937_, _18936_, _18932_);
  or (_18938_, _18863_, _03179_);
  and (_18940_, _18938_, _03183_);
  and (_18941_, _18940_, _18937_);
  and (_18942_, _18849_, _02799_);
  or (_18943_, _18942_, _02887_);
  or (_18944_, _18943_, _18941_);
  or (_18945_, _18863_, _02888_);
  and (_18946_, _18945_, _34655_);
  and (_18947_, _18946_, _18944_);
  or (_35840_[0], _18947_, _18848_);
  not (_18948_, \oc8051_golden_model_1.P3 [1]);
  nor (_18950_, _34655_, _18948_);
  or (_18951_, _18950_, rst);
  or (_18952_, _10565_, _08691_);
  or (_18953_, _04670_, \oc8051_golden_model_1.P3 [1]);
  and (_18954_, _18953_, _03148_);
  and (_18955_, _18954_, _18952_);
  and (_18956_, _16701_, _05337_);
  nor (_18957_, _05337_, _18948_);
  or (_18958_, _18957_, _02986_);
  or (_18959_, _18958_, _18956_);
  and (_18961_, _10574_, _04670_);
  not (_18962_, _18961_);
  and (_18963_, _18962_, _18953_);
  or (_18964_, _18963_, _03006_);
  nand (_18965_, _04670_, _02543_);
  and (_18966_, _18965_, _18953_);
  and (_18967_, _18966_, _03845_);
  nor (_18968_, _03845_, _18948_);
  or (_18969_, _18968_, _02948_);
  or (_18970_, _18969_, _18967_);
  and (_18972_, _18970_, _02976_);
  and (_18973_, _18972_, _18964_);
  nor (_18974_, _04670_, _18948_);
  nor (_18975_, _08691_, _04020_);
  or (_18976_, _18975_, _18974_);
  and (_18977_, _18976_, _02946_);
  and (_18978_, _10569_, _05337_);
  or (_18979_, _18978_, _18957_);
  and (_18980_, _18979_, _02884_);
  or (_18981_, _18980_, _18977_);
  or (_18983_, _18981_, _02880_);
  or (_18984_, _18983_, _18973_);
  or (_18985_, _18966_, _02992_);
  and (_18986_, _18985_, _18984_);
  or (_18987_, _18986_, _02877_);
  and (_18988_, _10572_, _05337_);
  or (_18989_, _18988_, _18957_);
  or (_18990_, _18989_, _02987_);
  and (_18991_, _18990_, _06246_);
  and (_18992_, _18991_, _18987_);
  and (_18994_, _18978_, _10568_);
  or (_18995_, _18994_, _18957_);
  and (_18996_, _18995_, _02871_);
  or (_18997_, _18996_, _02866_);
  or (_18998_, _18997_, _18992_);
  and (_18999_, _18998_, _18959_);
  or (_19000_, _18999_, _05535_);
  or (_19001_, _18976_, _02859_);
  and (_19002_, _19001_, _19000_);
  or (_19003_, _19002_, _02841_);
  and (_19005_, _06163_, _04670_);
  or (_19006_, _18974_, _02842_);
  or (_19007_, _19006_, _19005_);
  and (_19008_, _19007_, _02839_);
  and (_19009_, _19008_, _19003_);
  and (_19010_, _10674_, _04670_);
  or (_19011_, _19010_, _18974_);
  and (_19012_, _19011_, _02567_);
  or (_19013_, _19012_, _19009_);
  and (_19014_, _19013_, _03052_);
  or (_19016_, _10689_, _08691_);
  and (_19017_, _19016_, _03051_);
  nand (_19018_, _04670_, _03720_);
  and (_19019_, _19018_, _02834_);
  or (_19020_, _19019_, _19017_);
  and (_19021_, _19020_, _18953_);
  or (_19022_, _19021_, _19014_);
  and (_19023_, _19022_, _07150_);
  or (_19024_, _19023_, _18955_);
  and (_19025_, _19024_, _03138_);
  or (_19027_, _10688_, _08691_);
  and (_19028_, _18953_, _03022_);
  and (_19029_, _19028_, _19027_);
  or (_19030_, _18974_, _05038_);
  and (_19031_, _18966_, _03137_);
  and (_19032_, _19031_, _19030_);
  or (_19033_, _19032_, _19029_);
  or (_19034_, _19033_, _19025_);
  and (_19035_, _19034_, _03144_);
  or (_19036_, _18965_, _05038_);
  and (_19038_, _18953_, _03143_);
  and (_19039_, _19038_, _19036_);
  or (_19040_, _19039_, _03174_);
  or (_19041_, _19018_, _05038_);
  and (_19042_, _18953_, _03042_);
  and (_19043_, _19042_, _19041_);
  or (_19044_, _19043_, _19040_);
  or (_19045_, _19044_, _19035_);
  or (_19046_, _18963_, _03179_);
  and (_19047_, _19046_, _03183_);
  and (_19049_, _19047_, _19045_);
  and (_19050_, _18989_, _02799_);
  or (_19051_, _19050_, _02887_);
  or (_19052_, _19051_, _19049_);
  or (_19053_, _18974_, _02888_);
  or (_19054_, _19053_, _18961_);
  and (_19055_, _19054_, _34655_);
  and (_19056_, _19055_, _19052_);
  or (_35840_[1], _19056_, _18951_);
  not (_19057_, \oc8051_golden_model_1.P3 [2]);
  nor (_19059_, _34655_, _19057_);
  or (_19060_, _19059_, rst);
  nor (_19061_, _04670_, _19057_);
  nor (_19062_, _08691_, _04449_);
  or (_19063_, _19062_, _19061_);
  or (_19064_, _19063_, _02859_);
  nor (_19065_, _10788_, _08691_);
  or (_19066_, _19065_, _19061_);
  or (_19067_, _19066_, _03006_);
  and (_19068_, _04670_, \oc8051_golden_model_1.ACC [2]);
  or (_19070_, _19068_, _19061_);
  and (_19071_, _19070_, _03845_);
  nor (_19072_, _03845_, _19057_);
  or (_19073_, _19072_, _02948_);
  or (_19074_, _19073_, _19071_);
  and (_19075_, _19074_, _02976_);
  and (_19076_, _19075_, _19067_);
  and (_19077_, _19063_, _02946_);
  nor (_19078_, _05337_, _19057_);
  and (_19079_, _10792_, _05337_);
  or (_19081_, _19079_, _19078_);
  and (_19082_, _19081_, _02884_);
  or (_19083_, _19082_, _19077_);
  or (_19084_, _19083_, _02880_);
  or (_19085_, _19084_, _19076_);
  or (_19086_, _19070_, _02992_);
  and (_19087_, _19086_, _19085_);
  or (_19088_, _19087_, _02877_);
  and (_19089_, _10773_, _05337_);
  or (_19090_, _19089_, _19078_);
  or (_19092_, _19090_, _02987_);
  and (_19093_, _19092_, _06246_);
  and (_19094_, _19093_, _19088_);
  and (_19095_, _19079_, _10807_);
  or (_19096_, _19095_, _19078_);
  and (_19097_, _19096_, _02871_);
  or (_19098_, _19097_, _19094_);
  and (_19099_, _19098_, _02986_);
  and (_19100_, _16847_, _05337_);
  or (_19101_, _19078_, _19100_);
  and (_19103_, _19101_, _02866_);
  or (_19104_, _19103_, _05535_);
  or (_19105_, _19104_, _19099_);
  and (_19106_, _19105_, _19064_);
  or (_19107_, _19106_, _02841_);
  and (_19108_, _06167_, _04670_);
  or (_19109_, _19061_, _02842_);
  or (_19110_, _19109_, _19108_);
  and (_19111_, _19110_, _02839_);
  and (_19112_, _19111_, _19107_);
  nor (_19114_, _10881_, _08691_);
  or (_19115_, _19114_, _19061_);
  and (_19116_, _19115_, _02567_);
  or (_19117_, _19116_, _19112_);
  or (_19118_, _19117_, _08207_);
  and (_19119_, _10770_, _04670_);
  or (_19120_, _19061_, _07139_);
  or (_19121_, _19120_, _19119_);
  and (_19122_, _04670_, _05693_);
  or (_19123_, _19122_, _19061_);
  or (_19125_, _19123_, _07140_);
  and (_19126_, _19125_, _07150_);
  and (_19127_, _19126_, _19121_);
  and (_19128_, _19127_, _19118_);
  and (_19129_, _10766_, _04670_);
  or (_19130_, _19129_, _19061_);
  and (_19131_, _19130_, _03148_);
  or (_19132_, _19131_, _19128_);
  and (_19133_, _19132_, _03138_);
  or (_19134_, _19061_, _05135_);
  and (_19136_, _19070_, _03137_);
  and (_19137_, _19123_, _03022_);
  or (_19138_, _19137_, _19136_);
  and (_19139_, _19138_, _19134_);
  or (_19140_, _19139_, _03042_);
  or (_19141_, _19140_, _19133_);
  nor (_19142_, _10768_, _08691_);
  or (_19143_, _19061_, _03043_);
  or (_19144_, _19143_, _19142_);
  and (_19145_, _19144_, _07161_);
  and (_19147_, _19145_, _19141_);
  nor (_19148_, _10765_, _08691_);
  or (_19149_, _19148_, _19061_);
  and (_19150_, _19149_, _03143_);
  or (_19151_, _19150_, _03174_);
  or (_19152_, _19151_, _19147_);
  or (_19153_, _19066_, _03179_);
  and (_19154_, _19153_, _03183_);
  and (_19155_, _19154_, _19152_);
  and (_19156_, _19090_, _02799_);
  or (_19158_, _19156_, _02887_);
  or (_19159_, _19158_, _19155_);
  and (_19160_, _10941_, _04670_);
  or (_19161_, _19061_, _02888_);
  or (_19162_, _19161_, _19160_);
  and (_19163_, _19162_, _34655_);
  and (_19164_, _19163_, _19159_);
  or (_35840_[2], _19164_, _19060_);
  nor (_19165_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_19166_, _19165_, _04552_);
  and (_19168_, _08691_, \oc8051_golden_model_1.P3 [3]);
  nor (_19169_, _08691_, _04275_);
  or (_19170_, _19169_, _19168_);
  or (_19171_, _19170_, _02859_);
  and (_19172_, _16920_, _05337_);
  not (_19173_, _05337_);
  and (_19174_, _19173_, \oc8051_golden_model_1.P3 [3]);
  or (_19175_, _19174_, _02986_);
  or (_19176_, _19175_, _19172_);
  nor (_19177_, _10983_, _08691_);
  or (_19179_, _19177_, _19168_);
  or (_19180_, _19179_, _03006_);
  and (_19181_, _04670_, \oc8051_golden_model_1.ACC [3]);
  or (_19182_, _19181_, _19168_);
  and (_19183_, _19182_, _03845_);
  and (_19184_, _04194_, \oc8051_golden_model_1.P3 [3]);
  or (_19185_, _19184_, _02948_);
  or (_19186_, _19185_, _19183_);
  and (_19187_, _19186_, _02976_);
  and (_19188_, _19187_, _19180_);
  and (_19190_, _19170_, _02946_);
  and (_19191_, _10976_, _05337_);
  or (_19192_, _19191_, _19174_);
  and (_19193_, _19192_, _02884_);
  or (_19194_, _19193_, _19190_);
  or (_19195_, _19194_, _02880_);
  or (_19196_, _19195_, _19188_);
  or (_19197_, _19182_, _02992_);
  and (_19198_, _19197_, _19196_);
  or (_19199_, _19198_, _02877_);
  and (_19201_, _10979_, _05337_);
  or (_19202_, _19201_, _19174_);
  or (_19203_, _19202_, _02987_);
  and (_19204_, _19203_, _06246_);
  and (_19205_, _19204_, _19199_);
  or (_19206_, _19174_, _10975_);
  and (_19207_, _19206_, _02871_);
  and (_19208_, _19207_, _19192_);
  or (_19209_, _19208_, _02866_);
  or (_19210_, _19209_, _19205_);
  and (_19212_, _19210_, _19176_);
  or (_19213_, _19212_, _05535_);
  and (_19214_, _19213_, _19171_);
  or (_19215_, _19214_, _02841_);
  and (_19216_, _06166_, _04670_);
  or (_19217_, _19168_, _02842_);
  or (_19218_, _19217_, _19216_);
  and (_19219_, _19218_, _02839_);
  and (_19220_, _19219_, _19215_);
  nor (_19221_, _11076_, _08691_);
  or (_19223_, _19168_, _19221_);
  and (_19224_, _19223_, _02567_);
  or (_19225_, _19224_, _19220_);
  or (_19226_, _19225_, _08207_);
  and (_19227_, _10968_, _04670_);
  or (_19228_, _19168_, _07139_);
  or (_19229_, _19228_, _19227_);
  and (_19230_, _04670_, _05654_);
  or (_19231_, _19230_, _19168_);
  or (_19232_, _19231_, _07140_);
  and (_19234_, _19232_, _07150_);
  and (_19235_, _19234_, _19229_);
  and (_19236_, _19235_, _19226_);
  and (_19237_, _10964_, _04670_);
  or (_19238_, _19237_, _19168_);
  and (_19239_, _19238_, _03148_);
  or (_19240_, _19239_, _19236_);
  and (_19241_, _19240_, _03138_);
  or (_19242_, _19168_, _04993_);
  and (_19243_, _19182_, _03137_);
  and (_19245_, _19231_, _03022_);
  or (_19246_, _19245_, _19243_);
  and (_19247_, _19246_, _19242_);
  or (_19248_, _19247_, _03042_);
  or (_19249_, _19248_, _19241_);
  nor (_19250_, _10967_, _08691_);
  or (_19251_, _19168_, _03043_);
  or (_19252_, _19251_, _19250_);
  and (_19253_, _19252_, _07161_);
  and (_19254_, _19253_, _19249_);
  nor (_19256_, _10962_, _08691_);
  or (_19257_, _19256_, _19168_);
  and (_19258_, _19257_, _03143_);
  or (_19259_, _19258_, _03174_);
  or (_19260_, _19259_, _19254_);
  or (_19261_, _19179_, _03179_);
  and (_19262_, _19261_, _03183_);
  and (_19263_, _19262_, _19260_);
  and (_19264_, _19202_, _02799_);
  or (_19265_, _19264_, _02887_);
  or (_19267_, _19265_, _19263_);
  and (_19268_, _11136_, _04670_);
  or (_19269_, _19168_, _02888_);
  or (_19270_, _19269_, _19268_);
  and (_19271_, _19270_, _34655_);
  and (_19272_, _19271_, _19267_);
  or (_35840_[3], _19272_, _19166_);
  nor (_19273_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_19274_, _19273_, _04552_);
  and (_19275_, _08691_, \oc8051_golden_model_1.P3 [4]);
  nor (_19277_, _05192_, _08691_);
  or (_19278_, _19277_, _19275_);
  or (_19279_, _19278_, _02859_);
  and (_19280_, _19173_, \oc8051_golden_model_1.P3 [4]);
  and (_19281_, _11167_, _05337_);
  or (_19282_, _19281_, _19280_);
  or (_19283_, _19280_, _11201_);
  and (_19284_, _19283_, _02871_);
  and (_19285_, _19284_, _19282_);
  nor (_19286_, _11184_, _08691_);
  or (_19288_, _19286_, _19275_);
  or (_19289_, _19288_, _03006_);
  and (_19290_, _04670_, \oc8051_golden_model_1.ACC [4]);
  or (_19291_, _19290_, _19275_);
  and (_19292_, _19291_, _03845_);
  and (_19293_, _04194_, \oc8051_golden_model_1.P3 [4]);
  or (_19294_, _19293_, _02948_);
  or (_19295_, _19294_, _19292_);
  and (_19296_, _19295_, _02976_);
  and (_19297_, _19296_, _19289_);
  and (_19299_, _19278_, _02946_);
  and (_19300_, _19282_, _02884_);
  or (_19301_, _19300_, _19299_);
  or (_19302_, _19301_, _02880_);
  or (_19303_, _19302_, _19297_);
  or (_19304_, _19291_, _02992_);
  and (_19305_, _19304_, _19303_);
  or (_19306_, _19305_, _02877_);
  and (_19307_, _11165_, _05337_);
  or (_19308_, _19307_, _19280_);
  or (_19310_, _19308_, _02987_);
  and (_19311_, _19310_, _06246_);
  and (_19312_, _19311_, _19306_);
  or (_19313_, _19312_, _19285_);
  and (_19314_, _19313_, _02986_);
  and (_19315_, _17065_, _05337_);
  or (_19316_, _19315_, _19280_);
  and (_19317_, _19316_, _02866_);
  or (_19318_, _19317_, _05535_);
  or (_19319_, _19318_, _19314_);
  and (_19321_, _19319_, _19279_);
  or (_19322_, _19321_, _02841_);
  and (_19323_, _06171_, _04670_);
  or (_19324_, _19275_, _02842_);
  or (_19325_, _19324_, _19323_);
  and (_19326_, _19325_, _02839_);
  and (_19327_, _19326_, _19322_);
  nor (_19328_, _11271_, _08691_);
  or (_19329_, _19328_, _19275_);
  and (_19330_, _19329_, _02567_);
  or (_19332_, _19330_, _19327_);
  or (_19333_, _19332_, _08207_);
  and (_19334_, _11158_, _04670_);
  or (_19335_, _19275_, _07139_);
  or (_19336_, _19335_, _19334_);
  and (_19337_, _05618_, _04670_);
  or (_19338_, _19337_, _19275_);
  or (_19339_, _19338_, _07140_);
  and (_19340_, _19339_, _07150_);
  and (_19341_, _19340_, _19336_);
  and (_19343_, _19341_, _19333_);
  and (_19344_, _11154_, _04670_);
  or (_19345_, _19344_, _19275_);
  and (_19346_, _19345_, _03148_);
  or (_19347_, _19346_, _19343_);
  and (_19348_, _19347_, _03138_);
  or (_19349_, _19275_, _05240_);
  and (_19350_, _19291_, _03137_);
  and (_19351_, _19338_, _03022_);
  or (_19352_, _19351_, _19350_);
  and (_19354_, _19352_, _19349_);
  or (_19355_, _19354_, _03042_);
  or (_19356_, _19355_, _19348_);
  nor (_19357_, _11157_, _08691_);
  or (_19358_, _19275_, _03043_);
  or (_19359_, _19358_, _19357_);
  and (_19360_, _19359_, _07161_);
  and (_19361_, _19360_, _19356_);
  nor (_19362_, _11152_, _08691_);
  or (_19363_, _19362_, _19275_);
  and (_19365_, _19363_, _03143_);
  or (_19366_, _19365_, _03174_);
  or (_19367_, _19366_, _19361_);
  or (_19368_, _19288_, _03179_);
  and (_19369_, _19368_, _03183_);
  and (_19370_, _19369_, _19367_);
  and (_19371_, _19308_, _02799_);
  or (_19372_, _19371_, _02887_);
  or (_19373_, _19372_, _19370_);
  and (_19374_, _11338_, _04670_);
  or (_19376_, _19275_, _02888_);
  or (_19377_, _19376_, _19374_);
  and (_19378_, _19377_, _34655_);
  and (_19379_, _19378_, _19373_);
  or (_35840_[4], _19379_, _19274_);
  nor (_19380_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_19381_, _19380_, _04552_);
  and (_19382_, _19173_, \oc8051_golden_model_1.P3 [5]);
  and (_19383_, _11365_, _05337_);
  or (_19384_, _19383_, _19382_);
  or (_19386_, _19382_, _11397_);
  and (_19387_, _19386_, _02871_);
  and (_19388_, _19387_, _19384_);
  and (_19389_, _08691_, \oc8051_golden_model_1.P3 [5]);
  nor (_19390_, _11380_, _08691_);
  or (_19391_, _19390_, _19389_);
  or (_19392_, _19391_, _03006_);
  and (_19393_, _04670_, \oc8051_golden_model_1.ACC [5]);
  or (_19394_, _19393_, _19389_);
  and (_19395_, _19394_, _03845_);
  and (_19397_, _04194_, \oc8051_golden_model_1.P3 [5]);
  or (_19398_, _19397_, _02948_);
  or (_19399_, _19398_, _19395_);
  and (_19400_, _19399_, _02976_);
  and (_19401_, _19400_, _19392_);
  nor (_19402_, _04894_, _08691_);
  or (_19403_, _19402_, _19389_);
  and (_19404_, _19403_, _02946_);
  and (_19405_, _19384_, _02884_);
  or (_19406_, _19405_, _19404_);
  or (_19408_, _19406_, _02880_);
  or (_19409_, _19408_, _19401_);
  or (_19410_, _19394_, _02992_);
  and (_19411_, _19410_, _19409_);
  or (_19412_, _19411_, _02877_);
  and (_19413_, _11363_, _05337_);
  or (_19414_, _19413_, _19382_);
  or (_19415_, _19414_, _02987_);
  and (_19416_, _19415_, _06246_);
  and (_19417_, _19416_, _19412_);
  or (_19419_, _19417_, _19388_);
  and (_19420_, _19419_, _02986_);
  and (_19421_, _17171_, _05337_);
  or (_19422_, _19421_, _19382_);
  and (_19423_, _19422_, _02866_);
  or (_19424_, _19423_, _05535_);
  or (_19425_, _19424_, _19420_);
  or (_19426_, _19403_, _02859_);
  and (_19427_, _19426_, _19425_);
  or (_19428_, _19427_, _02841_);
  and (_19430_, _06170_, _04670_);
  or (_19431_, _19389_, _02842_);
  or (_19432_, _19431_, _19430_);
  and (_19433_, _19432_, _02839_);
  and (_19434_, _19433_, _19428_);
  nor (_19435_, _11467_, _08691_);
  or (_19436_, _19435_, _19389_);
  and (_19437_, _19436_, _02567_);
  or (_19438_, _19437_, _08207_);
  or (_19439_, _19438_, _19434_);
  and (_19441_, _11482_, _04670_);
  or (_19442_, _19389_, _07139_);
  or (_19443_, _19442_, _19441_);
  and (_19444_, _05671_, _04670_);
  or (_19445_, _19444_, _19389_);
  or (_19446_, _19445_, _07140_);
  and (_19447_, _19446_, _07150_);
  and (_19448_, _19447_, _19443_);
  and (_19449_, _19448_, _19439_);
  and (_19450_, _11356_, _04670_);
  or (_19452_, _19450_, _19389_);
  and (_19453_, _19452_, _03148_);
  or (_19454_, _19453_, _19449_);
  and (_19455_, _19454_, _03138_);
  or (_19456_, _19389_, _04945_);
  and (_19457_, _19394_, _03137_);
  and (_19458_, _19445_, _03022_);
  or (_19459_, _19458_, _19457_);
  and (_19460_, _19459_, _19456_);
  or (_19461_, _19460_, _03042_);
  or (_19463_, _19461_, _19455_);
  nor (_19464_, _11480_, _08691_);
  or (_19465_, _19389_, _03043_);
  or (_19466_, _19465_, _19464_);
  and (_19467_, _19466_, _07161_);
  and (_19468_, _19467_, _19463_);
  nor (_19469_, _11355_, _08691_);
  or (_19470_, _19469_, _19389_);
  and (_19471_, _19470_, _03143_);
  or (_19472_, _19471_, _03174_);
  or (_19474_, _19472_, _19468_);
  or (_19475_, _19391_, _03179_);
  and (_19476_, _19475_, _03183_);
  and (_19477_, _19476_, _19474_);
  and (_19478_, _19414_, _02799_);
  or (_19479_, _19478_, _02887_);
  or (_19480_, _19479_, _19477_);
  and (_19481_, _11541_, _04670_);
  or (_19482_, _19389_, _02888_);
  or (_19483_, _19482_, _19481_);
  and (_19485_, _19483_, _34655_);
  and (_19486_, _19485_, _19480_);
  or (_35840_[5], _19486_, _19381_);
  not (_19487_, \oc8051_golden_model_1.P3 [6]);
  nor (_19488_, _34655_, _19487_);
  or (_19489_, _19488_, rst);
  nor (_19490_, _05337_, _19487_);
  and (_19491_, _11564_, _05337_);
  or (_19492_, _19491_, _19490_);
  or (_19493_, _19490_, _11596_);
  and (_19495_, _19493_, _02871_);
  and (_19496_, _19495_, _19492_);
  nor (_19497_, _04670_, _19487_);
  nor (_19498_, _11567_, _08691_);
  or (_19499_, _19498_, _19497_);
  or (_19500_, _19499_, _03006_);
  and (_19501_, _04670_, \oc8051_golden_model_1.ACC [6]);
  or (_19502_, _19501_, _19497_);
  and (_19503_, _19502_, _03845_);
  nor (_19504_, _03845_, _19487_);
  or (_19506_, _19504_, _02948_);
  or (_19507_, _19506_, _19503_);
  and (_19508_, _19507_, _02976_);
  and (_19509_, _19508_, _19500_);
  nor (_19510_, _04790_, _08691_);
  or (_19511_, _19510_, _19497_);
  and (_19512_, _19511_, _02946_);
  and (_19513_, _19492_, _02884_);
  or (_19514_, _19513_, _19512_);
  or (_19515_, _19514_, _02880_);
  or (_19517_, _19515_, _19509_);
  or (_19518_, _19502_, _02992_);
  and (_19519_, _19518_, _19517_);
  or (_19520_, _19519_, _02877_);
  and (_19521_, _11562_, _05337_);
  or (_19522_, _19521_, _19490_);
  or (_19523_, _19522_, _02987_);
  and (_19524_, _19523_, _06246_);
  and (_19525_, _19524_, _19520_);
  or (_19526_, _19525_, _19496_);
  and (_19528_, _19526_, _02986_);
  and (_19529_, _17281_, _05337_);
  or (_19530_, _19529_, _19490_);
  and (_19531_, _19530_, _02866_);
  or (_19532_, _19531_, _05535_);
  or (_19533_, _19532_, _19528_);
  or (_19534_, _19511_, _02859_);
  and (_19535_, _19534_, _19533_);
  or (_19536_, _19535_, _02841_);
  and (_19537_, _06162_, _04670_);
  or (_19539_, _19497_, _02842_);
  or (_19540_, _19539_, _19537_);
  and (_19541_, _19540_, _02839_);
  and (_19542_, _19541_, _19536_);
  nor (_19543_, _11671_, _08691_);
  or (_19544_, _19543_, _19497_);
  and (_19545_, _19544_, _02567_);
  or (_19546_, _19545_, _08207_);
  or (_19547_, _19546_, _19542_);
  and (_19548_, _11560_, _04670_);
  or (_19550_, _19497_, _07139_);
  or (_19551_, _19550_, _19548_);
  and (_19552_, _11678_, _04670_);
  or (_19553_, _19552_, _19497_);
  or (_19554_, _19553_, _07140_);
  and (_19555_, _19554_, _07150_);
  and (_19556_, _19555_, _19551_);
  and (_19557_, _19556_, _19547_);
  and (_19558_, _11556_, _04670_);
  or (_19559_, _19558_, _19497_);
  and (_19561_, _19559_, _03148_);
  or (_19562_, _19561_, _19557_);
  and (_19563_, _19562_, _03138_);
  or (_19564_, _19497_, _04838_);
  and (_19565_, _19502_, _03137_);
  and (_19566_, _19553_, _03022_);
  or (_19567_, _19566_, _19565_);
  and (_19568_, _19567_, _19564_);
  or (_19569_, _19568_, _03042_);
  or (_19570_, _19569_, _19563_);
  nor (_19572_, _11558_, _08691_);
  or (_19573_, _19497_, _03043_);
  or (_19574_, _19573_, _19572_);
  and (_19575_, _19574_, _07161_);
  and (_19576_, _19575_, _19570_);
  nor (_19577_, _11555_, _08691_);
  or (_19578_, _19577_, _19497_);
  and (_19579_, _19578_, _03143_);
  or (_19580_, _19579_, _03174_);
  or (_19581_, _19580_, _19576_);
  or (_19583_, _19499_, _03179_);
  and (_19584_, _19583_, _03183_);
  and (_19585_, _19584_, _19581_);
  and (_19586_, _19522_, _02799_);
  or (_19587_, _19586_, _02887_);
  or (_19588_, _19587_, _19585_);
  and (_19589_, _11744_, _04670_);
  or (_19590_, _19497_, _02888_);
  or (_19591_, _19590_, _19589_);
  and (_19592_, _19591_, _34655_);
  and (_19594_, _19592_, _19588_);
  or (_35840_[6], _19594_, _19489_);
  and (_19595_, _08786_, _02247_);
  and (_19596_, _09692_, \oc8051_golden_model_1.PC [0]);
  and (_19597_, _03505_, \oc8051_golden_model_1.PC [0]);
  nor (_19598_, _19597_, _08896_);
  nor (_19599_, _19598_, _09692_);
  nor (_19600_, _19599_, _19596_);
  and (_19601_, _19600_, _02799_);
  and (_19602_, _09732_, _09724_);
  nor (_19604_, _19602_, _02247_);
  and (_19605_, _08803_, _08116_);
  nor (_19606_, _19605_, _02247_);
  not (_19607_, _08808_);
  nor (_19608_, _07763_, _02247_);
  and (_19609_, _07763_, _02247_);
  nor (_19610_, _19609_, _19608_);
  nor (_19611_, _19610_, _19607_);
  and (_19612_, _08815_, _03043_);
  nor (_19613_, _19612_, _02247_);
  not (_19615_, _02530_);
  and (_19616_, _09453_, _03023_);
  nor (_19617_, _19616_, _02247_);
  not (_19618_, _02524_);
  and (_19619_, _08823_, _07139_);
  nor (_19620_, _19619_, _02247_);
  not (_19621_, _09419_);
  not (_19622_, _09376_);
  and (_19623_, _02834_, _02247_);
  nor (_19624_, _03505_, _02589_);
  nor (_19626_, _09309_, _02247_);
  not (_19627_, _02589_);
  nor (_19628_, _03505_, _02591_);
  and (_19629_, _09200_, _09186_);
  nor (_19630_, _19629_, _02247_);
  nor (_19631_, _03505_, _02604_);
  not (_19632_, _07436_);
  and (_19633_, _09153_, _19632_);
  nor (_19634_, _19633_, _02247_);
  nor (_19635_, _19634_, _09169_);
  not (_19637_, _19635_);
  not (_19638_, _19633_);
  and (_19639_, _09145_, _02247_);
  nor (_19640_, _09145_, _02247_);
  nor (_19641_, _19640_, _19639_);
  and (_19642_, _19641_, _02603_);
  nor (_19643_, _19642_, _19638_);
  nor (_19644_, _19643_, _19637_);
  nor (_19645_, _19644_, _19631_);
  nor (_19646_, _19645_, _07433_);
  and (_19648_, _07433_, _02247_);
  nor (_19649_, _19648_, _09132_);
  not (_19650_, _19649_);
  nor (_19651_, _19650_, _19646_);
  nand (_19652_, _09011_, _09009_);
  and (_19653_, _02837_, _02247_);
  nor (_19654_, _19653_, _09073_);
  and (_19655_, _19654_, _19652_);
  and (_19656_, _05353_, _09010_);
  and (_19657_, _05351_, _05259_);
  and (_19659_, _19657_, _19656_);
  and (_19660_, _19659_, \oc8051_golden_model_1.PC [0]);
  or (_19661_, _19660_, _19655_);
  nor (_19662_, _19661_, _05361_);
  nor (_19663_, _19662_, _19651_);
  nor (_19664_, _19663_, _03840_);
  and (_19665_, _03840_, \oc8051_golden_model_1.PC [0]);
  nor (_19666_, _19665_, _02948_);
  not (_19667_, _19666_);
  nor (_19668_, _19667_, _19664_);
  not (_19670_, _19668_);
  nor (_19671_, _19598_, _09003_);
  and (_19672_, _05085_, _04992_);
  and (_19673_, _19672_, _09002_);
  and (_19674_, _19673_, _10785_);
  and (_19675_, _19674_, \oc8051_golden_model_1.PC [0]);
  or (_19676_, _19675_, _03006_);
  or (_19677_, _19676_, _19671_);
  and (_19678_, _19677_, _08997_);
  and (_19679_, _19678_, _19670_);
  nor (_19681_, _08997_, _02247_);
  nor (_19682_, _19681_, _04225_);
  not (_19683_, _19682_);
  nor (_19684_, _19683_, _19679_);
  nor (_19685_, _03505_, _02597_);
  not (_19686_, _19629_);
  nor (_19687_, _19686_, _19685_);
  not (_19688_, _19687_);
  nor (_19689_, _19688_, _19684_);
  or (_19690_, _19689_, _08989_);
  nor (_19692_, _19690_, _19630_);
  nor (_19693_, _03505_, _02595_);
  nor (_19694_, _19693_, _09210_);
  not (_19695_, _19694_);
  nor (_19696_, _19695_, _19692_);
  and (_19697_, _09242_, _02247_);
  not (_19698_, _19598_);
  nor (_19699_, _19698_, _09242_);
  or (_19700_, _19699_, _19697_);
  nor (_19701_, _19700_, _09209_);
  or (_19703_, _19701_, _08985_);
  nor (_19704_, _19703_, _19696_);
  or (_19705_, _19598_, _09918_);
  or (_19706_, _08981_, _02247_);
  and (_19707_, _19706_, _08985_);
  and (_19708_, _19707_, _19705_);
  or (_19709_, _19708_, _19704_);
  and (_19710_, _19709_, _09299_);
  and (_19711_, _09297_, _02247_);
  nor (_19712_, _19698_, _09297_);
  nor (_19714_, _19712_, _19711_);
  nor (_19715_, _19714_, _09299_);
  nor (_19716_, _19715_, _19710_);
  nor (_19717_, _19716_, _03029_);
  and (_19718_, _09276_, \oc8051_golden_model_1.PC [0]);
  nor (_19719_, _19598_, _09276_);
  or (_19720_, _19719_, _09279_);
  nor (_19721_, _19720_, _19718_);
  or (_19722_, _19721_, _19717_);
  and (_19723_, _19722_, _09250_);
  and (_19725_, _09249_, _02247_);
  or (_19726_, _19725_, _19723_);
  and (_19727_, _19726_, _02591_);
  or (_19728_, _19727_, _09310_);
  nor (_19729_, _19728_, _19628_);
  or (_19730_, _19729_, _19627_);
  nor (_19731_, _19730_, _19626_);
  and (_19732_, _09320_, _02571_);
  not (_19733_, _19732_);
  or (_19734_, _19733_, _19731_);
  nor (_19736_, _19734_, _19624_);
  nor (_19737_, _19732_, _02247_);
  nor (_19738_, _19737_, _02569_);
  not (_19739_, _19738_);
  nor (_19740_, _19739_, _19736_);
  nor (_19741_, _03505_, _04134_);
  and (_19742_, _09353_, _08211_);
  not (_19743_, _19742_);
  nor (_19744_, _19743_, _19741_);
  not (_19745_, _19744_);
  nor (_19747_, _19745_, _19740_);
  nor (_19748_, _19742_, _02247_);
  nor (_19749_, _19748_, _02516_);
  not (_19750_, _19749_);
  nor (_19751_, _19750_, _19747_);
  nor (_19752_, _03505_, _02517_);
  or (_19753_, _19752_, _09362_);
  or (_19754_, _19753_, _19751_);
  or (_19755_, _19654_, _09366_);
  and (_19756_, _19755_, _19754_);
  and (_19758_, _19756_, _07140_);
  or (_19759_, _19758_, _19623_);
  and (_19760_, _19759_, _19622_);
  and (_19761_, _09376_, _02689_);
  or (_19762_, _19761_, _19760_);
  and (_19763_, _19762_, _04131_);
  nor (_19764_, _03505_, _04131_);
  or (_19765_, _19764_, _19763_);
  and (_19766_, _19765_, _19621_);
  not (_19767_, _19619_);
  and (_19769_, _08166_, \oc8051_golden_model_1.PC [0]);
  and (_19770_, _19654_, _09447_);
  or (_19771_, _19770_, _19769_);
  and (_19772_, _19771_, _09419_);
  nor (_19773_, _19772_, _19767_);
  not (_19774_, _19773_);
  nor (_19775_, _19774_, _19766_);
  nor (_19776_, _19775_, _19620_);
  and (_19777_, _19776_, _19618_);
  nor (_19778_, _03505_, _19618_);
  or (_19780_, _19778_, _19777_);
  and (_19781_, _19780_, _09446_);
  not (_19782_, _19616_);
  nor (_19783_, _19654_, _09447_);
  nor (_19784_, _08166_, \oc8051_golden_model_1.PC [0]);
  nor (_19785_, _19784_, _09446_);
  not (_19786_, _19785_);
  nor (_19787_, _19786_, _19783_);
  nor (_19788_, _19787_, _19782_);
  not (_19789_, _19788_);
  nor (_19791_, _19789_, _19781_);
  nor (_19792_, _19791_, _19617_);
  and (_19793_, _19792_, _19615_);
  nor (_19794_, _03505_, _19615_);
  or (_19795_, _19794_, _19793_);
  and (_19796_, _19795_, _09470_);
  not (_19797_, _19612_);
  nor (_19798_, _19654_, \oc8051_golden_model_1.PSW [7]);
  and (_19799_, \oc8051_golden_model_1.PSW [7], _02247_);
  nor (_19800_, _19799_, _09470_);
  not (_19802_, _19800_);
  nor (_19803_, _19802_, _19798_);
  nor (_19804_, _19803_, _19797_);
  not (_19805_, _19804_);
  nor (_19806_, _19805_, _19796_);
  nor (_19807_, _19806_, _19613_);
  and (_19808_, _19807_, _02534_);
  nor (_19809_, _03505_, _02534_);
  or (_19810_, _19809_, _19808_);
  and (_19811_, _19810_, _19607_);
  and (_19813_, _08806_, _07996_);
  not (_19814_, _19813_);
  or (_19815_, _19814_, _19811_);
  nor (_19816_, _19815_, _19611_);
  nor (_19817_, _19813_, _02247_);
  nor (_19818_, _19817_, _03155_);
  not (_19819_, _19818_);
  nor (_19820_, _19819_, _19816_);
  and (_19821_, _06164_, _03155_);
  or (_19822_, _19821_, _19820_);
  and (_19824_, _19822_, _05790_);
  nor (_19825_, _03505_, _05790_);
  or (_19826_, _19825_, _19824_);
  and (_19827_, _19826_, _03223_);
  not (_19828_, _19605_);
  and (_19829_, _19698_, _09692_);
  nor (_19830_, _09692_, _02247_);
  or (_19831_, _19830_, _03223_);
  nor (_19832_, _19831_, _19829_);
  nor (_19833_, _19832_, _19828_);
  not (_19835_, _19833_);
  nor (_19836_, _19835_, _19827_);
  nor (_19837_, _19836_, _19606_);
  and (_19838_, _19837_, _02891_);
  and (_19839_, _06164_, _02890_);
  or (_19840_, _19839_, _19838_);
  and (_19841_, _19840_, _08788_);
  nor (_19842_, _03505_, _08788_);
  nor (_19843_, _19842_, _19841_);
  nor (_19844_, _19843_, _02889_);
  not (_19846_, _19602_);
  and (_19847_, _19600_, _02889_);
  nor (_19848_, _19847_, _19846_);
  not (_19849_, _19848_);
  nor (_19850_, _19849_, _19844_);
  nor (_19851_, _19850_, _19604_);
  nor (_19852_, _19851_, _04150_);
  and (_19853_, _04150_, _03505_);
  nor (_19854_, _19853_, _02799_);
  not (_19855_, _19854_);
  nor (_19857_, _19855_, _19852_);
  nor (_19858_, _19857_, _19601_);
  and (_19859_, _09755_, _09747_);
  not (_19860_, _19859_);
  nor (_19861_, _19860_, _19858_);
  nor (_19862_, _03036_, _02499_);
  not (_19863_, _19862_);
  nor (_19864_, _19859_, \oc8051_golden_model_1.PC [0]);
  nor (_19865_, _19864_, _19863_);
  not (_19866_, _19865_);
  nor (_19868_, _19866_, _19861_);
  and (_19869_, _19863_, _03505_);
  nor (_19870_, _19869_, _08786_);
  not (_19871_, _19870_);
  nor (_19872_, _19871_, _19868_);
  nor (_19873_, _19872_, _19595_);
  nand (_19874_, _19873_, _34655_);
  or (_19875_, _34655_, \oc8051_golden_model_1.PC [0]);
  and (_19876_, _19875_, _35796_);
  and (_35842_[0], _19876_, _19874_);
  and (_19878_, _08786_, _08894_);
  and (_19879_, _02887_, _02220_);
  and (_19880_, _03608_, _03297_);
  and (_19881_, _05256_, _02544_);
  or (_19882_, _19881_, _19880_);
  and (_19883_, _03174_, _02220_);
  nor (_19884_, _03299_, _03271_);
  and (_19885_, _19884_, _04520_);
  nor (_19886_, _19885_, _08894_);
  nor (_19887_, _08806_, _08894_);
  nor (_19889_, _08815_, _08894_);
  nor (_19890_, _09453_, _08894_);
  nor (_19891_, _08823_, _08894_);
  nor (_19892_, _09320_, _08894_);
  nor (_19893_, _09262_, _02220_);
  nand (_19894_, _09003_, _02544_);
  nor (_19895_, _08898_, _08896_);
  nor (_19896_, _19895_, _08899_);
  not (_19897_, _19896_);
  or (_19898_, _19897_, _09003_);
  nand (_19900_, _19898_, _19894_);
  nand (_19901_, _19900_, _02948_);
  nor (_19902_, _09075_, _09073_);
  nor (_19903_, _19902_, _09076_);
  and (_19904_, _19903_, _19652_);
  and (_19905_, _09012_, _02220_);
  nor (_19906_, _19905_, _19904_);
  nand (_19907_, _19906_, _09132_);
  and (_19908_, _03840_, _02544_);
  nor (_19909_, _19908_, _02948_);
  and (_19911_, _07436_, _02544_);
  nor (_19912_, _03720_, _02603_);
  not (_19913_, _09151_);
  and (_19914_, _09138_, \oc8051_golden_model_1.PC [0]);
  nor (_19915_, _19914_, _03845_);
  nor (_19916_, _19915_, _02220_);
  and (_19917_, _19915_, _02220_);
  or (_19918_, _19917_, _19916_);
  nor (_19919_, _19918_, _07423_);
  nor (_19920_, _09134_, _08894_);
  nor (_19922_, _19920_, _09135_);
  nor (_19923_, _19922_, _19919_);
  and (_19924_, _09134_, _02544_);
  nor (_19925_, _19924_, _03849_);
  not (_19926_, _19925_);
  nor (_19927_, _19926_, _19923_);
  nor (_19928_, _19927_, _19913_);
  not (_19929_, _19928_);
  nor (_19930_, _19929_, _19912_);
  nor (_19931_, _09151_, _08894_);
  not (_19933_, _19931_);
  and (_19934_, _19933_, _07420_);
  not (_19935_, _19934_);
  nor (_19936_, _19935_, _19930_);
  nor (_19937_, _07420_, _02544_);
  nor (_19938_, _19937_, _07410_);
  not (_19939_, _19938_);
  nor (_19940_, _19939_, _19936_);
  and (_19941_, _07410_, _02544_);
  nor (_19942_, _19941_, _02951_);
  not (_19944_, _19942_);
  nor (_19945_, _19944_, _19940_);
  and (_19946_, _02951_, _02220_);
  or (_19947_, _19946_, _07436_);
  nor (_19948_, _19947_, _19945_);
  or (_19949_, _19948_, _09169_);
  nor (_19950_, _19949_, _19911_);
  nor (_19951_, _03720_, _02601_);
  nor (_19952_, _19951_, _19950_);
  nor (_19953_, _19952_, _07433_);
  and (_19955_, _07433_, _08894_);
  nor (_19956_, _19955_, _03840_);
  nand (_19957_, _19956_, _05361_);
  or (_19958_, _19957_, _19953_);
  and (_19959_, _19958_, _19909_);
  nand (_19960_, _19959_, _19907_);
  and (_19961_, _19960_, _08997_);
  nand (_19962_, _19961_, _19901_);
  nor (_19963_, _08997_, _08894_);
  nor (_19964_, _19963_, _02884_);
  nand (_19966_, _19964_, _19962_);
  and (_19967_, _02884_, _02220_);
  nor (_19968_, _19967_, _04225_);
  nand (_19969_, _19968_, _19966_);
  and (_19970_, _03720_, _04225_);
  nor (_19971_, _19970_, _02946_);
  nand (_19972_, _19971_, _19969_);
  and (_19973_, _02946_, _02220_);
  nor (_19974_, _19973_, _09187_);
  nand (_19975_, _19974_, _19972_);
  nor (_19977_, _09186_, _08894_);
  nor (_19978_, _19977_, _02880_);
  nand (_19979_, _19978_, _19975_);
  and (_19980_, _02880_, _02220_);
  nor (_19981_, _19980_, _09193_);
  nand (_19982_, _19981_, _19979_);
  and (_19983_, _09193_, _02544_);
  nor (_19984_, _19983_, _02877_);
  nand (_19985_, _19984_, _19982_);
  and (_19986_, _02595_, \oc8051_golden_model_1.PC [1]);
  or (_19988_, _19986_, _08990_);
  nand (_19989_, _19988_, _19985_);
  and (_19990_, _03720_, _08989_);
  nor (_19991_, _19990_, _02876_);
  nand (_19992_, _19991_, _19989_);
  and (_19993_, _02876_, _02220_);
  nor (_19994_, _19993_, _09210_);
  nand (_19995_, _19994_, _19992_);
  and (_19996_, _09242_, _02544_);
  nor (_19997_, _19897_, _09242_);
  or (_19999_, _19997_, _19996_);
  nor (_20000_, _19999_, _09209_);
  nor (_20001_, _20000_, _08985_);
  nand (_20002_, _20001_, _19995_);
  or (_20003_, _19897_, _09918_);
  or (_20004_, _08981_, _08894_);
  nand (_20005_, _20004_, _20003_);
  nand (_20006_, _20005_, _08985_);
  and (_20007_, _20006_, _09299_);
  nand (_20008_, _20007_, _20002_);
  nor (_20010_, _19897_, _09297_);
  not (_20011_, _20010_);
  and (_20012_, _09297_, _02544_);
  nor (_20013_, _20012_, _09299_);
  and (_20014_, _20013_, _20011_);
  nor (_20015_, _20014_, _03029_);
  nand (_20016_, _20015_, _20008_);
  and (_20017_, _09276_, _08894_);
  nor (_20018_, _19896_, _09276_);
  or (_20019_, _20018_, _09279_);
  or (_20021_, _20019_, _20017_);
  and (_20022_, _20021_, _09250_);
  and (_20023_, _20022_, _20016_);
  and (_20024_, _09249_, _02544_);
  or (_20025_, _20024_, _20023_);
  nand (_20026_, _20025_, _06246_);
  and (_20027_, _02871_, \oc8051_golden_model_1.PC [1]);
  nor (_20028_, _20027_, _09257_);
  nand (_20029_, _20028_, _20026_);
  not (_20030_, _09262_);
  nor (_20032_, _03720_, _02591_);
  nor (_20033_, _20032_, _20030_);
  and (_20034_, _20033_, _20029_);
  or (_20035_, _20034_, _19893_);
  nand (_20036_, _20035_, _09309_);
  nor (_20037_, _09309_, _08894_);
  nor (_20038_, _20037_, _02941_);
  nand (_20039_, _20038_, _20036_);
  and (_20040_, _02941_, _02220_);
  nor (_20041_, _20040_, _19627_);
  nand (_20043_, _20041_, _20039_);
  and (_20044_, _03720_, _19627_);
  nor (_20045_, _20044_, _02940_);
  nand (_20046_, _20045_, _20043_);
  and (_20047_, _02940_, _02220_);
  nor (_20048_, _20047_, _09326_);
  and (_20049_, _20048_, _20046_);
  or (_20050_, _20049_, _19892_);
  nand (_20051_, _20050_, _09324_);
  nor (_20052_, _09324_, _02220_);
  nor (_20054_, _20052_, _07721_);
  and (_20055_, _20054_, _20051_);
  nor (_20056_, _02571_, _02544_);
  or (_20057_, _20056_, _02866_);
  nor (_20058_, _20057_, _20055_);
  and (_20059_, _02866_, \oc8051_golden_model_1.PC [1]);
  or (_20060_, _20059_, _20058_);
  nand (_20061_, _20060_, _04134_);
  and (_20062_, _03720_, _02569_);
  nor (_20063_, _20062_, _03046_);
  nand (_20064_, _20063_, _20061_);
  and (_20065_, _02860_, _08894_);
  or (_20066_, _20065_, _09345_);
  nand (_20067_, _20066_, _20064_);
  nor (_20068_, _02860_, _02220_);
  nor (_20069_, _20068_, _02567_);
  and (_20070_, _20069_, _20067_);
  nor (_20071_, _09352_, _02544_);
  nor (_20072_, _20071_, _09353_);
  or (_20073_, _20072_, _20070_);
  and (_20075_, _09352_, _02544_);
  nor (_20076_, _20075_, _02930_);
  nand (_20077_, _20076_, _20073_);
  and (_20078_, _02930_, _02220_);
  nor (_20079_, _20078_, _02516_);
  nand (_20080_, _20079_, _20077_);
  and (_20081_, _03720_, _02516_);
  nor (_20082_, _20081_, _09362_);
  nand (_20083_, _20082_, _20080_);
  and (_20084_, _19903_, _09362_);
  nor (_20086_, _20084_, _05749_);
  nand (_20087_, _20086_, _20083_);
  nor (_20088_, _05748_, _02220_);
  nor (_20089_, _20088_, _02834_);
  and (_20090_, _20089_, _20087_);
  and (_20091_, _02834_, _02544_);
  or (_20092_, _20091_, _07830_);
  nor (_20093_, _20092_, _20090_);
  and (_20094_, _07830_, \oc8051_golden_model_1.PC [1]);
  or (_20095_, _20094_, _20093_);
  nand (_20097_, _20095_, _19622_);
  nor (_20098_, _19622_, _02674_);
  nor (_20099_, _20098_, _02928_);
  nand (_20100_, _20099_, _20097_);
  and (_20101_, _02928_, _02220_);
  nor (_20102_, _20101_, _02522_);
  nand (_20103_, _20102_, _20100_);
  and (_20104_, _03720_, _02522_);
  nor (_20105_, _20104_, _09419_);
  nand (_20106_, _20105_, _20103_);
  and (_20107_, _08166_, _02220_);
  and (_20108_, _19903_, _09447_);
  or (_20109_, _20108_, _20107_);
  and (_20110_, _20109_, _09419_);
  nor (_20111_, _20110_, _09428_);
  and (_20112_, _20111_, _20106_);
  or (_20113_, _20112_, _19891_);
  nand (_20114_, _20113_, _08822_);
  nor (_20115_, _08822_, _02220_);
  nor (_20116_, _20115_, _03051_);
  and (_20118_, _20116_, _20114_);
  and (_20119_, _03051_, _02544_);
  or (_20120_, _20119_, _03148_);
  nor (_20121_, _20120_, _20118_);
  and (_20122_, _03148_, \oc8051_golden_model_1.PC [1]);
  or (_20123_, _20122_, _20121_);
  nand (_20124_, _20123_, _19618_);
  and (_20125_, _03720_, _02524_);
  nor (_20126_, _20125_, _09441_);
  nand (_20127_, _20126_, _20124_);
  not (_20129_, _09453_);
  nor (_20130_, _19903_, _09447_);
  nor (_20131_, _08166_, _02220_);
  nor (_20132_, _20131_, _09446_);
  not (_20133_, _20132_);
  nor (_20134_, _20133_, _20130_);
  nor (_20135_, _20134_, _20129_);
  and (_20136_, _20135_, _20127_);
  or (_20137_, _20136_, _19890_);
  nand (_20138_, _20137_, _09455_);
  nor (_20139_, _09455_, _02220_);
  nor (_20140_, _20139_, _03022_);
  and (_20141_, _20140_, _20138_);
  and (_20142_, _03022_, _02544_);
  or (_20143_, _20142_, _03137_);
  nor (_20144_, _20143_, _20141_);
  and (_20145_, _03137_, \oc8051_golden_model_1.PC [1]);
  or (_20146_, _20145_, _20144_);
  nand (_20147_, _20146_, _19615_);
  and (_20148_, _03720_, _02530_);
  nor (_20150_, _20148_, _08818_);
  nand (_20151_, _20150_, _20147_);
  nor (_20152_, _19903_, \oc8051_golden_model_1.PSW [7]);
  and (_20153_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor (_20154_, _20153_, _09470_);
  not (_20155_, _20154_);
  nor (_20156_, _20155_, _20152_);
  nor (_20157_, _20156_, _09468_);
  and (_20158_, _20157_, _20151_);
  or (_20159_, _20158_, _19889_);
  nand (_20161_, _20159_, _08812_);
  nor (_20162_, _08812_, _02220_);
  nor (_20163_, _20162_, _03042_);
  and (_20164_, _20163_, _20161_);
  and (_20165_, _03042_, _02544_);
  or (_20166_, _20165_, _03143_);
  nor (_20167_, _20166_, _20164_);
  and (_20168_, _03143_, \oc8051_golden_model_1.PC [1]);
  or (_20169_, _20168_, _20167_);
  nand (_20170_, _20169_, _02534_);
  and (_20171_, _03720_, _02533_);
  nor (_20172_, _20171_, _08808_);
  nand (_20173_, _20172_, _20170_);
  nor (_20174_, _19903_, _07288_);
  and (_20175_, _07288_, \oc8051_golden_model_1.PC [1]);
  nor (_20176_, _20175_, _19607_);
  not (_20177_, _20176_);
  nor (_20178_, _20177_, _20174_);
  nor (_20179_, _20178_, _09487_);
  and (_20180_, _20179_, _20173_);
  or (_20182_, _20180_, _19887_);
  nand (_20183_, _20182_, _07965_);
  nor (_20184_, _07965_, _02220_);
  nor (_20185_, _20184_, _07995_);
  and (_20186_, _20185_, _20183_);
  and (_20187_, _07995_, _08894_);
  or (_20188_, _20187_, _03155_);
  nor (_20189_, _20188_, _20186_);
  and (_20190_, _05900_, _03155_);
  or (_20191_, _20190_, _20189_);
  nand (_20193_, _20191_, _05790_);
  and (_20194_, _03720_, _02528_);
  nor (_20195_, _20194_, _03040_);
  nand (_20196_, _20195_, _20193_);
  not (_20197_, _07186_);
  and (_20198_, _19897_, _09692_);
  not (_20199_, _20198_);
  nor (_20200_, _09692_, _02544_);
  nor (_20201_, _20200_, _03223_);
  and (_20202_, _20201_, _20199_);
  nor (_20203_, _20202_, _20197_);
  nand (_20204_, _20203_, _20196_);
  nor (_20205_, _07186_, _08894_);
  and (_20206_, _08031_, _07188_);
  not (_20207_, _20206_);
  nor (_20208_, _20207_, _20205_);
  nand (_20209_, _20208_, _20204_);
  nor (_20210_, _20206_, _02544_);
  nor (_20211_, _20210_, _08112_);
  nand (_20212_, _20211_, _20209_);
  and (_20214_, _08112_, \oc8051_golden_model_1.PC [1]);
  nor (_20215_, _20214_, _08115_);
  nand (_20216_, _20215_, _20212_);
  and (_20217_, _08115_, _08894_);
  nor (_20218_, _20217_, _02890_);
  and (_20219_, _20218_, _20216_);
  and (_20220_, _05900_, _02890_);
  or (_20221_, _20220_, _20219_);
  nand (_20222_, _20221_, _08788_);
  and (_20223_, _03720_, _02510_);
  nor (_20225_, _20223_, _02889_);
  nand (_20226_, _20225_, _20222_);
  not (_20227_, _19885_);
  and (_20228_, _09692_, _08894_);
  nor (_20229_, _19896_, _09692_);
  nor (_20230_, _20229_, _20228_);
  and (_20231_, _20230_, _02889_);
  nor (_20232_, _20231_, _20227_);
  and (_20233_, _20232_, _20226_);
  or (_20234_, _20233_, _19886_);
  and (_20235_, _04522_, _05809_);
  nand (_20236_, _20235_, _20234_);
  nor (_20237_, _20235_, _08894_);
  nor (_20238_, _20237_, _03174_);
  and (_20239_, _20238_, _20236_);
  or (_20240_, _20239_, _19883_);
  nand (_20241_, _20240_, _09732_);
  nor (_20242_, _09732_, _02544_);
  nor (_20243_, _20242_, _04150_);
  nand (_20244_, _20243_, _20241_);
  and (_20246_, _04150_, _03720_);
  nor (_20247_, _20246_, _02799_);
  nand (_20248_, _20247_, _20244_);
  and (_20249_, _20230_, _02799_);
  nor (_20250_, _20249_, _05256_);
  and (_20251_, _20250_, _20248_);
  or (_20252_, _20251_, _19882_);
  and (_20253_, _19880_, _08894_);
  not (_20254_, _20253_);
  and (_20255_, _02962_, _02498_);
  nor (_20257_, _10743_, _20255_);
  and (_20258_, _20257_, _20254_);
  nand (_20259_, _20258_, _20252_);
  nor (_20260_, _20257_, _08894_);
  nor (_20261_, _20260_, _02887_);
  and (_20262_, _20261_, _20259_);
  or (_20263_, _20262_, _19879_);
  nand (_20264_, _20263_, _09755_);
  nor (_20265_, _09755_, _02544_);
  nor (_20266_, _20265_, _19863_);
  nand (_20267_, _20266_, _20264_);
  and (_20268_, _19863_, _03720_);
  nor (_20269_, _20268_, _08786_);
  and (_20270_, _20269_, _20267_);
  or (_20271_, _20270_, _19878_);
  or (_20272_, _20271_, _34659_);
  or (_20273_, _34655_, \oc8051_golden_model_1.PC [1]);
  and (_20274_, _20273_, _35796_);
  and (_35842_[1], _20274_, _20272_);
  and (_20275_, _08786_, _02553_);
  and (_20277_, _19863_, _03262_);
  nand (_20278_, _03174_, _02614_);
  nor (_20279_, _08803_, _02553_);
  nor (_20280_, _08806_, _02553_);
  nor (_20281_, _08815_, _02553_);
  nor (_20282_, _09453_, _02553_);
  nor (_20283_, _08823_, _02553_);
  nor (_20284_, _02858_, _02614_);
  and (_20285_, _02866_, _02620_);
  nor (_20286_, _09320_, _02553_);
  nor (_20288_, _09262_, _02614_);
  not (_20289_, _02553_);
  and (_20290_, _09249_, _20289_);
  and (_20291_, _08903_, _08900_);
  nor (_20292_, _20291_, _08904_);
  not (_20293_, _20292_);
  or (_20294_, _20293_, _09918_);
  nand (_20295_, _09918_, _08891_);
  and (_20296_, _20295_, _20294_);
  and (_20297_, _20296_, _08985_);
  nor (_20298_, _20292_, _09003_);
  and (_20299_, _09003_, _08892_);
  or (_20300_, _20299_, _20298_);
  and (_20301_, _20300_, _02948_);
  and (_20302_, _09080_, _09077_);
  nor (_20303_, _20302_, _09081_);
  nand (_20304_, _20303_, _19652_);
  nand (_20305_, _19659_, _02614_);
  and (_20306_, _20305_, _20304_);
  and (_20307_, _20306_, _09132_);
  or (_20309_, _03262_, _02601_);
  or (_20310_, _03262_, _02603_);
  nand (_20311_, _03845_, _02614_);
  and (_20312_, _20311_, _09135_);
  nor (_20313_, _09138_, \oc8051_golden_model_1.PC [2]);
  or (_20314_, _20313_, _03845_);
  and (_20315_, _20314_, _20312_);
  nor (_20316_, _09145_, _02553_);
  or (_20317_, _20316_, _03849_);
  or (_20318_, _20317_, _20315_);
  and (_20320_, _20318_, _09153_);
  and (_20321_, _20320_, _20310_);
  nor (_20322_, _09153_, _02553_);
  or (_20323_, _20322_, _02951_);
  or (_20324_, _20323_, _20321_);
  and (_20325_, _02951_, _02614_);
  nor (_20326_, _20325_, _07436_);
  and (_20327_, _20326_, _20324_);
  and (_20328_, _07436_, _20289_);
  or (_20329_, _20328_, _09169_);
  or (_20330_, _20329_, _20327_);
  and (_20331_, _20330_, _20309_);
  or (_20332_, _20331_, _07433_);
  nand (_20333_, _07433_, _02553_);
  and (_20334_, _20333_, _05361_);
  and (_20335_, _20334_, _20332_);
  or (_20336_, _20335_, _03840_);
  or (_20337_, _20336_, _20307_);
  nand (_20338_, _03840_, _02553_);
  and (_20339_, _20338_, _03006_);
  and (_20341_, _20339_, _20337_);
  or (_20342_, _20341_, _20301_);
  and (_20343_, _20342_, _08997_);
  nor (_20344_, _08997_, _02553_);
  or (_20345_, _20344_, _02884_);
  or (_20346_, _20345_, _20343_);
  nand (_20347_, _02884_, _02614_);
  and (_20348_, _20347_, _02597_);
  and (_20349_, _20348_, _20346_);
  and (_20350_, _03262_, _04225_);
  or (_20352_, _20350_, _02946_);
  or (_20353_, _20352_, _20349_);
  nand (_20354_, _02946_, _02614_);
  and (_20355_, _20354_, _09186_);
  and (_20356_, _20355_, _20353_);
  nor (_20357_, _09186_, _02553_);
  or (_20358_, _20357_, _02880_);
  or (_20359_, _20358_, _20356_);
  and (_20360_, _02880_, _02614_);
  nor (_20361_, _20360_, _09193_);
  and (_20362_, _20361_, _20359_);
  and (_20363_, _09193_, _20289_);
  or (_20364_, _20363_, _02877_);
  or (_20365_, _20364_, _20362_);
  nand (_20366_, _02877_, _02614_);
  and (_20367_, _20366_, _02595_);
  and (_20368_, _20367_, _20365_);
  and (_20369_, _03262_, _08989_);
  or (_20370_, _20369_, _02876_);
  or (_20371_, _20370_, _20368_);
  nand (_20373_, _02876_, _02614_);
  and (_20374_, _20373_, _09209_);
  and (_20375_, _20374_, _20371_);
  nor (_20376_, _20292_, _09242_);
  and (_20377_, _09242_, _08892_);
  or (_20378_, _20377_, _20376_);
  and (_20379_, _20378_, _09210_);
  or (_20380_, _20379_, _20375_);
  and (_20381_, _20380_, _08986_);
  or (_20382_, _20381_, _20297_);
  and (_20384_, _20382_, _09299_);
  nand (_20385_, _09297_, _08891_);
  or (_20386_, _20293_, _09297_);
  and (_20387_, _20386_, _02954_);
  and (_20388_, _20387_, _20385_);
  or (_20389_, _20388_, _03029_);
  or (_20390_, _20389_, _20384_);
  nor (_20391_, _20292_, _09276_);
  and (_20392_, _09276_, _08892_);
  or (_20393_, _20392_, _09279_);
  or (_20394_, _20393_, _20391_);
  and (_20395_, _20394_, _09250_);
  and (_20396_, _20395_, _20390_);
  or (_20397_, _20396_, _20290_);
  and (_20398_, _20397_, _06246_);
  and (_20399_, _02871_, _02620_);
  or (_20400_, _20399_, _09257_);
  or (_20401_, _20400_, _20398_);
  or (_20402_, _03262_, _02591_);
  and (_20403_, _20402_, _09262_);
  and (_20405_, _20403_, _20401_);
  or (_20406_, _20405_, _20288_);
  and (_20407_, _20406_, _09309_);
  nor (_20408_, _09309_, _02553_);
  or (_20409_, _20408_, _02941_);
  or (_20410_, _20409_, _20407_);
  nand (_20411_, _02941_, _02614_);
  and (_20412_, _20411_, _02589_);
  and (_20413_, _20412_, _20410_);
  and (_20414_, _03262_, _19627_);
  or (_20416_, _20414_, _02940_);
  or (_20417_, _20416_, _20413_);
  nand (_20418_, _02940_, _02614_);
  and (_20419_, _20418_, _09320_);
  and (_20420_, _20419_, _20417_);
  or (_20421_, _20420_, _20286_);
  and (_20422_, _20421_, _09324_);
  nor (_20423_, _09324_, _02614_);
  or (_20424_, _20423_, _07721_);
  or (_20425_, _20424_, _20422_);
  nor (_20426_, _20289_, _02571_);
  nor (_20427_, _20426_, _02866_);
  and (_20428_, _20427_, _20425_);
  or (_20429_, _20428_, _20285_);
  and (_20430_, _20429_, _04134_);
  and (_20431_, _03262_, _02569_);
  or (_20432_, _20431_, _03046_);
  or (_20433_, _20432_, _20430_);
  nand (_20434_, _08891_, _03046_);
  and (_20435_, _20434_, _02858_);
  and (_20437_, _20435_, _20433_);
  or (_20438_, _20437_, _20284_);
  and (_20439_, _20438_, _04195_);
  nor (_20440_, _04195_, _02614_);
  or (_20441_, _20440_, _02567_);
  or (_20442_, _20441_, _20439_);
  and (_20443_, _08891_, _02567_);
  nor (_20444_, _20443_, _09352_);
  and (_20445_, _20444_, _20442_);
  and (_20446_, _09352_, _20289_);
  or (_20448_, _20446_, _02930_);
  or (_20449_, _20448_, _20445_);
  nand (_20450_, _02930_, _02614_);
  and (_20451_, _20450_, _02517_);
  and (_20452_, _20451_, _20449_);
  and (_20453_, _03262_, _02516_);
  or (_20454_, _20453_, _09362_);
  or (_20455_, _20454_, _20452_);
  nand (_20456_, _20303_, _09362_);
  and (_20457_, _05747_, _02620_);
  or (_20458_, _20457_, _05748_);
  and (_20459_, _20458_, _20456_);
  and (_20460_, _20459_, _20455_);
  nor (_20461_, _05748_, _02614_);
  or (_20462_, _20461_, _20460_);
  and (_20463_, _20462_, _07140_);
  and (_20464_, _08892_, _02834_);
  or (_20465_, _20464_, _07830_);
  or (_20466_, _20465_, _20463_);
  nand (_20467_, _07830_, _02614_);
  and (_20469_, _20467_, _19622_);
  and (_20470_, _20469_, _20466_);
  and (_20471_, _09376_, _02585_);
  or (_20472_, _20471_, _02928_);
  or (_20473_, _20472_, _20470_);
  nand (_20474_, _02928_, _02614_);
  and (_20475_, _20474_, _04131_);
  and (_20476_, _20475_, _20473_);
  and (_20477_, _03262_, _02522_);
  or (_20478_, _20477_, _09419_);
  or (_20480_, _20478_, _20476_);
  nor (_20481_, _20303_, _08166_);
  nand (_20482_, _08166_, _02620_);
  nand (_20483_, _20482_, _09419_);
  or (_20484_, _20483_, _20481_);
  and (_20485_, _20484_, _08823_);
  and (_20486_, _20485_, _20480_);
  or (_20487_, _20486_, _20283_);
  and (_20488_, _20487_, _08822_);
  nor (_20489_, _08822_, _02614_);
  or (_20491_, _20489_, _03051_);
  or (_20492_, _20491_, _20488_);
  nand (_20493_, _08891_, _03051_);
  and (_20494_, _20493_, _07150_);
  and (_20495_, _20494_, _20492_);
  and (_20496_, _03148_, _02620_);
  or (_20497_, _20496_, _20495_);
  and (_20498_, _20497_, _19618_);
  and (_20499_, _03262_, _02524_);
  or (_20500_, _20499_, _09441_);
  or (_20501_, _20500_, _20498_);
  nor (_20502_, _20303_, _09447_);
  or (_20503_, _08166_, _02614_);
  nand (_20504_, _20503_, _09441_);
  or (_20505_, _20504_, _20502_);
  and (_20506_, _20505_, _09453_);
  and (_20507_, _20506_, _20501_);
  or (_20508_, _20507_, _20282_);
  and (_20509_, _20508_, _09455_);
  nor (_20510_, _09455_, _02614_);
  or (_20512_, _20510_, _03022_);
  or (_20513_, _20512_, _20509_);
  nand (_20514_, _08891_, _03022_);
  and (_20515_, _20514_, _06213_);
  and (_20516_, _20515_, _20513_);
  and (_20517_, _03137_, _02620_);
  or (_20518_, _20517_, _20516_);
  and (_20519_, _20518_, _19615_);
  and (_20520_, _03262_, _02530_);
  or (_20521_, _20520_, _08818_);
  or (_20523_, _20521_, _20519_);
  nor (_20524_, _20303_, \oc8051_golden_model_1.PSW [7]);
  or (_20525_, _02614_, _07288_);
  nand (_20526_, _20525_, _08818_);
  or (_20527_, _20526_, _20524_);
  and (_20528_, _20527_, _08815_);
  and (_20529_, _20528_, _20523_);
  or (_20530_, _20529_, _20281_);
  and (_20531_, _20530_, _08812_);
  nor (_20532_, _08812_, _02614_);
  or (_20533_, _20532_, _03042_);
  or (_20534_, _20533_, _20531_);
  nand (_20535_, _08891_, _03042_);
  and (_20536_, _20535_, _07161_);
  and (_20537_, _20536_, _20534_);
  and (_20538_, _03143_, _02620_);
  or (_20539_, _20538_, _20537_);
  and (_20540_, _20539_, _02534_);
  and (_20541_, _03262_, _02533_);
  or (_20542_, _20541_, _08808_);
  or (_20544_, _20542_, _20540_);
  or (_20545_, _20303_, _07288_);
  or (_20546_, _02614_, \oc8051_golden_model_1.PSW [7]);
  and (_20547_, _20546_, _08808_);
  and (_20548_, _20547_, _20545_);
  nor (_20549_, _20548_, _09487_);
  and (_20550_, _20549_, _20544_);
  or (_20551_, _20550_, _20280_);
  and (_20552_, _20551_, _07965_);
  nor (_20553_, _07965_, _02614_);
  or (_20555_, _20553_, _07995_);
  or (_20556_, _20555_, _20552_);
  not (_20557_, _03155_);
  nand (_20558_, _07995_, _02553_);
  and (_20559_, _20558_, _20557_);
  and (_20560_, _20559_, _20556_);
  and (_20561_, _06036_, _03155_);
  or (_20562_, _20561_, _20560_);
  and (_20563_, _20562_, _05790_);
  and (_20564_, _03262_, _02528_);
  or (_20566_, _20564_, _03040_);
  or (_20567_, _20566_, _20563_);
  nor (_20568_, _09692_, _08891_);
  and (_20569_, _20293_, _09692_);
  or (_20570_, _20569_, _03223_);
  or (_20571_, _20570_, _20568_);
  and (_20572_, _20571_, _08803_);
  and (_20573_, _20572_, _20567_);
  or (_20574_, _20573_, _20279_);
  and (_20575_, _20574_, _08789_);
  and (_20576_, _08112_, _02620_);
  or (_20577_, _20576_, _08115_);
  or (_20578_, _20577_, _20575_);
  nand (_20579_, _08115_, _02553_);
  and (_20580_, _20579_, _02891_);
  and (_20581_, _20580_, _20578_);
  and (_20582_, _06036_, _02890_);
  or (_20583_, _20582_, _20581_);
  and (_20584_, _20583_, _08788_);
  and (_20585_, _03262_, _02510_);
  or (_20587_, _20585_, _02889_);
  or (_20588_, _20587_, _20584_);
  nor (_20589_, _20292_, _09692_);
  and (_20590_, _09692_, _08892_);
  nor (_20591_, _20590_, _20589_);
  nand (_20592_, _20591_, _02889_);
  and (_20593_, _20592_, _09724_);
  and (_20594_, _20593_, _20588_);
  nor (_20595_, _09724_, _02553_);
  or (_20596_, _20595_, _03174_);
  or (_20598_, _20596_, _20594_);
  and (_20599_, _20598_, _20278_);
  nor (_20600_, _20599_, _09733_);
  nor (_20601_, _09732_, _20289_);
  nor (_20602_, _20601_, _04150_);
  not (_20603_, _20602_);
  nor (_20604_, _20603_, _20600_);
  and (_20605_, _04150_, _03262_);
  nor (_20606_, _20605_, _02799_);
  not (_20607_, _20606_);
  nor (_20608_, _20607_, _20604_);
  and (_20609_, _09747_, _03183_);
  nor (_20610_, _20591_, _09748_);
  nor (_20611_, _20610_, _20609_);
  nor (_20612_, _20611_, _20608_);
  nor (_20613_, _09747_, _02553_);
  nor (_20614_, _20613_, _02887_);
  not (_20615_, _20614_);
  nor (_20616_, _20615_, _20612_);
  and (_20617_, _09755_, _02888_);
  and (_20619_, _09755_, _02620_);
  nor (_20620_, _20619_, _20617_);
  nor (_20621_, _20620_, _20616_);
  nor (_20622_, _09755_, _02553_);
  nor (_20623_, _20622_, _20621_);
  nor (_20624_, _20623_, _19863_);
  or (_20625_, _20624_, _08786_);
  nor (_20626_, _20625_, _20277_);
  nor (_20627_, _20626_, _20275_);
  nand (_20628_, _20627_, _34655_);
  or (_20630_, _34655_, \oc8051_golden_model_1.PC [2]);
  and (_20631_, _20630_, _35796_);
  and (_35842_[2], _20631_, _20628_);
  and (_20632_, _08786_, _02636_);
  and (_20633_, _19863_, _03128_);
  nand (_20634_, _03174_, _02640_);
  nor (_20635_, _08803_, _02636_);
  and (_20636_, _05991_, _03155_);
  nor (_20637_, _08806_, _02636_);
  nor (_20638_, _08815_, _02636_);
  nor (_20640_, _09453_, _02636_);
  nor (_20641_, _08823_, _02636_);
  and (_20642_, _02866_, _02661_);
  nor (_20643_, _09320_, _02636_);
  nor (_20644_, _09262_, _02640_);
  and (_20645_, _09249_, _02628_);
  nand (_20646_, _09918_, _08886_);
  or (_20647_, _08889_, _08888_);
  and (_20648_, _20647_, _08905_);
  nor (_20649_, _20647_, _08905_);
  nor (_20651_, _20649_, _20648_);
  not (_20652_, _20651_);
  or (_20653_, _20652_, _09918_);
  and (_20654_, _20653_, _20646_);
  and (_20655_, _20654_, _08985_);
  nand (_20656_, _09242_, _08886_);
  or (_20657_, _20652_, _09242_);
  and (_20658_, _20657_, _20656_);
  and (_20659_, _20658_, _09210_);
  and (_20660_, _09003_, _08887_);
  nor (_20662_, _20651_, _09003_);
  or (_20663_, _20662_, _20660_);
  and (_20664_, _20663_, _02948_);
  or (_20665_, _09070_, _09069_);
  and (_20666_, _20665_, _09082_);
  nor (_20667_, _20665_, _09082_);
  nor (_20668_, _20667_, _20666_);
  nand (_20669_, _20668_, _19652_);
  nand (_20670_, _19659_, _02640_);
  and (_20671_, _20670_, _20669_);
  and (_20673_, _20671_, _09132_);
  or (_20674_, _03128_, _02601_);
  or (_20675_, _03128_, _02603_);
  nand (_20676_, _03845_, _02640_);
  and (_20677_, _20676_, _09135_);
  nor (_20678_, _09138_, \oc8051_golden_model_1.PC [3]);
  or (_20679_, _20678_, _03845_);
  and (_20680_, _20679_, _20677_);
  nor (_20681_, _09145_, _02636_);
  or (_20682_, _20681_, _03849_);
  or (_20684_, _20682_, _20680_);
  and (_20685_, _20684_, _09153_);
  and (_20686_, _20685_, _20675_);
  nor (_20687_, _09153_, _02636_);
  or (_20688_, _20687_, _02951_);
  or (_20689_, _20688_, _20686_);
  and (_20690_, _02951_, _02640_);
  nor (_20691_, _20690_, _07436_);
  and (_20692_, _20691_, _20689_);
  and (_20693_, _07436_, _02628_);
  or (_20695_, _20693_, _09169_);
  or (_20696_, _20695_, _20692_);
  and (_20697_, _20696_, _20674_);
  or (_20698_, _20697_, _07433_);
  nand (_20699_, _07433_, _02636_);
  and (_20700_, _20699_, _05361_);
  and (_20701_, _20700_, _20698_);
  or (_20702_, _20701_, _03840_);
  or (_20703_, _20702_, _20673_);
  nand (_20704_, _03840_, _02636_);
  and (_20706_, _20704_, _03006_);
  and (_20707_, _20706_, _20703_);
  or (_20708_, _20707_, _20664_);
  and (_20709_, _20708_, _08997_);
  nor (_20710_, _08997_, _02636_);
  or (_20711_, _20710_, _02884_);
  or (_20712_, _20711_, _20709_);
  nand (_20713_, _02884_, _02640_);
  and (_20714_, _20713_, _02597_);
  and (_20715_, _20714_, _20712_);
  and (_20716_, _03128_, _04225_);
  or (_20717_, _20716_, _02946_);
  or (_20718_, _20717_, _20715_);
  nand (_20719_, _02946_, _02640_);
  and (_20720_, _20719_, _09186_);
  and (_20721_, _20720_, _20718_);
  nor (_20722_, _09186_, _02636_);
  or (_20723_, _20722_, _02880_);
  or (_20724_, _20723_, _20721_);
  and (_20725_, _02880_, _02640_);
  nor (_20726_, _20725_, _09193_);
  and (_20727_, _20726_, _20724_);
  and (_20728_, _09193_, _02628_);
  or (_20729_, _20728_, _02877_);
  or (_20730_, _20729_, _20727_);
  nand (_20731_, _02877_, _02640_);
  and (_20732_, _20731_, _02595_);
  and (_20733_, _20732_, _20730_);
  and (_20734_, _03128_, _08989_);
  or (_20735_, _20734_, _02876_);
  or (_20737_, _20735_, _20733_);
  nand (_20738_, _02876_, _02640_);
  and (_20739_, _20738_, _09209_);
  and (_20740_, _20739_, _20737_);
  or (_20741_, _20740_, _20659_);
  and (_20742_, _20741_, _08986_);
  or (_20743_, _20742_, _20655_);
  and (_20744_, _20743_, _09299_);
  or (_20745_, _20652_, _09297_);
  nand (_20746_, _09297_, _08886_);
  and (_20748_, _20746_, _02954_);
  and (_20749_, _20748_, _20745_);
  or (_20750_, _20749_, _03029_);
  or (_20751_, _20750_, _20744_);
  nor (_20752_, _20651_, _09276_);
  and (_20753_, _09276_, _08887_);
  or (_20754_, _20753_, _09279_);
  or (_20755_, _20754_, _20752_);
  and (_20756_, _20755_, _09250_);
  and (_20757_, _20756_, _20751_);
  or (_20759_, _20757_, _20645_);
  and (_20760_, _20759_, _06246_);
  and (_20761_, _02871_, _02661_);
  or (_20762_, _20761_, _09257_);
  or (_20763_, _20762_, _20760_);
  or (_20764_, _03128_, _02591_);
  and (_20765_, _20764_, _09262_);
  and (_20766_, _20765_, _20763_);
  or (_20767_, _20766_, _20644_);
  and (_20768_, _20767_, _09309_);
  nor (_20770_, _09309_, _02636_);
  or (_20771_, _20770_, _02941_);
  or (_20772_, _20771_, _20768_);
  nand (_20773_, _02941_, _02640_);
  and (_20774_, _20773_, _02589_);
  and (_20775_, _20774_, _20772_);
  and (_20776_, _03128_, _19627_);
  or (_20777_, _20776_, _02940_);
  or (_20778_, _20777_, _20775_);
  nand (_20779_, _02940_, _02640_);
  and (_20781_, _20779_, _09320_);
  and (_20782_, _20781_, _20778_);
  or (_20783_, _20782_, _20643_);
  and (_20784_, _20783_, _09324_);
  nor (_20785_, _09324_, _02640_);
  or (_20786_, _20785_, _07721_);
  or (_20787_, _20786_, _20784_);
  nor (_20788_, _02571_, _02628_);
  nor (_20789_, _20788_, _02866_);
  and (_20790_, _20789_, _20787_);
  or (_20792_, _20790_, _20642_);
  and (_20793_, _20792_, _04134_);
  and (_20794_, _03128_, _02569_);
  or (_20795_, _20794_, _03046_);
  or (_20796_, _20795_, _20793_);
  nand (_20797_, _08886_, _03046_);
  and (_20798_, _20797_, _02860_);
  and (_20799_, _20798_, _20796_);
  nor (_20800_, _02860_, _02640_);
  or (_20801_, _20800_, _02567_);
  or (_20803_, _20801_, _20799_);
  nor (_20804_, _09352_, _08886_);
  or (_20805_, _20804_, _09353_);
  and (_20806_, _20805_, _20803_);
  and (_20807_, _09352_, _02628_);
  or (_20808_, _20807_, _02930_);
  or (_20809_, _20808_, _20806_);
  nand (_20810_, _02930_, _02640_);
  and (_20811_, _20810_, _02517_);
  and (_20812_, _20811_, _20809_);
  and (_20814_, _03128_, _02516_);
  or (_20815_, _20814_, _09362_);
  or (_20816_, _20815_, _20812_);
  nand (_20817_, _20668_, _09362_);
  and (_20818_, _20817_, _05748_);
  and (_20819_, _20818_, _20816_);
  nor (_20820_, _05748_, _02640_);
  or (_20821_, _20820_, _02834_);
  or (_20822_, _20821_, _20819_);
  nand (_20823_, _08886_, _02834_);
  and (_20825_, _20823_, _07831_);
  and (_20826_, _20825_, _20822_);
  and (_20827_, _07830_, _02661_);
  or (_20828_, _20827_, _20826_);
  and (_20829_, _20828_, _19622_);
  and (_20830_, _09376_, _02652_);
  or (_20831_, _20830_, _02928_);
  or (_20832_, _20831_, _20829_);
  nand (_20833_, _02928_, _02640_);
  and (_20834_, _20833_, _04131_);
  and (_20836_, _20834_, _20832_);
  and (_20837_, _03128_, _02522_);
  or (_20838_, _20837_, _09419_);
  or (_20839_, _20838_, _20836_);
  nor (_20840_, _20668_, _08166_);
  nand (_20841_, _08166_, _02661_);
  nand (_20842_, _20841_, _09419_);
  or (_20843_, _20842_, _20840_);
  and (_20844_, _20843_, _08823_);
  and (_20845_, _20844_, _20839_);
  or (_20847_, _20845_, _20641_);
  and (_20848_, _20847_, _08822_);
  nor (_20849_, _08822_, _02640_);
  or (_20850_, _20849_, _03051_);
  or (_20851_, _20850_, _20848_);
  nand (_20852_, _08886_, _03051_);
  and (_20853_, _20852_, _07150_);
  and (_20854_, _20853_, _20851_);
  and (_20855_, _03148_, _02661_);
  or (_20856_, _20855_, _20854_);
  and (_20858_, _20856_, _19618_);
  and (_20859_, _03128_, _02524_);
  or (_20860_, _20859_, _09441_);
  or (_20861_, _20860_, _20858_);
  nor (_20862_, _20668_, _09447_);
  or (_20863_, _08166_, _02640_);
  nand (_20864_, _20863_, _09441_);
  or (_20865_, _20864_, _20862_);
  and (_20866_, _20865_, _09453_);
  and (_20867_, _20866_, _20861_);
  or (_20869_, _20867_, _20640_);
  and (_20870_, _20869_, _09455_);
  nor (_20871_, _09455_, _02640_);
  or (_20872_, _20871_, _03022_);
  or (_20873_, _20872_, _20870_);
  nand (_20874_, _08886_, _03022_);
  and (_20875_, _20874_, _06213_);
  and (_20876_, _20875_, _20873_);
  and (_20877_, _03137_, _02661_);
  or (_20878_, _20877_, _20876_);
  and (_20880_, _20878_, _19615_);
  and (_20881_, _03128_, _02530_);
  or (_20882_, _20881_, _08818_);
  or (_20883_, _20882_, _20880_);
  nor (_20884_, _20668_, \oc8051_golden_model_1.PSW [7]);
  or (_20885_, _02640_, _07288_);
  nand (_20886_, _20885_, _08818_);
  or (_20887_, _20886_, _20884_);
  and (_20888_, _20887_, _08815_);
  and (_20889_, _20888_, _20883_);
  or (_20891_, _20889_, _20638_);
  and (_20892_, _20891_, _08812_);
  nor (_20893_, _08812_, _02640_);
  or (_20894_, _20893_, _03042_);
  or (_20895_, _20894_, _20892_);
  nand (_20896_, _08886_, _03042_);
  and (_20897_, _20896_, _07161_);
  and (_20898_, _20897_, _20895_);
  and (_20899_, _03143_, _02661_);
  or (_20900_, _20899_, _20898_);
  and (_20902_, _20900_, _02534_);
  and (_20903_, _03128_, _02533_);
  or (_20904_, _20903_, _08808_);
  or (_20905_, _20904_, _20902_);
  or (_20906_, _20668_, _07288_);
  or (_20907_, _02640_, \oc8051_golden_model_1.PSW [7]);
  and (_20908_, _20907_, _08808_);
  and (_20909_, _20908_, _20906_);
  nor (_20910_, _20909_, _09487_);
  and (_20911_, _20910_, _20905_);
  or (_20913_, _20911_, _20637_);
  and (_20914_, _20913_, _07965_);
  nor (_20915_, _07965_, _02640_);
  or (_20916_, _20915_, _07995_);
  or (_20917_, _20916_, _20914_);
  nand (_20918_, _07995_, _02636_);
  and (_20919_, _20918_, _20557_);
  and (_20920_, _20919_, _20917_);
  or (_20921_, _20920_, _20636_);
  and (_20922_, _20921_, _05790_);
  and (_20924_, _03128_, _02528_);
  or (_20925_, _20924_, _03040_);
  or (_20926_, _20925_, _20922_);
  nor (_20927_, _09692_, _08886_);
  and (_20928_, _20652_, _09692_);
  or (_20929_, _20928_, _03223_);
  or (_20930_, _20929_, _20927_);
  and (_20931_, _20930_, _08803_);
  and (_20932_, _20931_, _20926_);
  or (_20933_, _20932_, _20635_);
  and (_20935_, _20933_, _08789_);
  and (_20936_, _08112_, _02661_);
  or (_20937_, _20936_, _08115_);
  or (_20938_, _20937_, _20935_);
  nand (_20939_, _08115_, _02636_);
  and (_20940_, _20939_, _02891_);
  and (_20941_, _20940_, _20938_);
  and (_20942_, _05991_, _02890_);
  or (_20943_, _20942_, _20941_);
  and (_20944_, _20943_, _08788_);
  and (_20946_, _03128_, _02510_);
  or (_20947_, _20946_, _02889_);
  or (_20948_, _20947_, _20944_);
  and (_20949_, _09692_, _08887_);
  nor (_20950_, _20651_, _09692_);
  nor (_20951_, _20950_, _20949_);
  nand (_20952_, _20951_, _02889_);
  and (_20953_, _20952_, _09724_);
  and (_20954_, _20953_, _20948_);
  nor (_20955_, _09724_, _02636_);
  or (_20957_, _20955_, _03174_);
  or (_20958_, _20957_, _20954_);
  and (_20959_, _20958_, _20634_);
  nor (_20960_, _20959_, _09733_);
  nor (_20961_, _09732_, _02628_);
  nor (_20962_, _20961_, _04150_);
  not (_20963_, _20962_);
  nor (_20964_, _20963_, _20960_);
  and (_20965_, _04150_, _03128_);
  nor (_20966_, _20965_, _02799_);
  not (_20968_, _20966_);
  nor (_20969_, _20968_, _20964_);
  nor (_20970_, _20951_, _09748_);
  nor (_20971_, _20970_, _20609_);
  nor (_20972_, _20971_, _20969_);
  nor (_20973_, _09747_, _02636_);
  nor (_20974_, _20973_, _02887_);
  not (_20975_, _20974_);
  nor (_20976_, _20975_, _20972_);
  and (_20977_, _09755_, _02661_);
  nor (_20979_, _20977_, _20617_);
  nor (_20980_, _20979_, _20976_);
  nor (_20981_, _09755_, _02636_);
  nor (_20982_, _20981_, _20980_);
  nor (_20983_, _20982_, _19863_);
  or (_20984_, _20983_, _08786_);
  nor (_20985_, _20984_, _20633_);
  or (_20986_, _20985_, _20632_);
  or (_20987_, _20986_, _34659_);
  or (_20988_, _34655_, \oc8051_golden_model_1.PC [3]);
  and (_20990_, _20988_, _35796_);
  and (_35842_[3], _20990_, _20987_);
  not (_20991_, \oc8051_golden_model_1.PC [4]);
  nor (_20992_, _02234_, _20991_);
  and (_20993_, _02234_, _20991_);
  nor (_20994_, _20993_, _20992_);
  and (_20995_, _20994_, _08786_);
  not (_20996_, _20994_);
  nor (_20997_, _20996_, _09755_);
  nand (_20998_, _20996_, _09249_);
  nand (_21000_, _09067_, _02877_);
  or (_21001_, _20994_, _09186_);
  and (_21002_, _08910_, _08907_);
  nor (_21003_, _21002_, _08911_);
  not (_21004_, _21003_);
  nor (_21005_, _21004_, _09003_);
  and (_21006_, _09003_, _08882_);
  or (_21007_, _21006_, _21005_);
  and (_21008_, _21007_, _02948_);
  nor (_21009_, _09087_, _09085_);
  nor (_21011_, _21009_, _09088_);
  and (_21012_, _21011_, _19652_);
  and (_21013_, _09012_, _09066_);
  or (_21014_, _21013_, _21012_);
  or (_21015_, _21014_, _05361_);
  and (_21016_, _05617_, _03849_);
  nand (_21017_, _09067_, _03845_);
  nand (_21018_, _21017_, _09135_);
  or (_21019_, _09138_, _20991_);
  and (_21020_, _21019_, _04194_);
  or (_21022_, _21020_, _21018_);
  or (_21023_, _20996_, _09145_);
  and (_21024_, _21023_, _02603_);
  and (_21025_, _21024_, _21022_);
  or (_21026_, _21025_, _09154_);
  or (_21027_, _21026_, _21016_);
  or (_21028_, _20996_, _09153_);
  and (_21029_, _21028_, _03401_);
  and (_21030_, _21029_, _21027_);
  and (_21031_, _09067_, _02951_);
  or (_21033_, _21031_, _21030_);
  nand (_21034_, _21033_, _19632_);
  nand (_21035_, _20996_, _07436_);
  and (_21036_, _21035_, _21034_);
  or (_21037_, _21036_, _09169_);
  nand (_21038_, _05617_, _09169_);
  and (_21039_, _21038_, _09133_);
  and (_21040_, _21039_, _21037_);
  nand (_21041_, _20994_, _07433_);
  nand (_21042_, _21041_, _05361_);
  or (_21044_, _21042_, _21040_);
  and (_21045_, _21044_, _09176_);
  and (_21046_, _21045_, _21015_);
  or (_21047_, _21046_, _21008_);
  and (_21048_, _21047_, _08997_);
  and (_21049_, _20994_, _09181_);
  or (_21050_, _21049_, _02884_);
  or (_21051_, _21050_, _21048_);
  nand (_21052_, _09067_, _02884_);
  and (_21053_, _21052_, _02597_);
  and (_21055_, _21053_, _21051_);
  nor (_21056_, _05617_, _02597_);
  or (_21057_, _21056_, _02946_);
  or (_21058_, _21057_, _21055_);
  nand (_21059_, _09067_, _02946_);
  and (_21060_, _21059_, _21058_);
  or (_21061_, _21060_, _09187_);
  and (_21062_, _21061_, _21001_);
  or (_21063_, _21062_, _02880_);
  and (_21064_, _09067_, _02880_);
  nor (_21066_, _21064_, _09193_);
  and (_21067_, _21066_, _21063_);
  and (_21068_, _20994_, _09193_);
  or (_21069_, _21068_, _02877_);
  or (_21070_, _21069_, _21067_);
  and (_21071_, _21070_, _21000_);
  or (_21072_, _21071_, _08989_);
  nand (_21073_, _05617_, _08989_);
  and (_21074_, _21073_, _03962_);
  and (_21075_, _21074_, _21072_);
  nand (_21077_, _09066_, _02876_);
  nand (_21078_, _21077_, _09209_);
  or (_21079_, _21078_, _21075_);
  and (_21080_, _09242_, _08882_);
  nor (_21081_, _21004_, _09242_);
  or (_21082_, _21081_, _21080_);
  or (_21083_, _21082_, _09209_);
  and (_21084_, _21083_, _21079_);
  or (_21085_, _21084_, _08985_);
  and (_21086_, _21003_, _08981_);
  and (_21088_, _09918_, _08882_);
  or (_21089_, _21088_, _08986_);
  or (_21090_, _21089_, _21086_);
  and (_21091_, _21090_, _21085_);
  or (_21092_, _21091_, _02954_);
  nor (_21093_, _21004_, _09297_);
  and (_21094_, _09297_, _08882_);
  or (_21095_, _21094_, _09299_);
  or (_21096_, _21095_, _21093_);
  and (_21097_, _21096_, _09279_);
  and (_21099_, _21097_, _21092_);
  or (_21100_, _21003_, _09276_);
  nand (_21101_, _09276_, _08883_);
  and (_21102_, _21101_, _03029_);
  and (_21103_, _21102_, _21100_);
  or (_21104_, _21103_, _09249_);
  or (_21105_, _21104_, _21099_);
  and (_21106_, _21105_, _20998_);
  or (_21107_, _21106_, _02871_);
  nand (_21108_, _09067_, _02871_);
  and (_21110_, _21108_, _02591_);
  and (_21111_, _21110_, _21107_);
  nor (_21112_, _05617_, _02591_);
  or (_21113_, _21112_, _20030_);
  or (_21114_, _21113_, _21111_);
  or (_21115_, _09262_, _09066_);
  and (_21116_, _21115_, _09309_);
  and (_21117_, _21116_, _21114_);
  nor (_21118_, _20996_, _09309_);
  or (_21119_, _21118_, _02941_);
  or (_21121_, _21119_, _21117_);
  nand (_21122_, _09067_, _02941_);
  and (_21123_, _21122_, _21121_);
  or (_21124_, _21123_, _19627_);
  nand (_21125_, _05617_, _19627_);
  and (_21126_, _21125_, _10030_);
  and (_21127_, _21126_, _21124_);
  and (_21128_, _09066_, _02940_);
  or (_21129_, _21128_, _21127_);
  and (_21130_, _21129_, _09320_);
  nor (_21132_, _20996_, _09320_);
  or (_21133_, _21132_, _09325_);
  or (_21134_, _21133_, _21130_);
  or (_21135_, _09324_, _09066_);
  and (_21136_, _21135_, _02571_);
  and (_21137_, _21136_, _21134_);
  nor (_21138_, _20996_, _02571_);
  or (_21139_, _21138_, _02866_);
  or (_21140_, _21139_, _21137_);
  nand (_21141_, _09067_, _02866_);
  and (_21143_, _21141_, _21140_);
  or (_21144_, _21143_, _02569_);
  nand (_21145_, _05617_, _02569_);
  and (_21146_, _21145_, _08211_);
  and (_21147_, _21146_, _21144_);
  nand (_21148_, _08882_, _03046_);
  nand (_21149_, _21148_, _02860_);
  or (_21150_, _21149_, _21147_);
  or (_21151_, _09066_, _02860_);
  and (_21152_, _21151_, _02839_);
  and (_21154_, _21152_, _21150_);
  nor (_21155_, _09352_, _08882_);
  nor (_21156_, _21155_, _09353_);
  or (_21157_, _21156_, _21154_);
  nand (_21158_, _20996_, _09352_);
  and (_21159_, _21158_, _03508_);
  and (_21160_, _21159_, _21157_);
  and (_21161_, _09066_, _02930_);
  or (_21162_, _21161_, _02516_);
  or (_21163_, _21162_, _21160_);
  nand (_21165_, _05617_, _02516_);
  and (_21166_, _21165_, _09366_);
  and (_21167_, _21166_, _21163_);
  and (_21168_, _21011_, _09362_);
  or (_21169_, _21168_, _05749_);
  or (_21170_, _21169_, _21167_);
  or (_21171_, _09066_, _05748_);
  and (_21172_, _21171_, _07140_);
  and (_21173_, _21172_, _21170_);
  and (_21174_, _08882_, _02834_);
  or (_21176_, _21174_, _07830_);
  or (_21177_, _21176_, _21173_);
  nand (_21178_, _09067_, _07830_);
  and (_21179_, _21178_, _21177_);
  or (_21180_, _21179_, _09376_);
  and (_21181_, _09395_, _09392_);
  nor (_21182_, _21181_, _09396_);
  or (_21183_, _21182_, _19622_);
  and (_21184_, _21183_, _09778_);
  and (_21185_, _21184_, _21180_);
  and (_21187_, _09066_, _02928_);
  or (_21188_, _21187_, _02522_);
  or (_21189_, _21188_, _21185_);
  and (_21190_, _08823_, _19621_);
  nand (_21191_, _05617_, _02522_);
  and (_21192_, _21191_, _21190_);
  and (_21193_, _21192_, _21189_);
  or (_21194_, _21011_, _08166_);
  nand (_21195_, _09067_, _08166_);
  and (_21196_, _21195_, _09419_);
  and (_21198_, _21196_, _21194_);
  not (_21199_, _08822_);
  nor (_21200_, _20996_, _08823_);
  or (_21201_, _21200_, _21199_);
  or (_21202_, _21201_, _21198_);
  or (_21203_, _21202_, _21193_);
  or (_21204_, _09066_, _08822_);
  and (_21205_, _21204_, _07139_);
  and (_21206_, _21205_, _21203_);
  and (_21207_, _08882_, _03051_);
  or (_21209_, _21207_, _03148_);
  or (_21210_, _21209_, _21206_);
  nand (_21211_, _09067_, _03148_);
  and (_21212_, _21211_, _21210_);
  or (_21213_, _21212_, _02524_);
  and (_21214_, _09453_, _09446_);
  nand (_21215_, _05617_, _02524_);
  and (_21216_, _21215_, _21214_);
  and (_21217_, _21216_, _21213_);
  or (_21218_, _21011_, _09447_);
  or (_21220_, _09066_, _08166_);
  and (_21221_, _21220_, _09441_);
  and (_21222_, _21221_, _21218_);
  nor (_21223_, _20996_, _09453_);
  or (_21224_, _21223_, _09456_);
  or (_21225_, _21224_, _21222_);
  or (_21226_, _21225_, _21217_);
  or (_21227_, _09066_, _09455_);
  and (_21228_, _21227_, _03023_);
  and (_21229_, _21228_, _21226_);
  and (_21231_, _08882_, _03022_);
  or (_21232_, _21231_, _03137_);
  or (_21233_, _21232_, _21229_);
  nand (_21234_, _09067_, _03137_);
  and (_21235_, _21234_, _21233_);
  or (_21236_, _21235_, _02530_);
  nand (_21237_, _05617_, _02530_);
  and (_21238_, _21237_, _09470_);
  and (_21239_, _21238_, _21236_);
  or (_21240_, _21011_, \oc8051_golden_model_1.PSW [7]);
  or (_21242_, _09066_, _07288_);
  and (_21243_, _21242_, _08818_);
  and (_21244_, _21243_, _21240_);
  or (_21245_, _21244_, _21239_);
  and (_21246_, _21245_, _08815_);
  nor (_21247_, _20996_, _08815_);
  or (_21248_, _21247_, _13433_);
  or (_21249_, _21248_, _21246_);
  or (_21250_, _09066_, _08812_);
  and (_21251_, _21250_, _03043_);
  and (_21253_, _21251_, _21249_);
  and (_21254_, _08882_, _03042_);
  or (_21255_, _21254_, _03143_);
  or (_21256_, _21255_, _21253_);
  nand (_21257_, _09067_, _03143_);
  and (_21258_, _21257_, _21256_);
  or (_21259_, _21258_, _02533_);
  and (_21260_, _19607_, _08806_);
  nand (_21261_, _05617_, _02533_);
  and (_21262_, _21261_, _21260_);
  and (_21264_, _21262_, _21259_);
  or (_21265_, _21011_, _07288_);
  or (_21266_, _09066_, \oc8051_golden_model_1.PSW [7]);
  and (_21267_, _21266_, _08808_);
  and (_21268_, _21267_, _21265_);
  nor (_21269_, _20996_, _08806_);
  or (_21270_, _21269_, _07966_);
  or (_21271_, _21270_, _21268_);
  or (_21272_, _21271_, _21264_);
  or (_21273_, _09066_, _07965_);
  and (_21275_, _21273_, _07996_);
  and (_21276_, _21275_, _21272_);
  and (_21277_, _20994_, _07995_);
  or (_21278_, _21277_, _03155_);
  or (_21279_, _21278_, _21276_);
  or (_21280_, _06171_, _20557_);
  and (_21281_, _21280_, _21279_);
  or (_21282_, _21281_, _02528_);
  nand (_21283_, _05617_, _02528_);
  and (_21284_, _21283_, _03223_);
  and (_21286_, _21284_, _21282_);
  nor (_21287_, _09692_, _08883_);
  and (_21288_, _21003_, _09692_);
  or (_21289_, _21288_, _21287_);
  and (_21290_, _21289_, _03040_);
  or (_21291_, _21290_, _21286_);
  and (_21292_, _21291_, _08803_);
  not (_21293_, _03358_);
  and (_21294_, _07189_, _21293_);
  nor (_21295_, _20994_, _08112_);
  nor (_21297_, _21295_, _21294_);
  or (_21298_, _21297_, _21292_);
  nand (_21299_, _09067_, _08112_);
  and (_21300_, _21299_, _08116_);
  and (_21301_, _21300_, _21298_);
  and (_21302_, _20994_, _08115_);
  or (_21303_, _21302_, _02890_);
  or (_21304_, _21303_, _21301_);
  or (_21305_, _06171_, _02891_);
  and (_21306_, _21305_, _08788_);
  and (_21308_, _21306_, _21304_);
  nor (_21309_, _05617_, _08788_);
  or (_21310_, _21309_, _02889_);
  or (_21311_, _21310_, _21308_);
  and (_21312_, _09692_, _08883_);
  nor (_21313_, _21003_, _09692_);
  nor (_21314_, _21313_, _21312_);
  or (_21315_, _21314_, _03175_);
  and (_21316_, _21315_, _09724_);
  and (_21317_, _21316_, _21311_);
  nor (_21319_, _20996_, _09724_);
  or (_21320_, _21319_, _03174_);
  or (_21321_, _21320_, _21317_);
  nand (_21322_, _09067_, _03174_);
  and (_21323_, _21322_, _09732_);
  and (_21324_, _21323_, _21321_);
  nor (_21325_, _20996_, _09732_);
  or (_21326_, _21325_, _04150_);
  or (_21327_, _21326_, _21324_);
  nand (_21328_, _05617_, _04150_);
  and (_21330_, _21328_, _03183_);
  and (_21331_, _21330_, _21327_);
  and (_21332_, _21314_, _02799_);
  nor (_21333_, _21332_, _21331_);
  or (_21334_, _21333_, _09748_);
  or (_21335_, _20996_, _09747_);
  and (_21336_, _21335_, _02888_);
  and (_21337_, _21336_, _21334_);
  and (_21338_, _09067_, _02887_);
  nor (_21339_, _21338_, _09756_);
  not (_21341_, _21339_);
  nor (_21342_, _21341_, _21337_);
  or (_21343_, _21342_, _19863_);
  nor (_21344_, _21343_, _20997_);
  and (_21345_, _19863_, _05617_);
  nor (_21346_, _21345_, _08786_);
  not (_21347_, _21346_);
  nor (_21348_, _21347_, _21344_);
  nor (_21349_, _21348_, _20995_);
  nand (_21350_, _21349_, _34655_);
  or (_21352_, _34655_, \oc8051_golden_model_1.PC [4]);
  and (_21353_, _21352_, _35796_);
  and (_35842_[4], _21353_, _21350_);
  nor (_21354_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_21355_, _09061_, _02247_);
  nor (_21356_, _21355_, _21354_);
  and (_21357_, _21356_, _08786_);
  nor (_21358_, _21356_, _09755_);
  and (_21359_, _09061_, _03174_);
  and (_21360_, _06083_, _02890_);
  nor (_21362_, _21356_, _08803_);
  nor (_21363_, _21356_, _08806_);
  nor (_21364_, _21356_, _08815_);
  nor (_21365_, _21356_, _09453_);
  nor (_21366_, _21356_, _08823_);
  not (_21367_, _21356_);
  and (_21368_, _21367_, _09249_);
  and (_21369_, _09297_, _08877_);
  or (_21370_, _08880_, _08879_);
  not (_21371_, _21370_);
  nor (_21374_, _21371_, _08912_);
  and (_21375_, _21371_, _08912_);
  nor (_21376_, _21375_, _21374_);
  nor (_21377_, _21376_, _09297_);
  nor (_21378_, _21377_, _21369_);
  or (_21379_, _21378_, _09299_);
  not (_21380_, _21376_);
  and (_21381_, _21380_, _08981_);
  and (_21382_, _09918_, _08877_);
  or (_21383_, _21382_, _21381_);
  nor (_21386_, _21383_, _08986_);
  or (_21387_, _21380_, _09003_);
  nand (_21388_, _09003_, _08878_);
  and (_21389_, _21388_, _21387_);
  or (_21390_, _21389_, _03006_);
  or (_21391_, _09063_, _09064_);
  and (_21392_, _21391_, _09089_);
  nor (_21393_, _21391_, _09089_);
  nor (_21394_, _21393_, _21392_);
  and (_21395_, _21394_, _19652_);
  and (_21398_, _19659_, _09061_);
  nor (_21399_, _21398_, _21395_);
  nand (_21400_, _21399_, _09132_);
  nor (_21401_, _05649_, _02601_);
  and (_21402_, _09061_, _02951_);
  nor (_21403_, _05649_, _02603_);
  not (_21404_, _09135_);
  and (_21405_, _09061_, _03845_);
  nor (_21406_, _21405_, _21404_);
  nor (_21407_, _09138_, \oc8051_golden_model_1.PC [5]);
  nor (_21410_, _21407_, _03845_);
  not (_21411_, _21410_);
  and (_21412_, _21411_, _21406_);
  not (_21413_, _21412_);
  nor (_21414_, _21356_, _09145_);
  nor (_21415_, _21414_, _03849_);
  and (_21416_, _21415_, _21413_);
  nor (_21417_, _21416_, _09154_);
  not (_21418_, _21417_);
  nor (_21419_, _21418_, _21403_);
  nor (_21422_, _21356_, _09153_);
  nor (_21423_, _21422_, _02951_);
  not (_21424_, _21423_);
  nor (_21425_, _21424_, _21419_);
  or (_21426_, _21425_, _07436_);
  nor (_21427_, _21426_, _21402_);
  and (_21428_, _21367_, _07436_);
  nor (_21429_, _21428_, _09169_);
  not (_21430_, _21429_);
  nor (_21431_, _21430_, _21427_);
  nor (_21434_, _21431_, _21401_);
  nor (_21435_, _21434_, _07433_);
  and (_21436_, _21356_, _07433_);
  nor (_21437_, _21436_, _09132_);
  not (_21438_, _21437_);
  nor (_21439_, _21438_, _21435_);
  nor (_21440_, _21439_, _03840_);
  and (_21441_, _21440_, _21400_);
  and (_21442_, _21356_, _03840_);
  or (_21443_, _21442_, _02948_);
  or (_21445_, _21443_, _21441_);
  nand (_21446_, _21445_, _21390_);
  nand (_21447_, _21446_, _08997_);
  nor (_21448_, _21356_, _08997_);
  nor (_21449_, _21448_, _02884_);
  nand (_21450_, _21449_, _21447_);
  and (_21451_, _09061_, _02884_);
  nor (_21452_, _21451_, _04225_);
  nand (_21453_, _21452_, _21450_);
  and (_21454_, _05649_, _04225_);
  nor (_21456_, _21454_, _02946_);
  nand (_21457_, _21456_, _21453_);
  and (_21458_, _09061_, _02946_);
  nor (_21459_, _21458_, _09187_);
  nand (_21460_, _21459_, _21457_);
  nor (_21461_, _21356_, _09186_);
  nor (_21462_, _21461_, _02880_);
  nand (_21463_, _21462_, _21460_);
  and (_21464_, _09061_, _02880_);
  nor (_21465_, _21464_, _09193_);
  nand (_21467_, _21465_, _21463_);
  and (_21468_, _21367_, _09193_);
  nor (_21469_, _21468_, _02877_);
  and (_21470_, _21469_, _21467_);
  and (_21471_, _09061_, _02877_);
  or (_21472_, _21471_, _08989_);
  or (_21473_, _21472_, _21470_);
  and (_21474_, _05649_, _08989_);
  nor (_21475_, _21474_, _02876_);
  nand (_21476_, _21475_, _21473_);
  and (_21478_, _09061_, _02876_);
  nor (_21479_, _21478_, _09210_);
  nand (_21480_, _21479_, _21476_);
  and (_21481_, _09242_, _08877_);
  nor (_21482_, _21376_, _09242_);
  or (_21483_, _21482_, _09209_);
  or (_21484_, _21483_, _21481_);
  nand (_21485_, _21484_, _21480_);
  and (_21486_, _21485_, _08986_);
  or (_21487_, _21486_, _21386_);
  or (_21489_, _21487_, _02954_);
  and (_21490_, _21489_, _21379_);
  or (_21491_, _21490_, _03029_);
  and (_21492_, _09276_, _08877_);
  nor (_21493_, _21376_, _09276_);
  or (_21494_, _21493_, _21492_);
  and (_21495_, _21494_, _03029_);
  nor (_21496_, _21495_, _09249_);
  and (_21497_, _21496_, _21491_);
  or (_21498_, _21497_, _21368_);
  nand (_21500_, _21498_, _06246_);
  and (_21501_, _09062_, _02871_);
  nor (_21502_, _21501_, _09257_);
  nand (_21503_, _21502_, _21500_);
  nor (_21504_, _05649_, _02591_);
  nor (_21505_, _21504_, _20030_);
  and (_21506_, _21505_, _21503_);
  nor (_21507_, _09262_, _09061_);
  or (_21508_, _21507_, _21506_);
  nand (_21509_, _21508_, _09309_);
  nor (_21511_, _21356_, _09309_);
  nor (_21512_, _21511_, _02941_);
  nand (_21513_, _21512_, _21509_);
  and (_21514_, _09061_, _02941_);
  nor (_21515_, _21514_, _19627_);
  nand (_21516_, _21515_, _21513_);
  and (_21517_, _05649_, _19627_);
  nor (_21518_, _21517_, _02940_);
  nand (_21519_, _21518_, _21516_);
  and (_21520_, _09061_, _02940_);
  nor (_21522_, _21520_, _09326_);
  and (_21523_, _21522_, _21519_);
  nor (_21524_, _21356_, _09320_);
  or (_21525_, _21524_, _21523_);
  nand (_21526_, _21525_, _09324_);
  nor (_21527_, _09324_, _09061_);
  nor (_21528_, _21527_, _07721_);
  and (_21529_, _21528_, _21526_);
  nor (_21530_, _21367_, _02571_);
  or (_21531_, _21530_, _02866_);
  nor (_21533_, _21531_, _21529_);
  and (_21534_, _09062_, _02866_);
  or (_21535_, _21534_, _21533_);
  nand (_21536_, _21535_, _04134_);
  and (_21537_, _05649_, _02569_);
  nor (_21538_, _21537_, _03046_);
  nand (_21539_, _21538_, _21536_);
  and (_21540_, _08877_, _03046_);
  not (_21541_, _21540_);
  and (_21542_, _21541_, _02860_);
  nand (_21544_, _21542_, _21539_);
  nor (_21545_, _09061_, _02860_);
  nor (_21546_, _21545_, _02567_);
  and (_21547_, _21546_, _21544_);
  nor (_21548_, _09352_, _08877_);
  nor (_21549_, _21548_, _09353_);
  or (_21550_, _21549_, _21547_);
  and (_21551_, _21367_, _09352_);
  nor (_21552_, _21551_, _02930_);
  nand (_21553_, _21552_, _21550_);
  and (_21555_, _09061_, _02930_);
  nor (_21556_, _21555_, _02516_);
  nand (_21557_, _21556_, _21553_);
  and (_21558_, _05649_, _02516_);
  nor (_21559_, _21558_, _09362_);
  nand (_21560_, _21559_, _21557_);
  and (_21561_, _21394_, _09362_);
  nor (_21562_, _21561_, _05749_);
  nand (_21563_, _21562_, _21560_);
  nor (_21564_, _09061_, _05748_);
  nor (_21566_, _21564_, _02834_);
  and (_21567_, _21566_, _21563_);
  and (_21568_, _08877_, _02834_);
  or (_21569_, _21568_, _07830_);
  nor (_21570_, _21569_, _21567_);
  and (_21571_, _09062_, _07830_);
  or (_21572_, _21571_, _21570_);
  nand (_21573_, _21572_, _19622_);
  and (_21574_, _09397_, _09390_);
  nor (_21575_, _21574_, _09398_);
  nor (_21577_, _21575_, _19622_);
  nor (_21578_, _21577_, _02928_);
  nand (_21579_, _21578_, _21573_);
  and (_21580_, _09061_, _02928_);
  nor (_21581_, _21580_, _02522_);
  nand (_21582_, _21581_, _21579_);
  and (_21583_, _05649_, _02522_);
  nor (_21584_, _21583_, _09419_);
  nand (_21585_, _21584_, _21582_);
  and (_21586_, _09061_, _08166_);
  and (_21588_, _21394_, _09447_);
  or (_21589_, _21588_, _21586_);
  and (_21590_, _21589_, _09419_);
  nor (_21591_, _21590_, _09428_);
  and (_21592_, _21591_, _21585_);
  or (_21593_, _21592_, _21366_);
  nand (_21594_, _21593_, _08822_);
  nor (_21595_, _09061_, _08822_);
  nor (_21596_, _21595_, _03051_);
  and (_21597_, _21596_, _21594_);
  and (_21599_, _08877_, _03051_);
  or (_21600_, _21599_, _03148_);
  nor (_21601_, _21600_, _21597_);
  and (_21602_, _09062_, _03148_);
  or (_21603_, _21602_, _21601_);
  nand (_21604_, _21603_, _19618_);
  and (_21605_, _05649_, _02524_);
  nor (_21606_, _21605_, _09441_);
  nand (_21607_, _21606_, _21604_);
  nor (_21608_, _21394_, _09447_);
  nor (_21610_, _09061_, _08166_);
  nor (_21611_, _21610_, _09446_);
  not (_21612_, _21611_);
  nor (_21613_, _21612_, _21608_);
  nor (_21614_, _21613_, _20129_);
  and (_21615_, _21614_, _21607_);
  or (_21616_, _21615_, _21365_);
  nand (_21617_, _21616_, _09455_);
  nor (_21618_, _09061_, _09455_);
  nor (_21619_, _21618_, _03022_);
  and (_21621_, _21619_, _21617_);
  and (_21622_, _08877_, _03022_);
  or (_21623_, _21622_, _03137_);
  nor (_21624_, _21623_, _21621_);
  and (_21625_, _09062_, _03137_);
  or (_21626_, _21625_, _21624_);
  nand (_21627_, _21626_, _19615_);
  and (_21628_, _05649_, _02530_);
  nor (_21629_, _21628_, _08818_);
  nand (_21630_, _21629_, _21627_);
  nor (_21632_, _21394_, \oc8051_golden_model_1.PSW [7]);
  nor (_21633_, _09061_, _07288_);
  nor (_21634_, _21633_, _09470_);
  not (_21635_, _21634_);
  nor (_21636_, _21635_, _21632_);
  nor (_21637_, _21636_, _09468_);
  and (_21638_, _21637_, _21630_);
  or (_21639_, _21638_, _21364_);
  nand (_21640_, _21639_, _08812_);
  nor (_21641_, _09061_, _08812_);
  nor (_21643_, _21641_, _03042_);
  and (_21644_, _21643_, _21640_);
  and (_21645_, _08877_, _03042_);
  or (_21646_, _21645_, _03143_);
  nor (_21647_, _21646_, _21644_);
  and (_21648_, _09062_, _03143_);
  or (_21649_, _21648_, _21647_);
  nand (_21650_, _21649_, _02534_);
  and (_21651_, _05649_, _02533_);
  nor (_21652_, _21651_, _08808_);
  nand (_21654_, _21652_, _21650_);
  or (_21655_, _21394_, _07288_);
  or (_21656_, _09061_, \oc8051_golden_model_1.PSW [7]);
  and (_21657_, _21656_, _08808_);
  and (_21658_, _21657_, _21655_);
  nor (_21659_, _21658_, _09487_);
  and (_21660_, _21659_, _21654_);
  or (_21661_, _21660_, _21363_);
  nand (_21662_, _21661_, _07965_);
  nor (_21663_, _09061_, _07965_);
  nor (_21665_, _21663_, _07995_);
  and (_21666_, _21665_, _21662_);
  and (_21667_, _21356_, _07995_);
  or (_21668_, _21667_, _03155_);
  nor (_21669_, _21668_, _21666_);
  and (_21670_, _06083_, _03155_);
  or (_21671_, _21670_, _21669_);
  nand (_21672_, _21671_, _05790_);
  and (_21673_, _05649_, _02528_);
  nor (_21674_, _21673_, _03040_);
  nand (_21676_, _21674_, _21672_);
  nor (_21677_, _09692_, _08877_);
  and (_21678_, _21376_, _09692_);
  or (_21679_, _21678_, _03223_);
  or (_21680_, _21679_, _21677_);
  and (_21681_, _21680_, _08803_);
  and (_21682_, _21681_, _21676_);
  or (_21683_, _21682_, _21362_);
  nand (_21684_, _21683_, _08789_);
  and (_21685_, _09062_, _08112_);
  nor (_21687_, _21685_, _08115_);
  nand (_21688_, _21687_, _21684_);
  and (_21689_, _21356_, _08115_);
  nor (_21690_, _21689_, _02890_);
  and (_21691_, _21690_, _21688_);
  or (_21692_, _21691_, _21360_);
  nand (_21693_, _21692_, _08788_);
  and (_21694_, _05649_, _02510_);
  nor (_21695_, _21694_, _02889_);
  nand (_21696_, _21695_, _21693_);
  nor (_21698_, _21380_, _09692_);
  and (_21699_, _09692_, _08878_);
  nor (_21700_, _21699_, _21698_);
  and (_21701_, _21700_, _02889_);
  nor (_21702_, _21701_, _09725_);
  nand (_21703_, _21702_, _21696_);
  nor (_21704_, _21356_, _09724_);
  nor (_21705_, _21704_, _03174_);
  and (_21706_, _21705_, _21703_);
  or (_21707_, _21706_, _21359_);
  nand (_21709_, _21707_, _09732_);
  nor (_21710_, _21367_, _09732_);
  nor (_21711_, _21710_, _04150_);
  nand (_21712_, _21711_, _21709_);
  and (_21713_, _05649_, _04150_);
  nor (_21714_, _21713_, _02799_);
  nand (_21715_, _21714_, _21712_);
  and (_21716_, _21700_, _02799_);
  nor (_21717_, _21716_, _09748_);
  nand (_21718_, _21717_, _21715_);
  nor (_21720_, _21356_, _09747_);
  nor (_21721_, _21720_, _02887_);
  nand (_21722_, _21721_, _21718_);
  and (_21723_, _09061_, _02887_);
  nor (_21724_, _21723_, _09756_);
  and (_21725_, _21724_, _21722_);
  or (_21726_, _21725_, _21358_);
  nand (_21727_, _21726_, _19862_);
  and (_21728_, _19863_, _05649_);
  nor (_21729_, _21728_, _08786_);
  and (_21731_, _21729_, _21727_);
  or (_21732_, _21731_, _21357_);
  or (_21733_, _21732_, _34659_);
  or (_21734_, _34655_, \oc8051_golden_model_1.PC [5]);
  and (_21735_, _21734_, _35796_);
  and (_35842_[5], _21735_, _21733_);
  and (_21736_, _05264_, _08790_);
  nor (_21737_, _21736_, \oc8051_golden_model_1.PC [6]);
  nor (_21738_, _21737_, _08791_);
  and (_21739_, _21738_, _08786_);
  not (_21741_, _21738_);
  nor (_21742_, _21741_, _09755_);
  and (_21743_, _09055_, _02887_);
  or (_21744_, _21743_, _09756_);
  and (_21745_, _05585_, _04150_);
  and (_21746_, _21741_, _08115_);
  and (_21747_, _09470_, _08815_);
  and (_21748_, _08869_, _03051_);
  nor (_21749_, _21738_, _02571_);
  and (_21750_, _21741_, _09249_);
  and (_21752_, _09055_, _02877_);
  and (_21753_, _21741_, _09181_);
  and (_21754_, _05585_, _03849_);
  nand (_21755_, _09055_, _03845_);
  nand (_21756_, _21755_, _09135_);
  not (_21757_, \oc8051_golden_model_1.PC [6]);
  or (_21758_, _09138_, _21757_);
  and (_21759_, _21758_, _04194_);
  or (_21760_, _21759_, _21756_);
  or (_21761_, _21741_, _09145_);
  and (_21763_, _21761_, _02603_);
  and (_21764_, _21763_, _21760_);
  or (_21765_, _21764_, _09154_);
  or (_21766_, _21765_, _21754_);
  or (_21767_, _21741_, _09153_);
  and (_21768_, _21767_, _03401_);
  and (_21769_, _21768_, _21766_);
  and (_21770_, _09055_, _02951_);
  or (_21771_, _21770_, _21769_);
  and (_21772_, _21771_, _19632_);
  and (_21774_, _21741_, _07436_);
  or (_21775_, _21774_, _21772_);
  and (_21776_, _21775_, _02601_);
  and (_21777_, _05585_, _09169_);
  or (_21778_, _21777_, _07433_);
  or (_21779_, _21778_, _21776_);
  nand (_21780_, _21738_, _07433_);
  and (_21781_, _21780_, _05361_);
  and (_21782_, _21781_, _21779_);
  nor (_21783_, _09091_, _09058_);
  or (_21785_, _21783_, _09092_);
  or (_21786_, _21785_, _09012_);
  or (_21787_, _19652_, _09055_);
  and (_21788_, _21787_, _09132_);
  and (_21789_, _21788_, _21786_);
  or (_21790_, _21789_, _21782_);
  and (_21791_, _21790_, _09176_);
  and (_21792_, _08914_, _08874_);
  or (_21793_, _21792_, _08915_);
  or (_21794_, _21793_, _09003_);
  nand (_21796_, _09003_, _08868_);
  and (_21797_, _21796_, _02948_);
  and (_21798_, _21797_, _21794_);
  or (_21799_, _21798_, _21791_);
  and (_21800_, _21799_, _08997_);
  or (_21801_, _21800_, _21753_);
  and (_21802_, _21801_, _02934_);
  and (_21803_, _09055_, _02884_);
  or (_21804_, _21803_, _04225_);
  or (_21805_, _21804_, _21802_);
  or (_21807_, _05585_, _02597_);
  and (_21808_, _21807_, _07474_);
  and (_21809_, _21808_, _21805_);
  and (_21810_, _09055_, _02946_);
  or (_21811_, _21810_, _21809_);
  and (_21812_, _21811_, _09186_);
  nor (_21813_, _21738_, _09186_);
  or (_21814_, _21813_, _21812_);
  and (_21815_, _21814_, _02992_);
  and (_21816_, _09055_, _02880_);
  or (_21818_, _21816_, _09193_);
  or (_21819_, _21818_, _21815_);
  nand (_21820_, _21738_, _09193_);
  and (_21821_, _21820_, _02987_);
  and (_21822_, _21821_, _21819_);
  or (_21823_, _21822_, _21752_);
  and (_21824_, _21823_, _02595_);
  and (_21825_, _05585_, _08989_);
  or (_21826_, _21825_, _02876_);
  or (_21827_, _21826_, _21824_);
  nand (_21829_, _09054_, _02876_);
  and (_21830_, _21829_, _09209_);
  and (_21831_, _21830_, _21827_);
  nand (_21832_, _09242_, _08868_);
  or (_21833_, _21793_, _09242_);
  and (_21834_, _21833_, _21832_);
  and (_21835_, _21834_, _09210_);
  or (_21836_, _21835_, _21831_);
  and (_21837_, _21836_, _08986_);
  nand (_21838_, _09918_, _08868_);
  or (_21840_, _21793_, _09918_);
  and (_21841_, _21840_, _08985_);
  and (_21842_, _21841_, _21838_);
  or (_21843_, _21842_, _02954_);
  or (_21844_, _21843_, _21837_);
  nand (_21845_, _09297_, _08868_);
  or (_21846_, _21793_, _09297_);
  and (_21847_, _21846_, _21845_);
  or (_21848_, _21847_, _09299_);
  and (_21849_, _21848_, _21844_);
  or (_21851_, _21849_, _03029_);
  and (_21852_, _21793_, _09277_);
  and (_21853_, _09276_, _08869_);
  or (_21854_, _21853_, _09279_);
  or (_21855_, _21854_, _21852_);
  and (_21856_, _21855_, _09250_);
  and (_21857_, _21856_, _21851_);
  or (_21858_, _21857_, _21750_);
  and (_21859_, _21858_, _06246_);
  and (_21860_, _09055_, _02871_);
  or (_21862_, _21860_, _09257_);
  or (_21863_, _21862_, _21859_);
  or (_21864_, _05585_, _02591_);
  and (_21865_, _21864_, _09262_);
  and (_21866_, _21865_, _21863_);
  nor (_21867_, _09262_, _09054_);
  or (_21868_, _21867_, _21866_);
  and (_21869_, _21868_, _09309_);
  nor (_21870_, _21738_, _09309_);
  or (_21871_, _21870_, _02941_);
  or (_21873_, _21871_, _21869_);
  nand (_21874_, _09054_, _02941_);
  and (_21875_, _21874_, _02589_);
  and (_21876_, _21875_, _21873_);
  and (_21877_, _05585_, _19627_);
  or (_21878_, _21877_, _02940_);
  or (_21879_, _21878_, _21876_);
  nand (_21880_, _09054_, _02940_);
  and (_21881_, _21880_, _09320_);
  and (_21882_, _21881_, _21879_);
  nor (_21884_, _21738_, _09320_);
  or (_21885_, _21884_, _09325_);
  or (_21886_, _21885_, _21882_);
  or (_21887_, _09324_, _09055_);
  and (_21888_, _21887_, _02571_);
  and (_21889_, _21888_, _21886_);
  or (_21890_, _21889_, _21749_);
  and (_21891_, _21890_, _02986_);
  and (_21892_, _09055_, _02866_);
  or (_21893_, _21892_, _02569_);
  or (_21895_, _21893_, _21891_);
  or (_21896_, _05585_, _04134_);
  and (_21897_, _21896_, _08211_);
  and (_21898_, _21897_, _21895_);
  nand (_21899_, _08869_, _03046_);
  nand (_21900_, _21899_, _02860_);
  or (_21901_, _21900_, _21898_);
  or (_21902_, _09055_, _02860_);
  and (_21903_, _21902_, _02839_);
  and (_21904_, _21903_, _21901_);
  nor (_21906_, _09352_, _08869_);
  nor (_21907_, _21906_, _09353_);
  or (_21908_, _21907_, _21904_);
  nand (_21909_, _21738_, _09352_);
  and (_21910_, _21909_, _03508_);
  and (_21911_, _21910_, _21908_);
  and (_21912_, _09055_, _02930_);
  or (_21913_, _21912_, _21911_);
  and (_21914_, _21913_, _02517_);
  and (_21915_, _05585_, _02516_);
  or (_21917_, _21915_, _09362_);
  or (_21918_, _21917_, _21914_);
  or (_21919_, _21785_, _09366_);
  and (_21920_, _21919_, _05748_);
  and (_21921_, _21920_, _21918_);
  nor (_21922_, _09054_, _05748_);
  or (_21923_, _21922_, _21921_);
  and (_21924_, _21923_, _07140_);
  and (_21925_, _08869_, _02834_);
  or (_21926_, _21925_, _07830_);
  or (_21928_, _21926_, _21924_);
  nand (_21929_, _09054_, _07830_);
  and (_21930_, _21929_, _19622_);
  and (_21931_, _21930_, _21928_);
  and (_21932_, _09399_, _09386_);
  or (_21933_, _21932_, _09400_);
  and (_21934_, _21933_, _09376_);
  or (_21935_, _21934_, _02928_);
  or (_21936_, _21935_, _21931_);
  nand (_21937_, _09054_, _02928_);
  and (_21938_, _21937_, _04131_);
  and (_21939_, _21938_, _21936_);
  and (_21940_, _05585_, _02522_);
  or (_21941_, _21940_, _09419_);
  or (_21942_, _21941_, _21939_);
  and (_21943_, _21785_, _09447_);
  or (_21944_, _09054_, _09447_);
  nand (_21945_, _21944_, _09419_);
  or (_21946_, _21945_, _21943_);
  and (_21947_, _21946_, _08823_);
  and (_21950_, _21947_, _21942_);
  nor (_21951_, _21738_, _08823_);
  or (_21952_, _21951_, _21199_);
  or (_21953_, _21952_, _21950_);
  or (_21954_, _09055_, _08822_);
  and (_21955_, _21954_, _07139_);
  and (_21956_, _21955_, _21953_);
  or (_21957_, _21956_, _21748_);
  and (_21958_, _21957_, _07150_);
  and (_21959_, _09055_, _03148_);
  or (_21961_, _21959_, _02524_);
  or (_21962_, _21961_, _21958_);
  or (_21963_, _05585_, _19618_);
  nand (_21964_, _21963_, _21962_);
  nand (_21965_, _21964_, _21214_);
  or (_21966_, _21741_, _09453_);
  and (_21967_, _21785_, _08166_);
  or (_21968_, _09054_, _08166_);
  nand (_21969_, _21968_, _09441_);
  or (_21970_, _21969_, _21967_);
  and (_21972_, _21970_, _21966_);
  and (_21973_, _21972_, _21965_);
  or (_21974_, _21973_, _09456_);
  or (_21975_, _09055_, _09455_);
  and (_21976_, _21975_, _21974_);
  or (_21977_, _21976_, _03022_);
  nand (_21978_, _08868_, _03022_);
  and (_21979_, _21978_, _06213_);
  and (_21980_, _21979_, _21977_);
  and (_21981_, _09055_, _03137_);
  or (_21983_, _21981_, _02530_);
  or (_21984_, _21983_, _21980_);
  or (_21985_, _05585_, _19615_);
  nand (_21986_, _21985_, _21984_);
  nand (_21987_, _21986_, _21747_);
  or (_21988_, _21741_, _08815_);
  and (_21989_, _21785_, _07288_);
  or (_21990_, _09054_, _07288_);
  nand (_21991_, _21990_, _08818_);
  or (_21992_, _21991_, _21989_);
  and (_21994_, _21992_, _21988_);
  and (_21995_, _21994_, _21987_);
  or (_21996_, _21995_, _13433_);
  or (_21997_, _09055_, _08812_);
  and (_21998_, _21997_, _03043_);
  and (_21999_, _21998_, _21996_);
  and (_22000_, _08869_, _03042_);
  or (_22001_, _22000_, _03143_);
  or (_22002_, _22001_, _21999_);
  nand (_22003_, _09054_, _03143_);
  and (_22005_, _22003_, _02534_);
  and (_22006_, _22005_, _22002_);
  and (_22007_, _05585_, _02533_);
  nor (_22008_, _22007_, _22006_);
  nand (_22009_, _22008_, _21260_);
  or (_22010_, _21741_, _08806_);
  and (_22011_, _21785_, \oc8051_golden_model_1.PSW [7]);
  or (_22012_, _09054_, \oc8051_golden_model_1.PSW [7]);
  nand (_22013_, _22012_, _08808_);
  or (_22014_, _22013_, _22011_);
  and (_22016_, _22014_, _22010_);
  and (_22017_, _22016_, _22009_);
  or (_22018_, _22017_, _07966_);
  or (_22019_, _09055_, _07965_);
  and (_22020_, _22019_, _22018_);
  or (_22021_, _22020_, _07995_);
  nand (_22022_, _21738_, _07995_);
  and (_22023_, _22022_, _20557_);
  and (_22024_, _22023_, _22021_);
  and (_22025_, _05855_, _03155_);
  or (_22027_, _22025_, _22024_);
  and (_22028_, _22027_, _05790_);
  and (_22029_, _05585_, _02528_);
  or (_22030_, _22029_, _03040_);
  or (_22031_, _22030_, _22028_);
  nor (_22032_, _09692_, _08868_);
  and (_22033_, _21793_, _09692_);
  or (_22034_, _22033_, _03223_);
  or (_22035_, _22034_, _22032_);
  and (_22036_, _22035_, _08803_);
  and (_22038_, _22036_, _22031_);
  nor (_22039_, _21741_, _08112_);
  nor (_22040_, _22039_, _21294_);
  or (_22041_, _22040_, _22038_);
  nand (_22042_, _09054_, _08112_);
  and (_22043_, _22042_, _08116_);
  and (_22044_, _22043_, _22041_);
  or (_22045_, _22044_, _21746_);
  and (_22046_, _22045_, _02891_);
  and (_22047_, _05855_, _02890_);
  or (_22049_, _22047_, _02510_);
  or (_22050_, _22049_, _22046_);
  or (_22051_, _05585_, _08788_);
  and (_22052_, _22051_, _03175_);
  and (_22053_, _22052_, _22050_);
  nand (_22054_, _09692_, _08868_);
  or (_22055_, _21793_, _09692_);
  and (_22056_, _22055_, _22054_);
  and (_22057_, _22056_, _02889_);
  or (_22058_, _22057_, _22053_);
  and (_22060_, _22058_, _09724_);
  nor (_22061_, _21738_, _09724_);
  or (_22062_, _22061_, _22060_);
  and (_22063_, _22062_, _03179_);
  nand (_22064_, _09055_, _03174_);
  nand (_22065_, _22064_, _09732_);
  or (_22066_, _22065_, _22063_);
  or (_22067_, _21741_, _09732_);
  and (_22068_, _22067_, _03936_);
  and (_22069_, _22068_, _22066_);
  or (_22071_, _22069_, _21745_);
  and (_22072_, _22071_, _03183_);
  and (_22073_, _22056_, _02799_);
  or (_22074_, _22073_, _09748_);
  nor (_22075_, _22074_, _22072_);
  nor (_22076_, _21741_, _09747_);
  nor (_22077_, _22076_, _02887_);
  not (_22078_, _22077_);
  nor (_22079_, _22078_, _22075_);
  nor (_22080_, _22079_, _21744_);
  or (_22082_, _22080_, _19863_);
  nor (_22083_, _22082_, _21742_);
  and (_22084_, _19863_, _05585_);
  or (_22085_, _22084_, _08786_);
  nor (_22086_, _22085_, _22083_);
  or (_22087_, _22086_, _21739_);
  or (_22088_, _22087_, _34659_);
  or (_22089_, _34655_, \oc8051_golden_model_1.PC [6]);
  and (_22090_, _22089_, _35796_);
  and (_35842_[6], _22090_, _22088_);
  nor (_22092_, _08791_, \oc8051_golden_model_1.PC [7]);
  nor (_22093_, _22092_, _08792_);
  and (_22094_, _22093_, _08786_);
  and (_22095_, _19863_, _05302_);
  nand (_22096_, _05269_, _03174_);
  nor (_22097_, _22093_, _08803_);
  nor (_22098_, _22093_, _08806_);
  nor (_22099_, _22093_, _08815_);
  nor (_22100_, _22093_, _09453_);
  nor (_22101_, _22093_, _08823_);
  and (_22103_, _05507_, _02866_);
  nor (_22104_, _22093_, _09320_);
  nor (_22105_, _09262_, _05269_);
  not (_22106_, _22093_);
  and (_22107_, _22106_, _09249_);
  nand (_22108_, _09918_, _06146_);
  or (_22109_, _08864_, _08865_);
  and (_22110_, _22109_, _08916_);
  nor (_22111_, _22109_, _08916_);
  nor (_22112_, _22111_, _22110_);
  not (_22114_, _22112_);
  or (_22115_, _22114_, _09918_);
  and (_22116_, _22115_, _22108_);
  and (_22117_, _22116_, _08985_);
  and (_22118_, _09003_, _06147_);
  nor (_22119_, _22112_, _09003_);
  or (_22120_, _22119_, _22118_);
  and (_22121_, _22120_, _02948_);
  and (_22122_, _09093_, _09051_);
  nor (_22123_, _22122_, _09094_);
  nand (_22125_, _22123_, _19652_);
  nand (_22126_, _19659_, _05269_);
  and (_22127_, _22126_, _22125_);
  and (_22128_, _22127_, _09132_);
  or (_22129_, _05302_, _02603_);
  nand (_22130_, _05269_, _03845_);
  and (_22131_, _22130_, _09135_);
  nor (_22132_, _09138_, \oc8051_golden_model_1.PC [7]);
  or (_22133_, _22132_, _03845_);
  and (_22134_, _22133_, _22131_);
  nor (_22136_, _22093_, _09145_);
  or (_22137_, _22136_, _03849_);
  or (_22138_, _22137_, _22134_);
  and (_22139_, _22138_, _09153_);
  and (_22140_, _22139_, _22129_);
  nor (_22141_, _22093_, _09153_);
  or (_22142_, _22141_, _02951_);
  or (_22143_, _22142_, _22140_);
  and (_22144_, _05269_, _02951_);
  nor (_22145_, _22144_, _07436_);
  and (_22147_, _22145_, _22143_);
  and (_22148_, _22106_, _07436_);
  or (_22149_, _22148_, _09169_);
  or (_22150_, _22149_, _22147_);
  or (_22151_, _05302_, _02601_);
  and (_22152_, _22151_, _22150_);
  or (_22153_, _22152_, _07433_);
  nand (_22154_, _22093_, _07433_);
  and (_22155_, _22154_, _05361_);
  and (_22156_, _22155_, _22153_);
  or (_22158_, _22156_, _03840_);
  or (_22159_, _22158_, _22128_);
  nand (_22160_, _22093_, _03840_);
  and (_22161_, _22160_, _03006_);
  and (_22162_, _22161_, _22159_);
  or (_22163_, _22162_, _22121_);
  and (_22164_, _22163_, _08997_);
  nor (_22165_, _22093_, _08997_);
  or (_22166_, _22165_, _02884_);
  or (_22167_, _22166_, _22164_);
  nand (_22169_, _05269_, _02884_);
  and (_22170_, _22169_, _02597_);
  and (_22171_, _22170_, _22167_);
  and (_22172_, _05302_, _04225_);
  or (_22173_, _22172_, _02946_);
  or (_22174_, _22173_, _22171_);
  nand (_22175_, _05269_, _02946_);
  and (_22176_, _22175_, _09186_);
  and (_22177_, _22176_, _22174_);
  nor (_22178_, _22093_, _09186_);
  or (_22180_, _22178_, _02880_);
  or (_22181_, _22180_, _22177_);
  and (_22182_, _05269_, _02880_);
  nor (_22183_, _22182_, _09193_);
  and (_22184_, _22183_, _22181_);
  and (_22185_, _22106_, _09193_);
  or (_22186_, _22185_, _02877_);
  or (_22187_, _22186_, _22184_);
  nand (_22188_, _05269_, _02877_);
  and (_22189_, _22188_, _02595_);
  and (_22191_, _22189_, _22187_);
  and (_22192_, _05302_, _08989_);
  or (_22193_, _22192_, _02876_);
  or (_22194_, _22193_, _22191_);
  nand (_22195_, _05269_, _02876_);
  and (_22196_, _22195_, _09209_);
  and (_22197_, _22196_, _22194_);
  nand (_22198_, _09242_, _06146_);
  or (_22199_, _22114_, _09242_);
  and (_22200_, _22199_, _22198_);
  and (_22202_, _22200_, _09210_);
  or (_22203_, _22202_, _22197_);
  and (_22204_, _22203_, _08986_);
  or (_22205_, _22204_, _22117_);
  and (_22206_, _22205_, _09299_);
  or (_22207_, _22114_, _09297_);
  nand (_22208_, _09297_, _06146_);
  and (_22209_, _22208_, _02954_);
  and (_22210_, _22209_, _22207_);
  or (_22211_, _22210_, _03029_);
  or (_22214_, _22211_, _22206_);
  nor (_22215_, _22112_, _09276_);
  and (_22216_, _09276_, _06147_);
  or (_22217_, _22216_, _09279_);
  or (_22218_, _22217_, _22215_);
  and (_22219_, _22218_, _09250_);
  and (_22220_, _22219_, _22214_);
  or (_22221_, _22220_, _22107_);
  and (_22222_, _22221_, _06246_);
  and (_22223_, _05507_, _02871_);
  or (_22225_, _22223_, _09257_);
  or (_22226_, _22225_, _22222_);
  or (_22227_, _05302_, _02591_);
  and (_22228_, _22227_, _09262_);
  and (_22229_, _22228_, _22226_);
  or (_22230_, _22229_, _22105_);
  and (_22231_, _22230_, _09309_);
  nor (_22232_, _22093_, _09309_);
  or (_22233_, _22232_, _02941_);
  or (_22234_, _22233_, _22231_);
  nand (_22236_, _05269_, _02941_);
  and (_22237_, _22236_, _02589_);
  and (_22238_, _22237_, _22234_);
  and (_22239_, _05302_, _19627_);
  or (_22240_, _22239_, _02940_);
  or (_22241_, _22240_, _22238_);
  nand (_22242_, _05269_, _02940_);
  and (_22243_, _22242_, _09320_);
  and (_22244_, _22243_, _22241_);
  or (_22245_, _22244_, _22104_);
  and (_22247_, _22245_, _09324_);
  nor (_22248_, _09324_, _05269_);
  or (_22249_, _22248_, _07721_);
  or (_22250_, _22249_, _22247_);
  nor (_22251_, _22106_, _02571_);
  nor (_22252_, _22251_, _02866_);
  and (_22253_, _22252_, _22250_);
  or (_22254_, _22253_, _22103_);
  and (_22255_, _22254_, _04134_);
  and (_22256_, _05302_, _02569_);
  or (_22258_, _22256_, _03046_);
  or (_22259_, _22258_, _22255_);
  nand (_22260_, _06146_, _03046_);
  and (_22261_, _22260_, _02860_);
  and (_22262_, _22261_, _22259_);
  nor (_22263_, _05269_, _02860_);
  or (_22264_, _22263_, _02567_);
  or (_22265_, _22264_, _22262_);
  nor (_22266_, _09352_, _06146_);
  or (_22267_, _22266_, _09353_);
  and (_22269_, _22267_, _22265_);
  and (_22270_, _22106_, _09352_);
  or (_22271_, _22270_, _02930_);
  or (_22272_, _22271_, _22269_);
  nand (_22273_, _05269_, _02930_);
  and (_22274_, _22273_, _02517_);
  and (_22275_, _22274_, _22272_);
  and (_22276_, _05302_, _02516_);
  or (_22277_, _22276_, _09362_);
  or (_22278_, _22277_, _22275_);
  nand (_22280_, _22123_, _09362_);
  and (_22281_, _22280_, _05748_);
  and (_22282_, _22281_, _22278_);
  nor (_22283_, _05748_, _05269_);
  or (_22284_, _22283_, _02834_);
  or (_22285_, _22284_, _22282_);
  nand (_22286_, _06146_, _02834_);
  and (_22287_, _22286_, _07831_);
  and (_22288_, _22287_, _22285_);
  and (_22289_, _07830_, _05507_);
  or (_22291_, _22289_, _22288_);
  and (_22292_, _22291_, _19622_);
  or (_22293_, _09382_, _09381_);
  and (_22294_, _22293_, _09401_);
  nor (_22295_, _22293_, _09401_);
  or (_22296_, _22295_, _22294_);
  and (_22297_, _22296_, _09376_);
  or (_22298_, _22297_, _02928_);
  or (_22299_, _22298_, _22292_);
  nand (_22300_, _05269_, _02928_);
  and (_22302_, _22300_, _04131_);
  and (_22303_, _22302_, _22299_);
  and (_22304_, _05302_, _02522_);
  or (_22305_, _22304_, _09419_);
  or (_22306_, _22305_, _22303_);
  nor (_22307_, _22123_, _08166_);
  or (_22308_, _09447_, _05269_);
  nand (_22309_, _22308_, _09419_);
  or (_22310_, _22309_, _22307_);
  and (_22311_, _22310_, _08823_);
  and (_22313_, _22311_, _22306_);
  or (_22314_, _22313_, _22101_);
  and (_22315_, _22314_, _08822_);
  nor (_22316_, _08822_, _05269_);
  or (_22317_, _22316_, _03051_);
  or (_22318_, _22317_, _22315_);
  nand (_22319_, _06146_, _03051_);
  and (_22320_, _22319_, _07150_);
  and (_22321_, _22320_, _22318_);
  and (_22322_, _05507_, _03148_);
  or (_22324_, _22322_, _22321_);
  and (_22325_, _22324_, _19618_);
  and (_22326_, _05302_, _02524_);
  or (_22327_, _22326_, _09441_);
  or (_22328_, _22327_, _22325_);
  nor (_22329_, _22123_, _09447_);
  or (_22330_, _08166_, _05269_);
  nand (_22331_, _22330_, _09441_);
  or (_22332_, _22331_, _22329_);
  and (_22333_, _22332_, _09453_);
  and (_22335_, _22333_, _22328_);
  or (_22336_, _22335_, _22100_);
  and (_22337_, _22336_, _09455_);
  nor (_22338_, _09455_, _05269_);
  or (_22339_, _22338_, _03022_);
  or (_22340_, _22339_, _22337_);
  nand (_22341_, _06146_, _03022_);
  and (_22342_, _22341_, _06213_);
  and (_22343_, _22342_, _22340_);
  and (_22344_, _05507_, _03137_);
  or (_22346_, _22344_, _22343_);
  and (_22347_, _22346_, _19615_);
  and (_22348_, _05302_, _02530_);
  or (_22349_, _22348_, _08818_);
  or (_22350_, _22349_, _22347_);
  nor (_22351_, _22123_, \oc8051_golden_model_1.PSW [7]);
  or (_22352_, _05269_, _07288_);
  nand (_22353_, _22352_, _08818_);
  or (_22354_, _22353_, _22351_);
  and (_22355_, _22354_, _08815_);
  and (_22357_, _22355_, _22350_);
  or (_22358_, _22357_, _22099_);
  and (_22359_, _22358_, _08812_);
  nor (_22360_, _08812_, _05269_);
  or (_22361_, _22360_, _03042_);
  or (_22362_, _22361_, _22359_);
  nand (_22363_, _06146_, _03042_);
  and (_22364_, _22363_, _07161_);
  and (_22365_, _22364_, _22362_);
  and (_22366_, _05507_, _03143_);
  or (_22368_, _22366_, _22365_);
  and (_22369_, _22368_, _02534_);
  and (_22370_, _05302_, _02533_);
  or (_22371_, _22370_, _08808_);
  or (_22372_, _22371_, _22369_);
  or (_22373_, _22123_, _07288_);
  or (_22374_, _05269_, \oc8051_golden_model_1.PSW [7]);
  and (_22375_, _22374_, _08808_);
  and (_22376_, _22375_, _22373_);
  nor (_22377_, _22376_, _09487_);
  and (_22379_, _22377_, _22372_);
  or (_22380_, _22379_, _22098_);
  and (_22381_, _22380_, _07965_);
  nor (_22382_, _07965_, _05269_);
  or (_22383_, _22382_, _07995_);
  or (_22384_, _22383_, _22381_);
  nand (_22385_, _22093_, _07995_);
  and (_22386_, _22385_, _20557_);
  and (_22387_, _22386_, _22384_);
  and (_22388_, _05810_, _03155_);
  or (_22390_, _22388_, _22387_);
  and (_22391_, _22390_, _05790_);
  and (_22392_, _05302_, _02528_);
  or (_22393_, _22392_, _03040_);
  or (_22394_, _22393_, _22391_);
  nor (_22395_, _09692_, _06146_);
  and (_22396_, _22114_, _09692_);
  or (_22397_, _22396_, _03223_);
  or (_22398_, _22397_, _22395_);
  and (_22399_, _22398_, _08803_);
  and (_22401_, _22399_, _22394_);
  or (_22402_, _22401_, _22097_);
  and (_22403_, _22402_, _08789_);
  and (_22404_, _08112_, _05507_);
  or (_22405_, _22404_, _08115_);
  or (_22406_, _22405_, _22403_);
  nand (_22407_, _22093_, _08115_);
  and (_22408_, _22407_, _02891_);
  and (_22409_, _22408_, _22406_);
  and (_22410_, _05810_, _02890_);
  or (_22412_, _22410_, _22409_);
  and (_22413_, _22412_, _08788_);
  and (_22414_, _05302_, _02510_);
  or (_22415_, _22414_, _02889_);
  or (_22416_, _22415_, _22413_);
  and (_22417_, _09692_, _06147_);
  nor (_22418_, _22112_, _09692_);
  nor (_22419_, _22418_, _22417_);
  nand (_22420_, _22419_, _02889_);
  and (_22421_, _22420_, _09724_);
  and (_22423_, _22421_, _22416_);
  nor (_22424_, _22093_, _09724_);
  or (_22425_, _22424_, _03174_);
  or (_22426_, _22425_, _22423_);
  and (_22427_, _22426_, _22096_);
  nor (_22428_, _22427_, _09733_);
  nor (_22429_, _22106_, _09732_);
  nor (_22430_, _22429_, _04150_);
  not (_22431_, _22430_);
  nor (_22432_, _22431_, _22428_);
  and (_22434_, _05302_, _04150_);
  nor (_22435_, _22434_, _02799_);
  not (_22436_, _22435_);
  nor (_22437_, _22436_, _22432_);
  nor (_22438_, _22419_, _09748_);
  nor (_22439_, _22438_, _20609_);
  nor (_22440_, _22439_, _22437_);
  nor (_22441_, _22093_, _09747_);
  nor (_22442_, _22441_, _02887_);
  not (_22443_, _22442_);
  nor (_22445_, _22443_, _22440_);
  and (_22446_, _09755_, _05507_);
  nor (_22447_, _22446_, _20617_);
  nor (_22448_, _22447_, _22445_);
  nor (_22449_, _22093_, _09755_);
  nor (_22450_, _22449_, _22448_);
  nor (_22451_, _22450_, _19863_);
  or (_22452_, _22451_, _08786_);
  nor (_22453_, _22452_, _22095_);
  or (_22454_, _22453_, _22094_);
  or (_22456_, _22454_, _34659_);
  or (_22457_, _34655_, \oc8051_golden_model_1.PC [7]);
  and (_22458_, _22457_, _35796_);
  and (_35842_[7], _22458_, _22456_);
  and (_22459_, _03036_, _02833_);
  and (_22460_, _03034_, _02833_);
  nor (_22461_, _08808_, _02533_);
  and (_22462_, _08921_, _03022_);
  and (_22463_, _08921_, _03051_);
  or (_22464_, _22463_, _03148_);
  nor (_22466_, _09362_, _02516_);
  nor (_22467_, _08792_, \oc8051_golden_model_1.PC [8]);
  nor (_22468_, _22467_, _08793_);
  nor (_22469_, _22468_, _02571_);
  and (_22470_, _22468_, _09249_);
  and (_22471_, _09276_, _08920_);
  nor (_22472_, _08924_, _08918_);
  nor (_22473_, _22472_, _08925_);
  and (_22474_, _22473_, _09277_);
  or (_22475_, _22474_, _22471_);
  and (_22477_, _22475_, _03029_);
  or (_22478_, _22473_, _09297_);
  nand (_22479_, _09297_, _08921_);
  and (_22480_, _22479_, _02954_);
  and (_22481_, _22480_, _22478_);
  or (_22482_, _22481_, _22477_);
  or (_22483_, _22482_, _22470_);
  nor (_22484_, _02876_, _08989_);
  and (_22485_, _09097_, _02877_);
  and (_22486_, _09102_, _09095_);
  nor (_22488_, _22486_, _09103_);
  and (_22489_, _22488_, _19652_);
  and (_22490_, _19659_, _09097_);
  nor (_22491_, _22490_, _22489_);
  nand (_22492_, _22491_, _09132_);
  not (_22493_, _22468_);
  and (_22494_, _22493_, _03840_);
  nor (_22495_, _22494_, _02948_);
  and (_22496_, _22468_, _07436_);
  and (_22497_, _09153_, _09145_);
  or (_22499_, _22497_, _22468_);
  and (_22500_, _09153_, _02603_);
  nand (_22501_, _09098_, _03845_);
  or (_22502_, _03845_, \oc8051_golden_model_1.PC [8]);
  or (_22503_, _22502_, _09138_);
  and (_22504_, _22503_, _22501_);
  nor (_22505_, _22504_, _21404_);
  nand (_22506_, _22505_, _22500_);
  and (_22507_, _22506_, _22499_);
  or (_22508_, _22507_, _02951_);
  and (_22510_, _09098_, _02951_);
  nor (_22511_, _22510_, _07436_);
  and (_22512_, _22511_, _22508_);
  or (_22513_, _22512_, _09169_);
  nor (_22514_, _22513_, _22496_);
  nor (_22515_, _22514_, _07433_);
  and (_22516_, _22468_, _07433_);
  nor (_22517_, _22516_, _03840_);
  nand (_22518_, _22517_, _05361_);
  or (_22519_, _22518_, _22515_);
  and (_22521_, _22519_, _22495_);
  nand (_22522_, _22521_, _22492_);
  not (_22523_, _22473_);
  or (_22524_, _22523_, _09003_);
  nand (_22525_, _09003_, _08920_);
  and (_22526_, _22525_, _22524_);
  or (_22527_, _22526_, _03006_);
  and (_22528_, _22527_, _22522_);
  or (_22529_, _22528_, _08998_);
  or (_22530_, _22493_, _08997_);
  and (_22532_, _22530_, _02934_);
  and (_22533_, _22532_, _22529_);
  nor (_22534_, _02946_, _04225_);
  nand (_22535_, _09098_, _02884_);
  nand (_22536_, _22535_, _22534_);
  or (_22537_, _22536_, _22533_);
  and (_22538_, _09097_, _02946_);
  nor (_22539_, _22538_, _09187_);
  nand (_22540_, _22539_, _22537_);
  nor (_22541_, _22468_, _09186_);
  nor (_22543_, _22541_, _02880_);
  nand (_22544_, _22543_, _22540_);
  and (_22545_, _09097_, _02880_);
  nor (_22546_, _22545_, _09193_);
  nand (_22547_, _22546_, _22544_);
  and (_22548_, _22493_, _09193_);
  nor (_22549_, _22548_, _02877_);
  and (_22550_, _22549_, _22547_);
  or (_22551_, _22550_, _22485_);
  nand (_22552_, _22551_, _22484_);
  and (_22554_, _09097_, _02876_);
  nor (_22555_, _22554_, _09210_);
  and (_22556_, _22555_, _22552_);
  and (_22557_, _09242_, _08920_);
  nor (_22558_, _22523_, _09242_);
  or (_22559_, _22558_, _22557_);
  nor (_22560_, _22559_, _09209_);
  or (_22561_, _22560_, _22556_);
  nand (_22562_, _22561_, _08986_);
  and (_22563_, _09918_, _08920_);
  and (_22565_, _22473_, _08981_);
  nor (_22566_, _22565_, _22563_);
  nand (_22567_, _22566_, _08985_);
  and (_22568_, _22567_, _22562_);
  and (_22569_, _22568_, _09251_);
  or (_22570_, _22569_, _22483_);
  and (_22571_, _09262_, _06246_);
  and (_22572_, _22571_, _22570_);
  nor (_22573_, _22571_, _09098_);
  nand (_22574_, _09309_, _02591_);
  or (_22576_, _22574_, _22573_);
  or (_22577_, _22576_, _22572_);
  nor (_22578_, _22468_, _09309_);
  nor (_22579_, _22578_, _02941_);
  nand (_22580_, _22579_, _22577_);
  and (_22581_, _09097_, _02941_);
  nor (_22582_, _22581_, _19627_);
  nand (_22583_, _22582_, _22580_);
  nand (_22584_, _22583_, _10030_);
  and (_22585_, _09097_, _02940_);
  nor (_22587_, _22585_, _09326_);
  nand (_22588_, _22587_, _22584_);
  nor (_22589_, _22468_, _09320_);
  nor (_22590_, _22589_, _09325_);
  nand (_22591_, _22590_, _22588_);
  nor (_22592_, _09324_, _09098_);
  nor (_22593_, _22592_, _07721_);
  and (_22594_, _22593_, _22591_);
  or (_22595_, _22594_, _22469_);
  nand (_22596_, _22595_, _02986_);
  and (_22598_, _09098_, _02866_);
  nor (_22599_, _03046_, _02569_);
  not (_22600_, _22599_);
  nor (_22601_, _22600_, _22598_);
  nand (_22602_, _22601_, _22596_);
  and (_22603_, _08920_, _03046_);
  not (_22604_, _22603_);
  and (_22605_, _22604_, _02860_);
  nand (_22606_, _22605_, _22602_);
  nor (_22607_, _09097_, _02860_);
  nor (_22609_, _22607_, _02567_);
  and (_22610_, _22609_, _22606_);
  and (_22611_, _08920_, _02567_);
  or (_22612_, _22611_, _09352_);
  or (_22613_, _22612_, _22610_);
  and (_22614_, _22493_, _09352_);
  nor (_22615_, _22614_, _02930_);
  and (_22616_, _22615_, _22613_);
  and (_22617_, _09097_, _02930_);
  or (_22618_, _22617_, _22616_);
  nand (_22620_, _22618_, _22466_);
  and (_22621_, _22488_, _09362_);
  nor (_22622_, _22621_, _05749_);
  and (_22623_, _22622_, _22620_);
  nor (_22624_, _09097_, _05748_);
  or (_22625_, _22624_, _22623_);
  nand (_22626_, _22625_, _07140_);
  and (_22627_, _08921_, _02834_);
  nor (_22628_, _22627_, _07830_);
  nand (_22629_, _22628_, _22626_);
  and (_22631_, _09097_, _07830_);
  nor (_22632_, _22631_, _09376_);
  nand (_22633_, _22632_, _22629_);
  and (_22634_, _09403_, _09380_);
  nor (_22635_, _22634_, _09404_);
  nor (_22636_, _22635_, _19622_);
  nor (_22637_, _22636_, _02928_);
  nand (_22638_, _22637_, _22633_);
  and (_22639_, _09097_, _02928_);
  nor (_22640_, _22639_, _02522_);
  nand (_22642_, _22640_, _22638_);
  nand (_22643_, _22642_, _19621_);
  and (_22644_, _09097_, _08166_);
  and (_22645_, _22488_, _09447_);
  or (_22646_, _22645_, _22644_);
  and (_22647_, _22646_, _09419_);
  nor (_22648_, _22647_, _09428_);
  nand (_22649_, _22648_, _22643_);
  nor (_22650_, _22468_, _08823_);
  nor (_22651_, _22650_, _21199_);
  nand (_22653_, _22651_, _22649_);
  nor (_22654_, _09098_, _08822_);
  nor (_22655_, _22654_, _03051_);
  and (_22656_, _22655_, _22653_);
  or (_22657_, _22656_, _22464_);
  and (_22658_, _09097_, _03148_);
  nor (_22659_, _22658_, _02524_);
  nand (_22660_, _22659_, _22657_);
  nand (_22661_, _22660_, _09446_);
  nor (_22662_, _22488_, _09447_);
  nor (_22664_, _09097_, _08166_);
  nor (_22665_, _22664_, _09446_);
  not (_22666_, _22665_);
  nor (_22667_, _22666_, _22662_);
  nor (_22668_, _22667_, _20129_);
  nand (_22669_, _22668_, _22661_);
  nor (_22670_, _22468_, _09453_);
  nor (_22671_, _22670_, _09456_);
  nand (_22672_, _22671_, _22669_);
  nor (_22673_, _09098_, _09455_);
  nor (_22675_, _22673_, _03022_);
  and (_22676_, _22675_, _22672_);
  or (_22677_, _22676_, _22462_);
  nand (_22678_, _22677_, _06213_);
  nor (_22679_, _08818_, _02530_);
  and (_22680_, _09098_, _03137_);
  not (_22681_, _22680_);
  and (_22682_, _22681_, _22679_);
  nand (_22683_, _22682_, _22678_);
  or (_22684_, _22488_, \oc8051_golden_model_1.PSW [7]);
  or (_22686_, _09097_, _07288_);
  and (_22687_, _22686_, _08818_);
  and (_22688_, _22687_, _22684_);
  nor (_22689_, _22688_, _09468_);
  nand (_22690_, _22689_, _22683_);
  nor (_22691_, _22468_, _08815_);
  nor (_22692_, _22691_, _13433_);
  and (_22693_, _22692_, _22690_);
  nor (_22694_, _09098_, _08812_);
  or (_22695_, _22694_, _03042_);
  or (_22697_, _22695_, _22693_);
  and (_22698_, _08921_, _03042_);
  nor (_22699_, _22698_, _03143_);
  and (_22700_, _22699_, _22697_);
  and (_22701_, _09097_, _03143_);
  or (_22702_, _22701_, _22700_);
  nand (_22703_, _22702_, _22461_);
  or (_22704_, _22488_, _07288_);
  or (_22705_, _09097_, \oc8051_golden_model_1.PSW [7]);
  and (_22706_, _22705_, _08808_);
  and (_22708_, _22706_, _22704_);
  nor (_22709_, _22708_, _09487_);
  nand (_22710_, _22709_, _22703_);
  nor (_22711_, _22468_, _08806_);
  nor (_22712_, _22711_, _07966_);
  and (_22713_, _22712_, _22710_);
  nor (_22714_, _09098_, _07965_);
  or (_22715_, _22714_, _07995_);
  or (_22716_, _22715_, _22713_);
  and (_22717_, _22493_, _07995_);
  nor (_22719_, _22717_, _03155_);
  nand (_22720_, _22719_, _22716_);
  and (_22721_, _03838_, _03155_);
  nor (_22722_, _22721_, _02528_);
  nand (_22723_, _22722_, _22720_);
  nand (_22724_, _22723_, _03223_);
  and (_22725_, _22523_, _09692_);
  nor (_22726_, _09692_, _08920_);
  or (_22727_, _22726_, _03223_);
  or (_22728_, _22727_, _22725_);
  and (_22730_, _22728_, _08803_);
  nand (_22731_, _22730_, _22724_);
  nor (_22732_, _22468_, _08803_);
  nor (_22733_, _22732_, _08112_);
  and (_22734_, _22733_, _22731_);
  and (_22735_, _09097_, _08112_);
  or (_22736_, _22735_, _08115_);
  or (_22737_, _22736_, _22734_);
  and (_22738_, _22493_, _08115_);
  nor (_22739_, _22738_, _02890_);
  nand (_22741_, _22739_, _22737_);
  and (_22742_, _03838_, _02890_);
  nor (_22743_, _22742_, _02510_);
  nand (_22744_, _22743_, _22741_);
  nand (_22745_, _22744_, _03175_);
  and (_22746_, _09692_, _08921_);
  nor (_22747_, _22473_, _09692_);
  nor (_22748_, _22747_, _22746_);
  and (_22749_, _22748_, _02889_);
  nor (_22750_, _22749_, _09725_);
  nand (_22752_, _22750_, _22745_);
  nor (_22753_, _22468_, _09724_);
  nor (_22754_, _22753_, _03174_);
  nand (_22755_, _22754_, _22752_);
  and (_22756_, _09097_, _03174_);
  nor (_22757_, _22756_, _09733_);
  nand (_22758_, _22757_, _22755_);
  nor (_22759_, _22468_, _09732_);
  nor (_22760_, _22759_, _03034_);
  and (_22761_, _22760_, _22758_);
  or (_22763_, _22761_, _22460_);
  nor (_22764_, _02799_, _02505_);
  nand (_22765_, _22764_, _22763_);
  and (_22766_, _22748_, _02799_);
  nor (_22767_, _22766_, _09748_);
  nand (_22768_, _22767_, _22765_);
  nor (_22769_, _22468_, _09747_);
  nor (_22770_, _22769_, _02887_);
  nand (_22771_, _22770_, _22768_);
  and (_22772_, _09097_, _02887_);
  nor (_22774_, _22772_, _09756_);
  nand (_22775_, _22774_, _22771_);
  nor (_22776_, _22468_, _09755_);
  nor (_22777_, _22776_, _03036_);
  and (_22778_, _22777_, _22775_);
  or (_22779_, _22778_, _22459_);
  nor (_22780_, _08786_, _02499_);
  and (_22781_, _22780_, _22779_);
  and (_22782_, _22468_, _08786_);
  or (_22783_, _22782_, _22781_);
  or (_22785_, _22783_, _34659_);
  or (_22786_, _34655_, \oc8051_golden_model_1.PC [8]);
  and (_22787_, _22786_, _35796_);
  and (_35842_[8], _22787_, _22785_);
  nor (_22788_, _03687_, _03038_);
  nor (_22789_, _03687_, _06185_);
  nor (_22790_, _08793_, \oc8051_golden_model_1.PC [9]);
  nor (_22791_, _22790_, _08794_);
  nor (_22792_, _22791_, _08803_);
  nor (_22793_, _22791_, _08806_);
  and (_22795_, _08858_, _03042_);
  nor (_22796_, _22791_, _08815_);
  and (_22797_, _08858_, _03022_);
  nor (_22798_, _22791_, _09453_);
  and (_22799_, _08858_, _03051_);
  nor (_22800_, _22791_, _08823_);
  and (_22801_, _09043_, _02940_);
  nor (_22802_, _02940_, _19627_);
  and (_22803_, _09043_, _02941_);
  nor (_22804_, _08925_, _08922_);
  and (_22806_, _22804_, _08863_);
  nor (_22807_, _22804_, _08863_);
  nor (_22808_, _22807_, _22806_);
  not (_22809_, _22808_);
  or (_22810_, _22809_, _09918_);
  or (_22811_, _08981_, _08858_);
  and (_22812_, _22811_, _08985_);
  and (_22813_, _22812_, _22810_);
  nor (_22814_, _09103_, _09099_);
  and (_22815_, _22814_, _09047_);
  nor (_22817_, _22814_, _09047_);
  nor (_22818_, _22817_, _22815_);
  nor (_22819_, _22818_, _09012_);
  and (_22820_, _19659_, _09043_);
  or (_22821_, _22820_, _22819_);
  nor (_22822_, _22821_, _05361_);
  not (_22823_, _22791_);
  and (_22824_, _22823_, _03840_);
  nor (_22825_, _22824_, _02948_);
  and (_22826_, _22823_, _07436_);
  and (_22828_, _09043_, _02951_);
  nor (_22829_, _22791_, _22497_);
  and (_22830_, _09044_, _03845_);
  nor (_22831_, _03845_, \oc8051_golden_model_1.PC [9]);
  and (_22832_, _22831_, _09144_);
  nor (_22833_, _22832_, _22830_);
  nor (_22834_, _22833_, _21404_);
  and (_22835_, _22834_, _22500_);
  nor (_22836_, _22835_, _02951_);
  nor (_22837_, _22836_, _07436_);
  nor (_22839_, _22837_, _22829_);
  nor (_22840_, _22839_, _22828_);
  nor (_22841_, _22840_, _22826_);
  nor (_22842_, _22841_, _09169_);
  nor (_22843_, _22842_, _07433_);
  and (_22844_, _22791_, _07433_);
  nor (_22845_, _22844_, _03840_);
  nand (_22846_, _22845_, _05361_);
  or (_22847_, _22846_, _22843_);
  nand (_22848_, _22847_, _22825_);
  nor (_22850_, _22848_, _22822_);
  or (_22851_, _22809_, _19674_);
  nand (_22852_, _19673_, _10785_);
  or (_22853_, _22852_, _08858_);
  and (_22854_, _22853_, _02948_);
  and (_22855_, _22854_, _22851_);
  or (_22856_, _22855_, _08998_);
  nor (_22857_, _22856_, _22850_);
  nor (_22858_, _22791_, _08997_);
  nor (_22859_, _22858_, _02884_);
  not (_22861_, _22859_);
  nor (_22862_, _22861_, _22857_);
  and (_22863_, _09044_, _02597_);
  nor (_22864_, _22863_, _08993_);
  nor (_22865_, _22864_, _22862_);
  nor (_22866_, _22865_, _02946_);
  and (_22867_, _09043_, _02946_);
  nor (_22868_, _22867_, _09187_);
  not (_22869_, _22868_);
  nor (_22870_, _22869_, _22866_);
  nor (_22872_, _22791_, _09186_);
  nor (_22873_, _22872_, _02880_);
  not (_22874_, _22873_);
  nor (_22875_, _22874_, _22870_);
  and (_22876_, _09043_, _02880_);
  nor (_22877_, _22876_, _09193_);
  not (_22878_, _22877_);
  nor (_22879_, _22878_, _22875_);
  and (_22880_, _22823_, _09193_);
  nor (_22881_, _22880_, _02877_);
  not (_22882_, _22881_);
  nor (_22883_, _22882_, _22879_);
  and (_22884_, _09043_, _02877_);
  or (_22885_, _22884_, _22883_);
  or (_22886_, _22885_, _08989_);
  nand (_22887_, _22886_, _03962_);
  and (_22888_, _09043_, _02876_);
  nor (_22889_, _22888_, _09210_);
  nand (_22890_, _22889_, _22887_);
  and (_22891_, _09242_, _08858_);
  nor (_22894_, _22808_, _09242_);
  or (_22895_, _22894_, _22891_);
  nor (_22896_, _22895_, _09209_);
  nor (_22897_, _22896_, _08985_);
  and (_22898_, _22897_, _22890_);
  or (_22899_, _22898_, _22813_);
  nand (_22900_, _22899_, _09251_);
  nor (_22901_, _22808_, _09297_);
  and (_22902_, _09297_, _08858_);
  nor (_22903_, _22902_, _22901_);
  nor (_22905_, _22903_, _09299_);
  and (_22906_, _22808_, _09277_);
  and (_22907_, _09276_, _08859_);
  nor (_22908_, _22907_, _09279_);
  not (_22909_, _22908_);
  nor (_22910_, _22909_, _22906_);
  nor (_22911_, _22910_, _22905_);
  and (_22912_, _22791_, _09249_);
  nor (_22913_, _22912_, _02871_);
  and (_22914_, _22913_, _22911_);
  and (_22915_, _22914_, _22900_);
  and (_22916_, _09044_, _02871_);
  nor (_22917_, _22916_, _22915_);
  and (_22918_, _09262_, _02591_);
  nand (_22919_, _22918_, _22917_);
  nor (_22920_, _09262_, _09044_);
  nor (_22921_, _22920_, _09310_);
  nand (_22922_, _22921_, _22919_);
  nor (_22923_, _22791_, _09309_);
  nor (_22924_, _22923_, _02941_);
  and (_22926_, _22924_, _22922_);
  or (_22927_, _22926_, _22803_);
  and (_22928_, _22927_, _22802_);
  or (_22929_, _22928_, _22801_);
  nand (_22930_, _22929_, _09320_);
  nor (_22931_, _22823_, _09320_);
  nor (_22932_, _22931_, _09325_);
  nand (_22933_, _22932_, _22930_);
  nor (_22934_, _09324_, _09043_);
  nor (_22935_, _22934_, _07721_);
  nand (_22937_, _22935_, _22933_);
  nor (_22938_, _22823_, _02571_);
  nor (_22939_, _22938_, _02866_);
  nand (_22940_, _22939_, _22937_);
  and (_22941_, _09044_, _02866_);
  nor (_22942_, _22941_, _22600_);
  nand (_22943_, _22942_, _22940_);
  and (_22944_, _08858_, _03046_);
  not (_22945_, _22944_);
  and (_22946_, _22945_, _02860_);
  nand (_22947_, _22946_, _22943_);
  nor (_22948_, _09043_, _02860_);
  nor (_22949_, _22948_, _02567_);
  and (_22950_, _22949_, _22947_);
  nor (_22951_, _09352_, _08858_);
  nor (_22952_, _22951_, _09353_);
  or (_22953_, _22952_, _22950_);
  and (_22954_, _22823_, _09352_);
  nor (_22955_, _22954_, _02930_);
  and (_22956_, _22955_, _22953_);
  and (_22958_, _09043_, _02930_);
  or (_22959_, _22958_, _22956_);
  nand (_22960_, _22959_, _22466_);
  nor (_22961_, _22818_, _09366_);
  nor (_22962_, _22961_, _05749_);
  nand (_22963_, _22962_, _22960_);
  nor (_22964_, _09043_, _05748_);
  nor (_22965_, _22964_, _02834_);
  and (_22966_, _22965_, _22963_);
  and (_22967_, _08858_, _02834_);
  or (_22968_, _22967_, _07830_);
  nor (_22969_, _22968_, _22966_);
  and (_22970_, _09044_, _07830_);
  or (_22971_, _22970_, _22969_);
  nand (_22972_, _22971_, _19622_);
  nor (_22973_, _09404_, \oc8051_golden_model_1.DPH [1]);
  nor (_22974_, _22973_, _09405_);
  nor (_22975_, _22974_, _19622_);
  nor (_22976_, _22975_, _02928_);
  nand (_22977_, _22976_, _22972_);
  and (_22978_, _09043_, _02928_);
  nor (_22979_, _22978_, _02522_);
  nand (_22980_, _22979_, _22977_);
  nand (_22981_, _22980_, _19621_);
  and (_22982_, _09043_, _08166_);
  nor (_22983_, _22818_, _08166_);
  or (_22984_, _22983_, _22982_);
  and (_22985_, _22984_, _09419_);
  nor (_22986_, _22985_, _09428_);
  and (_22987_, _22986_, _22981_);
  or (_22988_, _22987_, _22800_);
  nand (_22989_, _22988_, _08822_);
  nor (_22990_, _09043_, _08822_);
  nor (_22991_, _22990_, _03051_);
  and (_22992_, _22991_, _22989_);
  or (_22993_, _22992_, _22799_);
  nand (_22994_, _22993_, _07150_);
  and (_22995_, _09043_, _03148_);
  nor (_22996_, _22995_, _02524_);
  nand (_22997_, _22996_, _22994_);
  nand (_22998_, _22997_, _09446_);
  and (_22999_, _22818_, _08166_);
  nor (_23000_, _09043_, _08166_);
  nor (_23001_, _23000_, _09446_);
  not (_23002_, _23001_);
  nor (_23003_, _23002_, _22999_);
  nor (_23004_, _23003_, _20129_);
  and (_23005_, _23004_, _22998_);
  or (_23006_, _23005_, _22798_);
  nand (_23007_, _23006_, _09455_);
  nor (_23008_, _09043_, _09455_);
  nor (_23009_, _23008_, _03022_);
  and (_23010_, _23009_, _23007_);
  or (_23011_, _23010_, _22797_);
  nand (_23012_, _23011_, _06213_);
  and (_23013_, _09043_, _03137_);
  nor (_23014_, _23013_, _02530_);
  nand (_23015_, _23014_, _23012_);
  nand (_23016_, _23015_, _09470_);
  and (_23017_, _22818_, _07288_);
  nor (_23020_, _09043_, _07288_);
  nor (_23021_, _23020_, _09470_);
  not (_23022_, _23021_);
  nor (_23023_, _23022_, _23017_);
  nor (_23024_, _23023_, _09468_);
  and (_23025_, _23024_, _23016_);
  or (_23026_, _23025_, _22796_);
  nand (_23027_, _23026_, _08812_);
  nor (_23028_, _09043_, _08812_);
  nor (_23029_, _23028_, _03042_);
  and (_23030_, _23029_, _23027_);
  or (_23031_, _23030_, _22795_);
  nand (_23032_, _23031_, _07161_);
  and (_23033_, _09043_, _03143_);
  nor (_23034_, _23033_, _02533_);
  nand (_23035_, _23034_, _23032_);
  nand (_23036_, _23035_, _19607_);
  nand (_23037_, _22818_, \oc8051_golden_model_1.PSW [7]);
  or (_23038_, _09043_, \oc8051_golden_model_1.PSW [7]);
  and (_23039_, _23038_, _08808_);
  and (_23040_, _23039_, _23037_);
  nor (_23041_, _23040_, _09487_);
  and (_23042_, _23041_, _23036_);
  or (_23043_, _23042_, _22793_);
  nand (_23044_, _23043_, _07965_);
  nor (_23045_, _09043_, _07965_);
  nor (_23046_, _23045_, _07995_);
  nand (_23047_, _23046_, _23044_);
  and (_23048_, _22791_, _07995_);
  nor (_23049_, _23048_, _03155_);
  nand (_23052_, _23049_, _23047_);
  nor (_23053_, _03040_, _02528_);
  not (_23054_, _23053_);
  and (_23055_, _04020_, _03155_);
  nor (_23056_, _23055_, _23054_);
  nand (_23057_, _23056_, _23052_);
  nor (_23058_, _09692_, _08858_);
  and (_23059_, _22808_, _09692_);
  or (_23060_, _23059_, _03223_);
  or (_23061_, _23060_, _23058_);
  and (_23063_, _23061_, _08803_);
  and (_23064_, _23063_, _23057_);
  or (_23065_, _23064_, _22792_);
  nand (_23066_, _23065_, _08789_);
  and (_23067_, _09044_, _08112_);
  nor (_23068_, _23067_, _08115_);
  nand (_23069_, _23068_, _23066_);
  and (_23070_, _22791_, _08115_);
  nor (_23071_, _23070_, _02890_);
  nand (_23072_, _23071_, _23069_);
  and (_23073_, _04020_, _02890_);
  nor (_23074_, _02889_, _02510_);
  not (_23075_, _23074_);
  nor (_23076_, _23075_, _23073_);
  nand (_23077_, _23076_, _23072_);
  nor (_23078_, _22809_, _09692_);
  and (_23079_, _09692_, _08859_);
  nor (_23080_, _23079_, _23078_);
  and (_23081_, _23080_, _02889_);
  nor (_23082_, _23081_, _09725_);
  nand (_23084_, _23082_, _23077_);
  nor (_23085_, _22791_, _09724_);
  nor (_23086_, _23085_, _03174_);
  nand (_23087_, _23086_, _23084_);
  and (_23088_, _09043_, _03174_);
  nor (_23089_, _23088_, _09733_);
  nand (_23090_, _23089_, _23087_);
  nor (_23091_, _22791_, _09732_);
  nor (_23092_, _23091_, _03034_);
  and (_23093_, _23092_, _23090_);
  or (_23095_, _23093_, _22789_);
  nand (_23096_, _23095_, _22764_);
  and (_23097_, _23080_, _02799_);
  nor (_23098_, _23097_, _09748_);
  nand (_23099_, _23098_, _23096_);
  nor (_23100_, _22791_, _09747_);
  nor (_23101_, _23100_, _02887_);
  nand (_23102_, _23101_, _23099_);
  and (_23103_, _09043_, _02887_);
  nor (_23104_, _23103_, _09756_);
  nand (_23106_, _23104_, _23102_);
  nor (_23107_, _22791_, _09755_);
  nor (_23108_, _23107_, _03036_);
  and (_23109_, _23108_, _23106_);
  or (_23110_, _23109_, _22788_);
  and (_23111_, _23110_, _22780_);
  and (_23112_, _22791_, _08786_);
  or (_23113_, _23112_, _23111_);
  or (_23114_, _23113_, _34659_);
  or (_23115_, _34655_, \oc8051_golden_model_1.PC [9]);
  and (_23117_, _23115_, _35796_);
  and (_35842_[9], _23117_, _23114_);
  nor (_23118_, _08794_, \oc8051_golden_model_1.PC [10]);
  nor (_23119_, _23118_, _08795_);
  and (_23120_, _23119_, _08786_);
  nor (_23121_, _23119_, _09724_);
  not (_23122_, _23119_);
  and (_23123_, _23122_, _07995_);
  nor (_23124_, _23119_, _08806_);
  nand (_23125_, _08852_, _03042_);
  nand (_23127_, _08852_, _03022_);
  nand (_23128_, _08852_, _03051_);
  and (_23129_, _08852_, _02567_);
  nor (_23130_, _23129_, _09352_);
  nand (_23131_, _09037_, _02940_);
  and (_23132_, _23119_, _09193_);
  nand (_23133_, _09037_, _02946_);
  and (_23134_, _09036_, _02884_);
  and (_23135_, _09003_, _08851_);
  not (_23136_, _08855_);
  nor (_23138_, _08929_, _08926_);
  nor (_23139_, _23138_, _23136_);
  and (_23140_, _23138_, _23136_);
  nor (_23141_, _23140_, _23139_);
  not (_23142_, _23141_);
  nor (_23143_, _23142_, _09003_);
  or (_23144_, _23143_, _23135_);
  and (_23145_, _23144_, _02948_);
  nor (_23146_, _09107_, _09104_);
  not (_23147_, _23146_);
  and (_23148_, _23147_, _09040_);
  nor (_23149_, _23147_, _09040_);
  nor (_23150_, _23149_, _23148_);
  and (_23151_, _23150_, _19652_);
  and (_23152_, _09012_, _09036_);
  or (_23153_, _23152_, _23151_);
  or (_23154_, _23153_, _05361_);
  nand (_23155_, _23122_, _03840_);
  and (_23156_, _23155_, _03006_);
  or (_23157_, _23119_, _22497_);
  nand (_23159_, _09037_, _03845_);
  or (_23160_, _03845_, \oc8051_golden_model_1.PC [10]);
  or (_23161_, _23160_, _09138_);
  and (_23162_, _23161_, _23159_);
  nor (_23163_, _23162_, _21404_);
  nand (_23164_, _23163_, _22500_);
  and (_23165_, _23164_, _23157_);
  or (_23166_, _23165_, _02951_);
  and (_23167_, _09037_, _02951_);
  nor (_23168_, _23167_, _07436_);
  and (_23170_, _23168_, _23166_);
  and (_23171_, _23119_, _07436_);
  or (_23172_, _23171_, _09169_);
  or (_23173_, _23172_, _23170_);
  and (_23174_, _23173_, _09133_);
  and (_23175_, _23119_, _07433_);
  nor (_23176_, _23175_, _03840_);
  nand (_23177_, _23176_, _05361_);
  or (_23178_, _23177_, _23174_);
  and (_23179_, _23178_, _23156_);
  and (_23181_, _23179_, _23154_);
  or (_23182_, _23181_, _08998_);
  or (_23183_, _23182_, _23145_);
  or (_23184_, _23119_, _08997_);
  and (_23185_, _23184_, _02934_);
  and (_23186_, _23185_, _23183_);
  nor (_23187_, _23186_, _23134_);
  nand (_23188_, _23187_, _22534_);
  and (_23189_, _23188_, _23133_);
  and (_23190_, _23189_, _09186_);
  nor (_23192_, _23122_, _09186_);
  or (_23193_, _23192_, _02880_);
  or (_23194_, _23193_, _23190_);
  and (_23195_, _09037_, _02880_);
  nor (_23196_, _23195_, _09193_);
  and (_23197_, _23196_, _23194_);
  or (_23198_, _23197_, _23132_);
  and (_23199_, _23198_, _02987_);
  and (_23200_, _09036_, _02877_);
  or (_23201_, _23200_, _08989_);
  or (_23203_, _23201_, _23199_);
  and (_23204_, _23203_, _03962_);
  nand (_23205_, _09036_, _02876_);
  nand (_23206_, _23205_, _09209_);
  or (_23207_, _23206_, _23204_);
  and (_23208_, _09242_, _08851_);
  nor (_23209_, _23142_, _09242_);
  or (_23210_, _23209_, _23208_);
  or (_23211_, _23210_, _09209_);
  and (_23212_, _23211_, _23207_);
  or (_23213_, _23212_, _08985_);
  and (_23214_, _23141_, _08981_);
  and (_23215_, _09918_, _08851_);
  or (_23216_, _23215_, _08986_);
  or (_23217_, _23216_, _23214_);
  and (_23218_, _23217_, _09299_);
  and (_23219_, _23218_, _23213_);
  and (_23220_, _09297_, _08851_);
  nor (_23221_, _23142_, _09297_);
  or (_23222_, _23221_, _23220_);
  and (_23224_, _23222_, _02954_);
  or (_23225_, _23224_, _23219_);
  and (_23226_, _23225_, _09279_);
  or (_23227_, _23141_, _09276_);
  nand (_23228_, _09276_, _08852_);
  and (_23229_, _23228_, _03029_);
  and (_23230_, _23229_, _23227_);
  or (_23231_, _23230_, _09249_);
  or (_23232_, _23231_, _23226_);
  nand (_23233_, _23122_, _09249_);
  and (_23235_, _23233_, _22571_);
  and (_23236_, _23235_, _23232_);
  nor (_23237_, _22571_, _09037_);
  or (_23238_, _23237_, _22574_);
  or (_23239_, _23238_, _23236_);
  or (_23240_, _23119_, _09309_);
  and (_23241_, _23240_, _09799_);
  and (_23242_, _23241_, _23239_);
  nand (_23243_, _09036_, _02941_);
  nand (_23244_, _23243_, _22802_);
  or (_23246_, _23244_, _23242_);
  and (_23247_, _23246_, _23131_);
  or (_23248_, _23247_, _09326_);
  or (_23249_, _23119_, _09320_);
  and (_23250_, _23249_, _09324_);
  and (_23251_, _23250_, _23248_);
  nor (_23252_, _09324_, _09037_);
  or (_23253_, _23252_, _07721_);
  or (_23254_, _23253_, _23251_);
  nor (_23255_, _23119_, _02571_);
  nor (_23257_, _23255_, _02866_);
  and (_23258_, _23257_, _23254_);
  nand (_23259_, _09036_, _02866_);
  nand (_23260_, _23259_, _22599_);
  or (_23261_, _23260_, _23258_);
  nand (_23262_, _08852_, _03046_);
  and (_23263_, _23262_, _02860_);
  and (_23264_, _23263_, _23261_);
  nor (_23265_, _09037_, _02860_);
  or (_23266_, _23265_, _02567_);
  or (_23268_, _23266_, _23264_);
  and (_23269_, _23268_, _23130_);
  and (_23270_, _23119_, _09352_);
  or (_23271_, _23270_, _23269_);
  and (_23272_, _23271_, _03508_);
  nand (_23273_, _09036_, _02930_);
  nand (_23274_, _23273_, _22466_);
  or (_23275_, _23274_, _23272_);
  or (_23276_, _23150_, _09366_);
  and (_23277_, _23276_, _05748_);
  and (_23278_, _23277_, _23275_);
  nor (_23279_, _09037_, _05748_);
  or (_23280_, _23279_, _02834_);
  or (_23281_, _23280_, _23278_);
  nand (_23282_, _08852_, _02834_);
  and (_23283_, _23282_, _07831_);
  and (_23284_, _23283_, _23281_);
  and (_23285_, _09036_, _07830_);
  or (_23286_, _23285_, _09376_);
  or (_23287_, _23286_, _23284_);
  nor (_23289_, _09405_, \oc8051_golden_model_1.DPH [2]);
  nor (_23290_, _23289_, _09406_);
  or (_23291_, _23290_, _19622_);
  and (_23292_, _23291_, _23287_);
  or (_23293_, _23292_, _02928_);
  nand (_23294_, _09037_, _02928_);
  nor (_23295_, _09419_, _02522_);
  and (_23296_, _23295_, _23294_);
  and (_23297_, _23296_, _23293_);
  or (_23298_, _23150_, _08166_);
  or (_23300_, _09036_, _09447_);
  and (_23301_, _23300_, _09419_);
  and (_23302_, _23301_, _23298_);
  or (_23303_, _23302_, _09428_);
  or (_23304_, _23303_, _23297_);
  or (_23305_, _23119_, _08823_);
  and (_23306_, _23305_, _08822_);
  and (_23307_, _23306_, _23304_);
  nor (_23308_, _09037_, _08822_);
  or (_23309_, _23308_, _03051_);
  or (_23311_, _23309_, _23307_);
  and (_23312_, _23311_, _23128_);
  or (_23313_, _23312_, _03148_);
  nand (_23314_, _09037_, _03148_);
  nor (_23315_, _09441_, _02524_);
  and (_23316_, _23315_, _23314_);
  and (_23317_, _23316_, _23313_);
  or (_23318_, _23150_, _09447_);
  or (_23319_, _09036_, _08166_);
  and (_23320_, _23319_, _09441_);
  and (_23322_, _23320_, _23318_);
  or (_23323_, _23322_, _20129_);
  or (_23324_, _23323_, _23317_);
  or (_23325_, _23119_, _09453_);
  and (_23326_, _23325_, _09455_);
  and (_23327_, _23326_, _23324_);
  nor (_23328_, _09037_, _09455_);
  or (_23329_, _23328_, _03022_);
  or (_23330_, _23329_, _23327_);
  and (_23331_, _23330_, _23127_);
  or (_23333_, _23331_, _03137_);
  nand (_23334_, _09037_, _03137_);
  and (_23335_, _23334_, _22679_);
  and (_23336_, _23335_, _23333_);
  or (_23337_, _23150_, \oc8051_golden_model_1.PSW [7]);
  or (_23338_, _09036_, _07288_);
  and (_23339_, _23338_, _08818_);
  and (_23340_, _23339_, _23337_);
  or (_23341_, _23340_, _09468_);
  or (_23342_, _23341_, _23336_);
  or (_23343_, _23119_, _08815_);
  and (_23344_, _23343_, _08812_);
  and (_23345_, _23344_, _23342_);
  nor (_23346_, _09037_, _08812_);
  or (_23347_, _23346_, _03042_);
  or (_23348_, _23347_, _23345_);
  and (_23349_, _23348_, _23125_);
  or (_23350_, _23349_, _03143_);
  nand (_23351_, _09037_, _03143_);
  and (_23352_, _23351_, _22461_);
  and (_23354_, _23352_, _23350_);
  or (_23355_, _23150_, _07288_);
  or (_23356_, _09036_, \oc8051_golden_model_1.PSW [7]);
  and (_23357_, _23356_, _08808_);
  and (_23358_, _23357_, _23355_);
  or (_23359_, _23358_, _09487_);
  nor (_23360_, _23359_, _23354_);
  or (_23361_, _23360_, _07966_);
  nor (_23362_, _23361_, _23124_);
  nor (_23363_, _09037_, _07965_);
  nor (_23365_, _23363_, _07995_);
  not (_23366_, _23365_);
  nor (_23367_, _23366_, _23362_);
  nor (_23368_, _23367_, _23123_);
  nor (_23369_, _23368_, _03155_);
  and (_23370_, _04449_, _03155_);
  nor (_23371_, _23370_, _23054_);
  not (_23372_, _23371_);
  nor (_23373_, _23372_, _23369_);
  not (_23374_, _08803_);
  nor (_23376_, _09692_, _08851_);
  and (_23377_, _23142_, _09692_);
  or (_23378_, _23377_, _03223_);
  nor (_23379_, _23378_, _23376_);
  or (_23380_, _23379_, _23374_);
  nor (_23381_, _23380_, _23373_);
  nor (_23382_, _23122_, _08112_);
  nor (_23383_, _23382_, _21294_);
  nor (_23384_, _23383_, _23381_);
  and (_23385_, _09036_, _08112_);
  nor (_23387_, _23385_, _08115_);
  not (_23388_, _23387_);
  nor (_23389_, _23388_, _23384_);
  and (_23390_, _23122_, _08115_);
  nor (_23391_, _23390_, _23389_);
  nor (_23392_, _23391_, _02890_);
  and (_23393_, _04449_, _02890_);
  nor (_23394_, _23393_, _23075_);
  not (_23395_, _23394_);
  nor (_23396_, _23395_, _23392_);
  and (_23398_, _09692_, _08852_);
  nor (_23399_, _23141_, _09692_);
  nor (_23400_, _23399_, _23398_);
  and (_23401_, _23400_, _02889_);
  nor (_23402_, _23401_, _09725_);
  not (_23403_, _23402_);
  nor (_23404_, _23403_, _23396_);
  nor (_23405_, _23404_, _23121_);
  nor (_23406_, _23405_, _03174_);
  and (_23407_, _09037_, _03174_);
  nor (_23409_, _23407_, _09733_);
  not (_23410_, _23409_);
  nor (_23411_, _23410_, _23406_);
  nor (_23412_, _23122_, _09732_);
  nor (_23413_, _23412_, _03034_);
  not (_23414_, _23413_);
  nor (_23415_, _23414_, _23411_);
  not (_23416_, _22764_);
  and (_23417_, _03356_, _03034_);
  nor (_23418_, _23417_, _23416_);
  not (_23420_, _23418_);
  nor (_23421_, _23420_, _23415_);
  and (_23422_, _23400_, _02799_);
  nor (_23423_, _23422_, _23421_);
  or (_23424_, _23423_, _09748_);
  or (_23425_, _23122_, _09747_);
  and (_23426_, _23425_, _02888_);
  and (_23427_, _23426_, _23424_);
  and (_23428_, _09037_, _02887_);
  nor (_23429_, _23428_, _09756_);
  not (_23430_, _23429_);
  or (_23431_, _23430_, _23427_);
  nor (_23432_, _23122_, _09755_);
  nor (_23433_, _23432_, _03036_);
  nand (_23434_, _23433_, _23431_);
  not (_23435_, _22780_);
  and (_23436_, _03356_, _03036_);
  nor (_23437_, _23436_, _23435_);
  and (_23438_, _23437_, _23434_);
  or (_23439_, _23438_, _23120_);
  or (_23441_, _23439_, _34659_);
  or (_23442_, _34655_, \oc8051_golden_model_1.PC [10]);
  and (_23443_, _23442_, _35796_);
  and (_35842_[10], _23443_, _23441_);
  nor (_23444_, _08795_, \oc8051_golden_model_1.PC [11]);
  nor (_23445_, _23444_, _08796_);
  or (_23446_, _23445_, _08803_);
  or (_23447_, _23445_, _08806_);
  or (_23448_, _09030_, _08809_);
  and (_23449_, _23448_, _19607_);
  or (_23451_, _23445_, _08815_);
  or (_23452_, _23445_, _09453_);
  or (_23453_, _23445_, _08823_);
  not (_23454_, _09360_);
  nor (_23455_, _23139_, _08853_);
  and (_23456_, _23455_, _08848_);
  nor (_23457_, _23455_, _08848_);
  or (_23458_, _23457_, _23456_);
  and (_23459_, _23458_, _08981_);
  and (_23460_, _09918_, _08844_);
  or (_23462_, _23460_, _08986_);
  or (_23463_, _23462_, _23459_);
  nor (_23464_, _08991_, _09031_);
  or (_23465_, _08994_, _09030_);
  nand (_23466_, _09003_, _08845_);
  or (_23467_, _23458_, _09003_);
  and (_23468_, _23467_, _02948_);
  and (_23469_, _23468_, _23466_);
  nor (_23470_, _23148_, _09038_);
  nor (_23471_, _23470_, _09034_);
  and (_23473_, _23470_, _09034_);
  or (_23474_, _23473_, _23471_);
  and (_23475_, _23474_, _19652_);
  and (_23476_, _09012_, _09030_);
  or (_23477_, _23476_, _05361_);
  or (_23478_, _23477_, _23475_);
  nor (_23479_, _09031_, _02601_);
  or (_23480_, _23445_, _09145_);
  or (_23481_, _09138_, \oc8051_golden_model_1.PC [11]);
  nand (_23482_, _09135_, _04194_);
  or (_23484_, _23482_, _23481_);
  and (_23485_, _23484_, _23480_);
  or (_23486_, _23485_, _03849_);
  nor (_23487_, _03845_, _03849_);
  or (_23488_, _23487_, _09030_);
  and (_23489_, _23488_, _09153_);
  and (_23490_, _23489_, _23486_);
  not (_23491_, _23445_);
  nor (_23492_, _23491_, _09153_);
  or (_23493_, _23492_, _23490_);
  and (_23494_, _23493_, _03401_);
  and (_23495_, _09030_, _02951_);
  or (_23496_, _23495_, _07436_);
  or (_23497_, _23496_, _23494_);
  nand (_23498_, _23491_, _07436_);
  and (_23499_, _23498_, _02601_);
  and (_23500_, _23499_, _23497_);
  or (_23501_, _23500_, _23479_);
  and (_23502_, _23501_, _09133_);
  nand (_23503_, _23445_, _07433_);
  nand (_23505_, _23503_, _05361_);
  or (_23506_, _23505_, _23502_);
  and (_23507_, _23506_, _09176_);
  and (_23508_, _23507_, _23478_);
  or (_23509_, _23508_, _23469_);
  and (_23510_, _23509_, _08997_);
  not (_23511_, _08994_);
  and (_23512_, _23445_, _09181_);
  or (_23513_, _23512_, _23511_);
  or (_23514_, _23513_, _23510_);
  and (_23516_, _23514_, _23465_);
  or (_23517_, _23516_, _09187_);
  or (_23518_, _23445_, _09186_);
  and (_23519_, _23518_, _02992_);
  and (_23520_, _23519_, _23517_);
  and (_23521_, _09030_, _02880_);
  or (_23522_, _23521_, _09193_);
  or (_23523_, _23522_, _23520_);
  nand (_23524_, _23491_, _09193_);
  and (_23525_, _23524_, _08991_);
  and (_23527_, _23525_, _23523_);
  or (_23528_, _23527_, _23464_);
  and (_23529_, _23528_, _09209_);
  nand (_23530_, _09242_, _08845_);
  or (_23531_, _23458_, _09242_);
  and (_23532_, _23531_, _09210_);
  and (_23533_, _23532_, _23530_);
  or (_23534_, _23533_, _08985_);
  or (_23535_, _23534_, _23529_);
  and (_23536_, _23535_, _09251_);
  and (_23538_, _23536_, _23463_);
  or (_23539_, _23458_, _09276_);
  nand (_23540_, _09276_, _08845_);
  and (_23541_, _23540_, _03029_);
  and (_23542_, _23541_, _23539_);
  or (_23543_, _23458_, _09297_);
  nand (_23544_, _09297_, _08845_);
  and (_23545_, _23544_, _02954_);
  and (_23546_, _23545_, _23543_);
  or (_23547_, _23546_, _23542_);
  nand (_23549_, _23445_, _09249_);
  nand (_23550_, _23549_, _09263_);
  or (_23551_, _23550_, _23547_);
  or (_23552_, _23551_, _23538_);
  or (_23553_, _09263_, _09030_);
  and (_23554_, _23553_, _09309_);
  and (_23555_, _23554_, _23552_);
  nor (_23556_, _23491_, _09309_);
  or (_23557_, _23556_, _09317_);
  or (_23558_, _23557_, _23555_);
  or (_23560_, _09316_, _09030_);
  and (_23561_, _23560_, _09320_);
  and (_23562_, _23561_, _23558_);
  nor (_23563_, _23491_, _09320_);
  or (_23564_, _23563_, _09325_);
  or (_23565_, _23564_, _23562_);
  or (_23566_, _09324_, _09030_);
  and (_23567_, _23566_, _02571_);
  and (_23568_, _23567_, _23565_);
  or (_23569_, _23491_, _02571_);
  nand (_23571_, _23569_, _09335_);
  or (_23572_, _23571_, _23568_);
  or (_23573_, _09335_, _09030_);
  and (_23574_, _23573_, _08211_);
  and (_23575_, _23574_, _23572_);
  nand (_23576_, _08844_, _03046_);
  nand (_23577_, _23576_, _02860_);
  or (_23578_, _23577_, _23575_);
  or (_23579_, _09030_, _02860_);
  and (_23580_, _23579_, _02839_);
  and (_23582_, _23580_, _23578_);
  nor (_23583_, _09352_, _08844_);
  nor (_23584_, _23583_, _09353_);
  or (_23585_, _23584_, _23582_);
  nand (_23586_, _23491_, _09352_);
  and (_23587_, _23586_, _23585_);
  or (_23588_, _23587_, _23454_);
  or (_23589_, _09360_, _09030_);
  and (_23590_, _23589_, _09366_);
  and (_23591_, _23590_, _23588_);
  and (_23593_, _23474_, _09362_);
  or (_23594_, _23593_, _05749_);
  or (_23595_, _23594_, _23591_);
  or (_23596_, _09030_, _05748_);
  and (_23597_, _23596_, _07140_);
  and (_23598_, _23597_, _23595_);
  and (_23599_, _08844_, _02834_);
  or (_23600_, _23599_, _07830_);
  or (_23601_, _23600_, _23598_);
  nand (_23602_, _09031_, _07830_);
  and (_23604_, _23602_, _19622_);
  and (_23605_, _23604_, _23601_);
  nor (_23606_, _09406_, \oc8051_golden_model_1.DPH [3]);
  nor (_23607_, _23606_, _09407_);
  and (_23608_, _23607_, _09376_);
  or (_23609_, _23608_, _09416_);
  or (_23610_, _23609_, _23605_);
  or (_23611_, _09415_, _09030_);
  and (_23612_, _23611_, _19621_);
  and (_23613_, _23612_, _23610_);
  or (_23615_, _23474_, _08166_);
  or (_23616_, _09030_, _09447_);
  and (_23617_, _23616_, _09419_);
  and (_23618_, _23617_, _23615_);
  or (_23619_, _23618_, _09428_);
  or (_23620_, _23619_, _23613_);
  and (_23621_, _23620_, _23453_);
  or (_23622_, _23621_, _21199_);
  or (_23623_, _09030_, _08822_);
  and (_23624_, _23623_, _07139_);
  and (_23626_, _23624_, _23622_);
  nand (_23627_, _08844_, _03051_);
  nand (_23628_, _23627_, _09437_);
  or (_23629_, _23628_, _23626_);
  or (_23630_, _09437_, _09030_);
  and (_23631_, _23630_, _09446_);
  and (_23632_, _23631_, _23629_);
  or (_23633_, _23474_, _09447_);
  or (_23634_, _09030_, _08166_);
  and (_23635_, _23634_, _09441_);
  and (_23637_, _23635_, _23633_);
  or (_23638_, _23637_, _20129_);
  or (_23639_, _23638_, _23632_);
  and (_23640_, _23639_, _23452_);
  or (_23641_, _23640_, _09456_);
  or (_23642_, _09030_, _09455_);
  and (_23643_, _23642_, _03023_);
  and (_23644_, _23643_, _23641_);
  nand (_23645_, _08844_, _03022_);
  nand (_23646_, _23645_, _08819_);
  or (_23648_, _23646_, _23644_);
  or (_23649_, _09030_, _08819_);
  and (_23650_, _23649_, _09470_);
  and (_23651_, _23650_, _23648_);
  or (_23652_, _23474_, \oc8051_golden_model_1.PSW [7]);
  or (_23653_, _09030_, _07288_);
  and (_23654_, _23653_, _08818_);
  and (_23655_, _23654_, _23652_);
  or (_23656_, _23655_, _09468_);
  or (_23657_, _23656_, _23651_);
  and (_23659_, _23657_, _23451_);
  or (_23660_, _23659_, _13433_);
  or (_23661_, _09030_, _08812_);
  and (_23662_, _23661_, _03043_);
  and (_23663_, _23662_, _23660_);
  nand (_23664_, _08844_, _03042_);
  nand (_23665_, _23664_, _08809_);
  or (_23666_, _23665_, _23663_);
  and (_23667_, _23666_, _23449_);
  or (_23668_, _23474_, _07288_);
  or (_23670_, _09030_, \oc8051_golden_model_1.PSW [7]);
  and (_23671_, _23670_, _08808_);
  and (_23672_, _23671_, _23668_);
  or (_23673_, _23672_, _09487_);
  or (_23674_, _23673_, _23667_);
  and (_23675_, _23674_, _23447_);
  or (_23676_, _23675_, _07966_);
  or (_23677_, _09030_, _07965_);
  and (_23678_, _23677_, _07996_);
  and (_23679_, _23678_, _23676_);
  and (_23681_, _23445_, _07995_);
  or (_23682_, _23681_, _03155_);
  or (_23683_, _23682_, _23679_);
  nand (_23684_, _04275_, _03155_);
  and (_23685_, _23684_, _23683_);
  or (_23686_, _23685_, _02528_);
  nand (_23687_, _09031_, _02528_);
  and (_23688_, _23687_, _03223_);
  and (_23689_, _23688_, _23686_);
  not (_23690_, _09692_);
  or (_23692_, _23458_, _23690_);
  or (_23693_, _09692_, _08844_);
  and (_23694_, _23693_, _03040_);
  and (_23695_, _23694_, _23692_);
  or (_23696_, _23695_, _23374_);
  or (_23697_, _23696_, _23689_);
  and (_23698_, _23697_, _23446_);
  or (_23699_, _23698_, _08112_);
  nand (_23700_, _09031_, _08112_);
  and (_23701_, _23700_, _08116_);
  and (_23703_, _23701_, _23699_);
  and (_23704_, _23445_, _08115_);
  or (_23705_, _23704_, _02890_);
  or (_23706_, _23705_, _23703_);
  nand (_23707_, _04275_, _02890_);
  and (_23708_, _23707_, _23706_);
  or (_23709_, _23708_, _02510_);
  nand (_23710_, _09031_, _02510_);
  and (_23711_, _23710_, _03175_);
  and (_23712_, _23711_, _23709_);
  or (_23714_, _23458_, _09692_);
  nand (_23715_, _09692_, _08845_);
  and (_23716_, _23715_, _23714_);
  and (_23717_, _23716_, _02889_);
  or (_23718_, _23717_, _09725_);
  or (_23719_, _23718_, _23712_);
  or (_23720_, _23445_, _09724_);
  and (_23721_, _23720_, _03179_);
  and (_23722_, _23721_, _23719_);
  nand (_23723_, _09030_, _03174_);
  nand (_23725_, _23723_, _09732_);
  or (_23726_, _23725_, _23722_);
  or (_23727_, _23445_, _09732_);
  and (_23728_, _23727_, _06185_);
  and (_23729_, _23728_, _23726_);
  and (_23730_, _03034_, _02794_);
  or (_23731_, _23730_, _02505_);
  or (_23732_, _23731_, _23729_);
  nand (_23733_, _09031_, _02505_);
  and (_23734_, _23733_, _03183_);
  and (_23736_, _23734_, _23732_);
  and (_23737_, _23716_, _02799_);
  or (_23738_, _23737_, _09748_);
  or (_23739_, _23738_, _23736_);
  or (_23740_, _23445_, _09747_);
  and (_23741_, _23740_, _02888_);
  and (_23742_, _23741_, _23739_);
  nand (_23743_, _09030_, _02887_);
  nand (_23744_, _23743_, _09755_);
  or (_23745_, _23744_, _23742_);
  or (_23747_, _23445_, _09755_);
  and (_23748_, _23747_, _03038_);
  and (_23749_, _23748_, _23745_);
  and (_23750_, _03036_, _02794_);
  or (_23751_, _23750_, _02499_);
  or (_23752_, _23751_, _23749_);
  nand (_23753_, _09031_, _02499_);
  and (_23754_, _23753_, _08787_);
  and (_23755_, _23754_, _23752_);
  and (_23756_, _23445_, _08786_);
  or (_23758_, _23756_, _23755_);
  or (_23759_, _23758_, _34659_);
  or (_23760_, _34655_, \oc8051_golden_model_1.PC [11]);
  and (_23761_, _23760_, _35796_);
  and (_35842_[11], _23761_, _23759_);
  and (_23762_, _09026_, _02499_);
  nand (_23763_, _09027_, _02887_);
  nor (_23764_, _09027_, _07965_);
  nor (_23765_, _09415_, _09027_);
  and (_23766_, _08841_, _02567_);
  nor (_23768_, _23766_, _09352_);
  nor (_23769_, _08936_, _08934_);
  nor (_23770_, _23769_, _08937_);
  and (_23771_, _23770_, _08981_);
  and (_23772_, _09918_, _08840_);
  or (_23773_, _23772_, _23771_);
  and (_23774_, _23773_, _08985_);
  nor (_23775_, _08796_, \oc8051_golden_model_1.PC [12]);
  nor (_23776_, _23775_, _08797_);
  and (_23777_, _23776_, _09193_);
  or (_23779_, _23776_, _09186_);
  or (_23780_, _23770_, _09003_);
  nand (_23781_, _09003_, _08841_);
  and (_23782_, _23781_, _23780_);
  or (_23783_, _23782_, _03006_);
  nor (_23784_, _09114_, _09112_);
  nor (_23785_, _23784_, _09115_);
  and (_23786_, _23785_, _19652_);
  and (_23787_, _09012_, _09026_);
  or (_23788_, _23787_, _05361_);
  or (_23790_, _23788_, _23786_);
  not (_23791_, _23776_);
  nor (_23792_, _23791_, _09153_);
  nor (_23793_, _23791_, _09145_);
  not (_23794_, \oc8051_golden_model_1.PC [12]);
  nor (_23795_, _03845_, _23794_);
  and (_23796_, _23795_, _09135_);
  and (_23797_, _23796_, _09144_);
  and (_23798_, _23797_, _09153_);
  or (_23799_, _23798_, _23793_);
  and (_23801_, _23799_, _02603_);
  or (_23802_, _23801_, _23792_);
  and (_23803_, _23802_, _03401_);
  nand (_23804_, _23487_, _03401_);
  and (_23805_, _23804_, _09026_);
  or (_23806_, _23805_, _23803_);
  and (_23807_, _23806_, _19632_);
  and (_23808_, _23776_, _07436_);
  or (_23809_, _23808_, _09169_);
  or (_23810_, _23809_, _23807_);
  nor (_23812_, _09026_, _02601_);
  nor (_23813_, _23812_, _07433_);
  and (_23814_, _23813_, _23810_);
  nand (_23815_, _23776_, _07433_);
  nand (_23816_, _23815_, _05361_);
  or (_23817_, _23816_, _23814_);
  and (_23818_, _23817_, _05371_);
  and (_23819_, _23818_, _23790_);
  and (_23820_, _23776_, _03840_);
  or (_23821_, _23820_, _02948_);
  or (_23823_, _23821_, _23819_);
  and (_23824_, _23823_, _23783_);
  or (_23825_, _23824_, _08998_);
  or (_23826_, _23776_, _08997_);
  and (_23827_, _23826_, _08994_);
  and (_23828_, _23827_, _23825_);
  or (_23829_, _08994_, _09027_);
  nand (_23830_, _23829_, _09186_);
  or (_23831_, _23830_, _23828_);
  and (_23832_, _23831_, _23779_);
  or (_23834_, _23832_, _02880_);
  and (_23835_, _09027_, _02880_);
  nor (_23836_, _23835_, _09193_);
  and (_23837_, _23836_, _23834_);
  or (_23838_, _23837_, _23777_);
  and (_23839_, _23838_, _08991_);
  or (_23840_, _08991_, _09027_);
  nand (_23841_, _23840_, _09209_);
  or (_23842_, _23841_, _23839_);
  or (_23843_, _23770_, _09242_);
  nand (_23845_, _09242_, _08841_);
  and (_23846_, _23845_, _23843_);
  or (_23847_, _23846_, _09209_);
  and (_23848_, _23847_, _08986_);
  and (_23849_, _23848_, _23842_);
  or (_23850_, _23849_, _02954_);
  or (_23851_, _23850_, _23774_);
  not (_23852_, _09297_);
  and (_23853_, _23770_, _23852_);
  and (_23854_, _09297_, _08840_);
  or (_23856_, _23854_, _09299_);
  or (_23857_, _23856_, _23853_);
  and (_23858_, _23857_, _09279_);
  and (_23859_, _23858_, _23851_);
  or (_23860_, _23770_, _09276_);
  nand (_23861_, _09276_, _08841_);
  and (_23862_, _23861_, _03029_);
  and (_23863_, _23862_, _23860_);
  or (_23864_, _23863_, _09249_);
  or (_23865_, _23864_, _23859_);
  nand (_23867_, _23791_, _09249_);
  and (_23868_, _23867_, _09263_);
  and (_23869_, _23868_, _23865_);
  nor (_23870_, _09263_, _09027_);
  or (_23871_, _23870_, _09310_);
  or (_23872_, _23871_, _23869_);
  or (_23873_, _23776_, _09309_);
  and (_23874_, _23873_, _09316_);
  and (_23875_, _23874_, _23872_);
  nor (_23876_, _09316_, _09027_);
  or (_23878_, _23876_, _09326_);
  or (_23879_, _23878_, _23875_);
  or (_23880_, _23776_, _09320_);
  and (_23881_, _23880_, _09324_);
  and (_23882_, _23881_, _23879_);
  nor (_23883_, _09324_, _09027_);
  or (_23884_, _23883_, _07721_);
  or (_23885_, _23884_, _23882_);
  and (_23886_, _23776_, _09335_);
  or (_23887_, _23886_, _09336_);
  and (_23889_, _23887_, _23885_);
  nor (_23890_, _09335_, _09027_);
  or (_23891_, _23890_, _03046_);
  or (_23892_, _23891_, _23889_);
  nand (_23893_, _08841_, _03046_);
  and (_23894_, _23893_, _02860_);
  and (_23895_, _23894_, _23892_);
  nor (_23896_, _09027_, _02860_);
  or (_23897_, _23896_, _02567_);
  or (_23898_, _23897_, _23895_);
  and (_23900_, _23898_, _23768_);
  and (_23901_, _23776_, _09352_);
  or (_23902_, _23901_, _23454_);
  or (_23903_, _23902_, _23900_);
  or (_23904_, _09360_, _09026_);
  and (_23905_, _23904_, _09366_);
  and (_23906_, _23905_, _23903_);
  and (_23907_, _23785_, _09362_);
  or (_23908_, _23907_, _23906_);
  and (_23909_, _23908_, _05748_);
  nor (_23911_, _09027_, _05748_);
  or (_23912_, _23911_, _02834_);
  or (_23913_, _23912_, _23909_);
  nand (_23914_, _08841_, _02834_);
  and (_23915_, _23914_, _07831_);
  and (_23916_, _23915_, _23913_);
  and (_23917_, _09026_, _07830_);
  or (_23918_, _23917_, _09376_);
  or (_23919_, _23918_, _23916_);
  nor (_23920_, _09407_, \oc8051_golden_model_1.DPH [4]);
  nor (_23922_, _23920_, _09408_);
  or (_23923_, _23922_, _19622_);
  and (_23924_, _23923_, _09415_);
  and (_23925_, _23924_, _23919_);
  or (_23926_, _23925_, _23765_);
  and (_23927_, _23926_, _21190_);
  or (_23928_, _23785_, _08166_);
  or (_23929_, _09026_, _09447_);
  and (_23930_, _23929_, _09419_);
  and (_23931_, _23930_, _23928_);
  nor (_23933_, _23791_, _08823_);
  or (_23934_, _23933_, _23931_);
  or (_23935_, _23934_, _23927_);
  and (_23936_, _23935_, _08822_);
  nor (_23937_, _09027_, _08822_);
  or (_23938_, _23937_, _03051_);
  or (_23939_, _23938_, _23936_);
  nand (_23940_, _08841_, _03051_);
  and (_23941_, _23940_, _09437_);
  and (_23942_, _23941_, _23939_);
  nor (_23944_, _09437_, _09027_);
  or (_23945_, _23944_, _23942_);
  and (_23946_, _23945_, _21214_);
  nor (_23947_, _23791_, _09453_);
  or (_23948_, _23785_, _09447_);
  or (_23949_, _09026_, _08166_);
  and (_23950_, _23949_, _09441_);
  and (_23951_, _23950_, _23948_);
  or (_23952_, _23951_, _23947_);
  or (_23953_, _23952_, _23946_);
  and (_23955_, _23953_, _09455_);
  nor (_23956_, _09027_, _09455_);
  or (_23957_, _23956_, _03022_);
  or (_23958_, _23957_, _23955_);
  nand (_23959_, _08841_, _03022_);
  and (_23960_, _23959_, _08819_);
  and (_23961_, _23960_, _23958_);
  nor (_23962_, _09027_, _08819_);
  or (_23963_, _23962_, _23961_);
  and (_23964_, _23963_, _21747_);
  nor (_23966_, _23791_, _08815_);
  or (_23967_, _23785_, \oc8051_golden_model_1.PSW [7]);
  or (_23968_, _09026_, _07288_);
  and (_23969_, _23968_, _08818_);
  and (_23970_, _23969_, _23967_);
  or (_23971_, _23970_, _23966_);
  or (_23972_, _23971_, _23964_);
  and (_23973_, _23972_, _08812_);
  nor (_23974_, _09027_, _08812_);
  or (_23975_, _23974_, _03042_);
  or (_23977_, _23975_, _23973_);
  nand (_23978_, _08841_, _03042_);
  and (_23979_, _23978_, _08809_);
  and (_23980_, _23979_, _23977_);
  nor (_23981_, _09027_, _08809_);
  or (_23982_, _23981_, _23980_);
  and (_23983_, _23982_, _21260_);
  nor (_23984_, _23791_, _08806_);
  or (_23985_, _23785_, _07288_);
  or (_23986_, _09026_, \oc8051_golden_model_1.PSW [7]);
  and (_23988_, _23986_, _08808_);
  and (_23989_, _23988_, _23985_);
  or (_23990_, _23989_, _23984_);
  or (_23991_, _23990_, _23983_);
  and (_23992_, _23991_, _07965_);
  or (_23993_, _23992_, _23764_);
  and (_23994_, _23993_, _07996_);
  and (_23995_, _23776_, _07995_);
  or (_23996_, _23995_, _03155_);
  or (_23997_, _23996_, _23994_);
  nand (_23999_, _05192_, _03155_);
  and (_24000_, _23999_, _23997_);
  or (_24001_, _24000_, _02528_);
  nand (_24002_, _09027_, _02528_);
  and (_24003_, _24002_, _03223_);
  and (_24004_, _24003_, _24001_);
  or (_24005_, _09692_, _08840_);
  or (_24006_, _23770_, _23690_);
  and (_24007_, _24006_, _03040_);
  and (_24008_, _24007_, _24005_);
  or (_24010_, _24008_, _23374_);
  or (_24011_, _24010_, _24004_);
  nor (_24012_, _23791_, _08112_);
  or (_24013_, _24012_, _21294_);
  and (_24014_, _24013_, _24011_);
  and (_24015_, _09026_, _08112_);
  or (_24016_, _24015_, _08115_);
  or (_24017_, _24016_, _24014_);
  nand (_24018_, _23791_, _08115_);
  and (_24019_, _24018_, _24017_);
  or (_24021_, _24019_, _02890_);
  nand (_24022_, _05192_, _02890_);
  and (_24023_, _24022_, _08788_);
  and (_24024_, _24023_, _24021_);
  and (_24025_, _09026_, _02510_);
  or (_24026_, _24025_, _02889_);
  or (_24027_, _24026_, _24024_);
  nand (_24028_, _09692_, _08841_);
  or (_24029_, _23770_, _09692_);
  and (_24030_, _24029_, _24028_);
  or (_24032_, _24030_, _03175_);
  and (_24033_, _24032_, _24027_);
  or (_24034_, _24033_, _09725_);
  or (_24035_, _23776_, _09724_);
  and (_24036_, _24035_, _24034_);
  or (_24037_, _24036_, _03174_);
  nand (_24038_, _09027_, _03174_);
  and (_24039_, _24038_, _09732_);
  and (_24040_, _24039_, _24037_);
  nor (_24041_, _23791_, _09732_);
  or (_24043_, _24041_, _03034_);
  or (_24044_, _24043_, _24040_);
  nand (_24045_, _03647_, _03034_);
  and (_24046_, _24045_, _09742_);
  and (_24047_, _24046_, _24044_);
  and (_24048_, _09026_, _02505_);
  or (_24049_, _24048_, _02799_);
  or (_24050_, _24049_, _24047_);
  or (_24051_, _24030_, _03183_);
  and (_24052_, _24051_, _09747_);
  and (_24054_, _24052_, _24050_);
  nor (_24055_, _23791_, _09747_);
  or (_24056_, _24055_, _02887_);
  or (_24057_, _24056_, _24054_);
  and (_24058_, _24057_, _23763_);
  or (_24059_, _24058_, _09756_);
  or (_24060_, _23776_, _09755_);
  and (_24061_, _24060_, _03038_);
  and (_24062_, _24061_, _24059_);
  nor (_24063_, _03647_, _03038_);
  nor (_24065_, _24063_, _24062_);
  nor (_24066_, _24065_, _02499_);
  nor (_24067_, _24066_, _23762_);
  nor (_24068_, _24067_, _08786_);
  and (_24069_, _23776_, _08786_);
  nor (_24070_, _24069_, _24068_);
  nand (_24071_, _24070_, _34655_);
  or (_24072_, _34655_, \oc8051_golden_model_1.PC [12]);
  and (_24073_, _24072_, _35796_);
  and (_35842_[12], _24073_, _24071_);
  nor (_24076_, _08797_, \oc8051_golden_model_1.PC [13]);
  nor (_24077_, _24076_, _08798_);
  or (_24078_, _24077_, _08803_);
  or (_24079_, _24077_, _08806_);
  or (_24080_, _09021_, _08809_);
  and (_24081_, _24080_, _19607_);
  or (_24082_, _24077_, _08815_);
  or (_24083_, _09021_, _08819_);
  and (_24084_, _24083_, _09470_);
  or (_24085_, _24077_, _08823_);
  or (_24088_, _08837_, _08836_);
  nand (_24089_, _24088_, _08938_);
  or (_24090_, _24088_, _08938_);
  and (_24091_, _24090_, _24089_);
  and (_24092_, _24091_, _08981_);
  and (_24093_, _09918_, _08834_);
  or (_24094_, _24093_, _24092_);
  or (_24095_, _24094_, _08986_);
  nor (_24096_, _08991_, _09022_);
  or (_24097_, _08994_, _09021_);
  nand (_24100_, _09003_, _08835_);
  or (_24101_, _24091_, _09003_);
  and (_24102_, _24101_, _02948_);
  and (_24103_, _24102_, _24100_);
  or (_24104_, _09024_, _09023_);
  nand (_24105_, _24104_, _09116_);
  or (_24106_, _24104_, _09116_);
  and (_24107_, _24106_, _24105_);
  and (_24108_, _24107_, _19652_);
  and (_24109_, _09012_, _09021_);
  or (_24112_, _24109_, _05361_);
  or (_24113_, _24112_, _24108_);
  and (_24114_, _09021_, _09169_);
  or (_24115_, _24077_, _22497_);
  or (_24116_, _23487_, _09021_);
  or (_24117_, _03849_, \oc8051_golden_model_1.PC [13]);
  or (_24118_, _24117_, _09138_);
  or (_24119_, _24118_, _23482_);
  and (_24120_, _24119_, _24116_);
  or (_24121_, _24120_, _09154_);
  and (_24124_, _24121_, _03401_);
  and (_24125_, _24124_, _24115_);
  and (_24126_, _09021_, _02951_);
  or (_24127_, _24126_, _07436_);
  or (_24128_, _24127_, _24125_);
  not (_24129_, _24077_);
  nand (_24130_, _24129_, _07436_);
  and (_24131_, _24130_, _02601_);
  and (_24132_, _24131_, _24128_);
  or (_24133_, _24132_, _24114_);
  and (_24136_, _24133_, _09133_);
  nand (_24137_, _24077_, _07433_);
  nand (_24138_, _24137_, _05361_);
  or (_24139_, _24138_, _24136_);
  and (_24140_, _24139_, _09176_);
  and (_24141_, _24140_, _24113_);
  or (_24142_, _24141_, _24103_);
  and (_24143_, _24142_, _08997_);
  and (_24144_, _24077_, _09181_);
  or (_24145_, _24144_, _23511_);
  or (_24148_, _24145_, _24143_);
  and (_24149_, _24148_, _24097_);
  or (_24150_, _24149_, _09187_);
  or (_24151_, _24077_, _09186_);
  and (_24152_, _24151_, _02992_);
  and (_24153_, _24152_, _24150_);
  and (_24154_, _09021_, _02880_);
  or (_24155_, _24154_, _09193_);
  or (_24156_, _24155_, _24153_);
  nand (_24157_, _24129_, _09193_);
  and (_24159_, _24157_, _08991_);
  and (_24160_, _24159_, _24156_);
  or (_24161_, _24160_, _24096_);
  and (_24162_, _24161_, _09209_);
  nand (_24163_, _09242_, _08835_);
  or (_24164_, _24091_, _09242_);
  and (_24165_, _24164_, _09210_);
  and (_24166_, _24165_, _24163_);
  or (_24167_, _24166_, _08985_);
  or (_24168_, _24167_, _24162_);
  and (_24170_, _24168_, _09251_);
  and (_24171_, _24170_, _24095_);
  or (_24172_, _24091_, _09276_);
  nand (_24173_, _09276_, _08835_);
  and (_24174_, _24173_, _03029_);
  and (_24175_, _24174_, _24172_);
  or (_24176_, _24091_, _09297_);
  nand (_24177_, _09297_, _08835_);
  and (_24178_, _24177_, _02954_);
  and (_24179_, _24178_, _24176_);
  or (_24181_, _24179_, _24175_);
  nand (_24182_, _24077_, _09249_);
  nand (_24183_, _24182_, _09263_);
  or (_24184_, _24183_, _24181_);
  or (_24185_, _24184_, _24171_);
  or (_24186_, _09263_, _09021_);
  and (_24187_, _24186_, _09309_);
  and (_24188_, _24187_, _24185_);
  nor (_24189_, _24129_, _09309_);
  or (_24190_, _24189_, _09317_);
  or (_24192_, _24190_, _24188_);
  or (_24193_, _09316_, _09021_);
  and (_24194_, _24193_, _09320_);
  and (_24195_, _24194_, _24192_);
  nor (_24196_, _24129_, _09320_);
  or (_24197_, _24196_, _09325_);
  or (_24198_, _24197_, _24195_);
  or (_24199_, _09324_, _09021_);
  and (_24200_, _24199_, _02571_);
  and (_24201_, _24200_, _24198_);
  nand (_24203_, _24077_, _07721_);
  nand (_24204_, _24203_, _09335_);
  or (_24205_, _24204_, _24201_);
  or (_24206_, _09335_, _09021_);
  and (_24207_, _24206_, _08211_);
  and (_24208_, _24207_, _24205_);
  nand (_24209_, _08834_, _03046_);
  nand (_24210_, _24209_, _02860_);
  or (_24211_, _24210_, _24208_);
  or (_24212_, _09021_, _02860_);
  and (_24214_, _24212_, _02839_);
  and (_24215_, _24214_, _24211_);
  nor (_24216_, _09352_, _08834_);
  nor (_24217_, _24216_, _09353_);
  or (_24218_, _24217_, _24215_);
  nand (_24219_, _24129_, _09352_);
  and (_24220_, _24219_, _24218_);
  or (_24221_, _24220_, _23454_);
  or (_24222_, _09360_, _09021_);
  and (_24223_, _24222_, _09366_);
  and (_24225_, _24223_, _24221_);
  and (_24226_, _24107_, _09362_);
  or (_24227_, _24226_, _05749_);
  or (_24228_, _24227_, _24225_);
  or (_24229_, _09021_, _05748_);
  and (_24230_, _24229_, _07140_);
  and (_24231_, _24230_, _24228_);
  and (_24232_, _08834_, _02834_);
  or (_24233_, _24232_, _07830_);
  or (_24234_, _24233_, _24231_);
  nand (_24236_, _09022_, _07830_);
  and (_24237_, _24236_, _19622_);
  and (_24238_, _24237_, _24234_);
  nor (_24239_, _09408_, \oc8051_golden_model_1.DPH [5]);
  nor (_24240_, _24239_, _09409_);
  and (_24241_, _24240_, _09376_);
  or (_24242_, _24241_, _09416_);
  or (_24243_, _24242_, _24238_);
  or (_24244_, _09415_, _09021_);
  and (_24245_, _24244_, _19621_);
  and (_24247_, _24245_, _24243_);
  or (_24248_, _24107_, _08166_);
  or (_24249_, _09021_, _09447_);
  and (_24250_, _24249_, _09419_);
  and (_24251_, _24250_, _24248_);
  or (_24252_, _24251_, _09428_);
  or (_24253_, _24252_, _24247_);
  and (_24254_, _24253_, _24085_);
  or (_24255_, _24254_, _21199_);
  or (_24256_, _09021_, _08822_);
  and (_24258_, _24256_, _07139_);
  and (_24259_, _24258_, _24255_);
  nand (_24260_, _08834_, _03051_);
  nand (_24261_, _24260_, _09437_);
  or (_24262_, _24261_, _24259_);
  or (_24263_, _09437_, _09021_);
  and (_24264_, _24263_, _09446_);
  and (_24265_, _24264_, _24262_);
  or (_24266_, _24107_, _09447_);
  or (_24267_, _09021_, _08166_);
  and (_24269_, _24267_, _09441_);
  and (_24270_, _24269_, _24266_);
  or (_24271_, _24270_, _24265_);
  and (_24272_, _24271_, _09453_);
  nor (_24273_, _24129_, _09453_);
  or (_24274_, _24273_, _09456_);
  or (_24275_, _24274_, _24272_);
  or (_24276_, _09021_, _09455_);
  and (_24277_, _24276_, _03023_);
  and (_24278_, _24277_, _24275_);
  nand (_24280_, _08834_, _03022_);
  nand (_24281_, _24280_, _08819_);
  or (_24282_, _24281_, _24278_);
  and (_24283_, _24282_, _24084_);
  or (_24284_, _24107_, \oc8051_golden_model_1.PSW [7]);
  or (_24285_, _09021_, _07288_);
  and (_24286_, _24285_, _08818_);
  and (_24287_, _24286_, _24284_);
  or (_24288_, _24287_, _09468_);
  or (_24289_, _24288_, _24283_);
  and (_24291_, _24289_, _24082_);
  or (_24292_, _24291_, _13433_);
  or (_24293_, _09021_, _08812_);
  and (_24294_, _24293_, _03043_);
  and (_24295_, _24294_, _24292_);
  nand (_24296_, _08834_, _03042_);
  nand (_24297_, _24296_, _08809_);
  or (_24298_, _24297_, _24295_);
  and (_24299_, _24298_, _24081_);
  or (_24300_, _24107_, _07288_);
  or (_24302_, _09021_, \oc8051_golden_model_1.PSW [7]);
  and (_24303_, _24302_, _08808_);
  and (_24304_, _24303_, _24300_);
  or (_24305_, _24304_, _09487_);
  or (_24306_, _24305_, _24299_);
  and (_24307_, _24306_, _24079_);
  or (_24308_, _24307_, _07966_);
  or (_24309_, _09021_, _07965_);
  and (_24310_, _24309_, _07996_);
  and (_24311_, _24310_, _24308_);
  and (_24313_, _24077_, _07995_);
  or (_24314_, _24313_, _03155_);
  or (_24315_, _24314_, _24311_);
  nand (_24316_, _04894_, _03155_);
  and (_24317_, _24316_, _24315_);
  or (_24318_, _24317_, _02528_);
  nand (_24319_, _09022_, _02528_);
  and (_24320_, _24319_, _03223_);
  and (_24321_, _24320_, _24318_);
  or (_24322_, _24091_, _23690_);
  or (_24324_, _09692_, _08834_);
  and (_24325_, _24324_, _03040_);
  and (_24326_, _24325_, _24322_);
  or (_24327_, _24326_, _23374_);
  or (_24328_, _24327_, _24321_);
  and (_24329_, _24328_, _24078_);
  or (_24330_, _24329_, _08112_);
  nand (_24331_, _09022_, _08112_);
  and (_24332_, _24331_, _08116_);
  and (_24333_, _24332_, _24330_);
  and (_24335_, _24077_, _08115_);
  or (_24336_, _24335_, _02890_);
  or (_24337_, _24336_, _24333_);
  nand (_24338_, _04894_, _02890_);
  and (_24339_, _24338_, _24337_);
  or (_24340_, _24339_, _02510_);
  nand (_24341_, _09022_, _02510_);
  and (_24342_, _24341_, _03175_);
  and (_24343_, _24342_, _24340_);
  or (_24344_, _24091_, _09692_);
  nand (_24346_, _09692_, _08835_);
  and (_24347_, _24346_, _24344_);
  and (_24348_, _24347_, _02889_);
  or (_24349_, _24348_, _09725_);
  or (_24350_, _24349_, _24343_);
  or (_24351_, _24077_, _09724_);
  and (_24352_, _24351_, _03179_);
  and (_24353_, _24352_, _24350_);
  nand (_24354_, _09021_, _03174_);
  nand (_24355_, _24354_, _09732_);
  or (_24357_, _24355_, _24353_);
  or (_24358_, _24077_, _09732_);
  and (_24359_, _24358_, _06185_);
  and (_24360_, _24359_, _24357_);
  nor (_24361_, _03220_, _06185_);
  or (_24362_, _24361_, _02505_);
  or (_24363_, _24362_, _24360_);
  nand (_24364_, _09022_, _02505_);
  and (_24365_, _24364_, _03183_);
  and (_24366_, _24365_, _24363_);
  and (_24368_, _24347_, _02799_);
  or (_24369_, _24368_, _09748_);
  or (_24370_, _24369_, _24366_);
  or (_24371_, _24077_, _09747_);
  and (_24372_, _24371_, _02888_);
  and (_24373_, _24372_, _24370_);
  nand (_24374_, _09021_, _02887_);
  nand (_24375_, _24374_, _09755_);
  or (_24376_, _24375_, _24373_);
  or (_24377_, _24077_, _09755_);
  and (_24379_, _24377_, _03038_);
  and (_24380_, _24379_, _24376_);
  nor (_24381_, _03220_, _03038_);
  or (_24382_, _24381_, _02499_);
  or (_24383_, _24382_, _24380_);
  nand (_24384_, _09022_, _02499_);
  and (_24385_, _24384_, _08787_);
  and (_24386_, _24385_, _24383_);
  and (_24387_, _24077_, _08786_);
  or (_24388_, _24387_, _24386_);
  or (_24390_, _24388_, _34659_);
  or (_24391_, _34655_, \oc8051_golden_model_1.PC [13]);
  and (_24392_, _24391_, _35796_);
  and (_35842_[13], _24392_, _24390_);
  nand (_24393_, _09015_, _02499_);
  nor (_24394_, _09015_, _02888_);
  nor (_24395_, _09016_, _07965_);
  nor (_24396_, _09415_, _09016_);
  or (_24397_, _08826_, _02839_);
  and (_24398_, _24397_, _09357_);
  or (_24400_, _09263_, _09015_);
  and (_24401_, _09242_, _08826_);
  and (_24402_, _08940_, _08832_);
  nor (_24403_, _24402_, _08941_);
  not (_24404_, _24403_);
  nor (_24405_, _24404_, _09242_);
  or (_24406_, _24405_, _24401_);
  or (_24407_, _24406_, _09209_);
  or (_24408_, _09015_, _02992_);
  nor (_24409_, _09119_, _09019_);
  nor (_24411_, _24409_, _09120_);
  and (_24412_, _24411_, _19652_);
  and (_24413_, _09012_, _09015_);
  or (_24414_, _24413_, _24412_);
  or (_24415_, _24414_, _05361_);
  or (_24416_, _23804_, _09169_);
  and (_24417_, _24416_, _09015_);
  nor (_24418_, _08798_, \oc8051_golden_model_1.PC [14]);
  nor (_24419_, _24418_, _08799_);
  nand (_24420_, _22497_, _19632_);
  and (_24422_, _24420_, _24419_);
  or (_24423_, _07436_, _02951_);
  not (_24424_, _24423_);
  nand (_24425_, _02603_, \oc8051_golden_model_1.PC [14]);
  nor (_24426_, _24425_, _03845_);
  and (_24427_, _24426_, _09145_);
  and (_24428_, _24427_, _24424_);
  and (_24429_, _24428_, _09153_);
  or (_24430_, _24429_, _24422_);
  and (_24431_, _24430_, _02601_);
  or (_24433_, _24431_, _24417_);
  and (_24434_, _24433_, _09133_);
  nand (_24435_, _24419_, _07433_);
  nand (_24436_, _24435_, _05361_);
  or (_24437_, _24436_, _24434_);
  and (_24438_, _24437_, _24415_);
  or (_24439_, _24438_, _03840_);
  or (_24440_, _24419_, _05371_);
  and (_24441_, _24440_, _03006_);
  and (_24442_, _24441_, _24439_);
  or (_24444_, _24403_, _09003_);
  and (_24445_, _24444_, _02948_);
  or (_24446_, _22852_, _08826_);
  and (_24447_, _24446_, _24445_);
  or (_24448_, _24447_, _08998_);
  or (_24449_, _24448_, _24442_);
  or (_24450_, _24419_, _08997_);
  and (_24451_, _24450_, _24449_);
  or (_24452_, _24451_, _23511_);
  or (_24453_, _08994_, _09015_);
  and (_24455_, _24453_, _09186_);
  and (_24456_, _24455_, _24452_);
  not (_24457_, _24419_);
  nor (_24458_, _24457_, _09186_);
  or (_24459_, _24458_, _02880_);
  or (_24460_, _24459_, _24456_);
  and (_24461_, _24460_, _24408_);
  or (_24462_, _24461_, _09193_);
  or (_24463_, _24419_, _09200_);
  and (_24464_, _24463_, _08991_);
  and (_24466_, _24464_, _24462_);
  or (_24467_, _08991_, _09016_);
  nand (_24468_, _24467_, _09209_);
  or (_24469_, _24468_, _24466_);
  and (_24470_, _24469_, _24407_);
  or (_24471_, _24470_, _08985_);
  and (_24472_, _09918_, _08826_);
  and (_24473_, _24403_, _08981_);
  or (_24474_, _24473_, _24472_);
  or (_24475_, _24474_, _08986_);
  and (_24477_, _24475_, _24471_);
  and (_24478_, _24477_, _09251_);
  or (_24479_, _24403_, _09276_);
  nand (_24480_, _09276_, _08828_);
  and (_24481_, _24480_, _03029_);
  and (_24482_, _24481_, _24479_);
  nand (_24483_, _09297_, _08828_);
  or (_24484_, _24403_, _09297_);
  and (_24485_, _24484_, _02954_);
  and (_24486_, _24485_, _24483_);
  or (_24488_, _24486_, _24482_);
  nand (_24489_, _24419_, _09249_);
  nand (_24490_, _24489_, _09263_);
  or (_24491_, _24490_, _24488_);
  or (_24492_, _24491_, _24478_);
  and (_24493_, _24492_, _24400_);
  or (_24494_, _24493_, _09310_);
  or (_24495_, _24419_, _09309_);
  and (_24496_, _24495_, _09316_);
  and (_24497_, _24496_, _24494_);
  nor (_24499_, _09316_, _09016_);
  or (_24500_, _24499_, _09326_);
  or (_24501_, _24500_, _24497_);
  or (_24502_, _24419_, _09320_);
  and (_24503_, _24502_, _09324_);
  and (_24504_, _24503_, _24501_);
  nor (_24505_, _09324_, _09016_);
  or (_24506_, _24505_, _07721_);
  or (_24507_, _24506_, _24504_);
  or (_24508_, _24419_, _02571_);
  and (_24511_, _24508_, _09335_);
  and (_24512_, _24511_, _24507_);
  nor (_24513_, _09335_, _09016_);
  or (_24514_, _24513_, _03046_);
  or (_24515_, _24514_, _24512_);
  or (_24516_, _08826_, _08211_);
  and (_24517_, _24516_, _02860_);
  and (_24518_, _24517_, _24515_);
  nor (_24519_, _09016_, _02860_);
  or (_24520_, _24519_, _02567_);
  or (_24522_, _24520_, _24518_);
  and (_24523_, _24522_, _24398_);
  and (_24524_, _24419_, _09352_);
  or (_24525_, _24524_, _23454_);
  or (_24526_, _24525_, _24523_);
  or (_24527_, _09360_, _09015_);
  and (_24528_, _24527_, _09366_);
  and (_24529_, _24528_, _24526_);
  and (_24530_, _24411_, _09362_);
  or (_24531_, _24530_, _05749_);
  or (_24533_, _24531_, _24529_);
  or (_24534_, _09015_, _05748_);
  and (_24535_, _24534_, _24533_);
  or (_24536_, _24535_, _02834_);
  or (_24537_, _08826_, _07140_);
  and (_24538_, _24537_, _07831_);
  and (_24539_, _24538_, _24536_);
  and (_24540_, _09015_, _07830_);
  or (_24541_, _24540_, _09376_);
  or (_24542_, _24541_, _24539_);
  nor (_24544_, _09409_, \oc8051_golden_model_1.DPH [6]);
  nor (_24545_, _24544_, _09410_);
  or (_24546_, _24545_, _19622_);
  and (_24547_, _24546_, _09415_);
  and (_24548_, _24547_, _24542_);
  or (_24549_, _24548_, _24396_);
  and (_24550_, _24549_, _21190_);
  or (_24551_, _24411_, _08166_);
  or (_24552_, _09015_, _09447_);
  and (_24553_, _24552_, _09419_);
  and (_24555_, _24553_, _24551_);
  nor (_24556_, _24457_, _08823_);
  or (_24557_, _24556_, _24555_);
  or (_24558_, _24557_, _24550_);
  and (_24559_, _24558_, _08822_);
  nor (_24560_, _09016_, _08822_);
  or (_24561_, _24560_, _03051_);
  or (_24562_, _24561_, _24559_);
  or (_24563_, _08826_, _07139_);
  and (_24564_, _24563_, _09437_);
  and (_24566_, _24564_, _24562_);
  nor (_24567_, _09437_, _09016_);
  or (_24568_, _24567_, _24566_);
  and (_24569_, _24568_, _21214_);
  nor (_24570_, _24457_, _09453_);
  or (_24571_, _24411_, _09447_);
  or (_24572_, _09015_, _08166_);
  and (_24573_, _24572_, _09441_);
  and (_24574_, _24573_, _24571_);
  or (_24575_, _24574_, _24570_);
  or (_24577_, _24575_, _24569_);
  and (_24578_, _24577_, _09455_);
  nor (_24579_, _09016_, _09455_);
  or (_24580_, _24579_, _03022_);
  or (_24581_, _24580_, _24578_);
  or (_24582_, _08826_, _03023_);
  and (_24583_, _24582_, _08819_);
  and (_24584_, _24583_, _24581_);
  nor (_24585_, _09016_, _08819_);
  or (_24586_, _24585_, _24584_);
  and (_24588_, _24586_, _21747_);
  nor (_24589_, _24457_, _08815_);
  or (_24590_, _24411_, \oc8051_golden_model_1.PSW [7]);
  or (_24591_, _09015_, _07288_);
  and (_24592_, _24591_, _08818_);
  and (_24593_, _24592_, _24590_);
  or (_24594_, _24593_, _24589_);
  or (_24595_, _24594_, _24588_);
  and (_24596_, _24595_, _08812_);
  nor (_24597_, _09016_, _08812_);
  or (_24599_, _24597_, _03042_);
  or (_24600_, _24599_, _24596_);
  or (_24601_, _08826_, _03043_);
  and (_24602_, _24601_, _08809_);
  and (_24603_, _24602_, _24600_);
  nor (_24604_, _09016_, _08809_);
  or (_24605_, _24604_, _24603_);
  and (_24606_, _24605_, _21260_);
  nor (_24607_, _24457_, _08806_);
  or (_24608_, _24411_, _07288_);
  or (_24610_, _09015_, \oc8051_golden_model_1.PSW [7]);
  and (_24611_, _24610_, _08808_);
  and (_24612_, _24611_, _24608_);
  or (_24613_, _24612_, _24607_);
  or (_24614_, _24613_, _24606_);
  and (_24615_, _24614_, _07965_);
  or (_24616_, _24615_, _24395_);
  and (_24617_, _24616_, _07996_);
  and (_24618_, _24419_, _07995_);
  or (_24619_, _24618_, _03155_);
  or (_24621_, _24619_, _24617_);
  nand (_24622_, _04790_, _03155_);
  and (_24623_, _24622_, _24621_);
  or (_24624_, _24623_, _02528_);
  or (_24625_, _09015_, _05790_);
  and (_24626_, _24625_, _03223_);
  and (_24627_, _24626_, _24624_);
  or (_24628_, _09692_, _08826_);
  nand (_24629_, _24404_, _09692_);
  and (_24630_, _24629_, _03040_);
  and (_24632_, _24630_, _24628_);
  or (_24633_, _24632_, _23374_);
  or (_24634_, _24633_, _24627_);
  and (_24635_, _24419_, _08789_);
  or (_24636_, _24635_, _21294_);
  and (_24637_, _24636_, _24634_);
  and (_24638_, _09015_, _08112_);
  or (_24639_, _24638_, _08115_);
  or (_24640_, _24639_, _24637_);
  or (_24641_, _24419_, _08116_);
  and (_24643_, _24641_, _24640_);
  or (_24644_, _24643_, _02890_);
  nand (_24645_, _04790_, _02890_);
  and (_24646_, _24645_, _08788_);
  and (_24647_, _24646_, _24644_);
  and (_24648_, _09015_, _02510_);
  or (_24649_, _24648_, _02889_);
  or (_24650_, _24649_, _24647_);
  and (_24651_, _09692_, _08828_);
  nor (_24652_, _24403_, _09692_);
  nor (_24654_, _24652_, _24651_);
  or (_24655_, _24654_, _03175_);
  and (_24656_, _24655_, _24650_);
  nor (_24657_, _24656_, _09725_);
  nor (_24658_, _24419_, _09724_);
  nor (_24659_, _24658_, _24657_);
  nor (_24660_, _24659_, _03174_);
  nor (_24661_, _09015_, _03179_);
  nor (_24662_, _24661_, _09733_);
  not (_24663_, _24662_);
  nor (_24665_, _24663_, _24660_);
  and (_24666_, _24419_, _09733_);
  nor (_24667_, _24666_, _03034_);
  not (_24668_, _24667_);
  nor (_24669_, _24668_, _24665_);
  and (_24670_, _03034_, _02924_);
  or (_24671_, _24670_, _02505_);
  nor (_24672_, _24671_, _24669_);
  and (_24673_, _09015_, _02505_);
  or (_24674_, _24673_, _02799_);
  nor (_24676_, _24674_, _24672_);
  nor (_24677_, _24654_, _03183_);
  nor (_24678_, _24677_, _09748_);
  not (_24679_, _24678_);
  nor (_24680_, _24679_, _24676_);
  nor (_24681_, _24457_, _09747_);
  nor (_24682_, _24681_, _02887_);
  not (_24683_, _24682_);
  nor (_24684_, _24683_, _24680_);
  nor (_24685_, _24684_, _24394_);
  nor (_24687_, _24685_, _09756_);
  nor (_24688_, _24419_, _09755_);
  nor (_24689_, _24688_, _03036_);
  not (_24690_, _24689_);
  nor (_24691_, _24690_, _24687_);
  nor (_24692_, _03038_, _02924_);
  nor (_24693_, _24692_, _24691_);
  or (_24694_, _24693_, _02499_);
  and (_24695_, _24694_, _24393_);
  nor (_24696_, _24695_, _08786_);
  and (_24698_, _24419_, _08786_);
  nor (_24699_, _24698_, _24696_);
  nand (_24700_, _24699_, _34655_);
  or (_24701_, _34655_, \oc8051_golden_model_1.PC [14]);
  and (_24702_, _24701_, _35796_);
  and (_35842_[14], _24702_, _24700_);
  nor (_24703_, _06905_, _06904_);
  nor (_24704_, _24703_, _06807_);
  and (_24705_, _24703_, _06807_);
  nor (_24706_, _24705_, _24704_);
  nor (_24708_, _06825_, _06824_);
  nor (_24709_, _24708_, _13763_);
  and (_24710_, _24708_, _13763_);
  nor (_24711_, _24710_, _24709_);
  and (_24712_, _24711_, _24706_);
  nor (_24713_, _24711_, _24706_);
  nor (_24714_, _24713_, _24712_);
  or (_24715_, _24714_, _05364_);
  nand (_24716_, _24714_, _05364_);
  and (_24717_, _24716_, _24715_);
  or (_24719_, _24717_, _03936_);
  and (_24720_, _07439_, _02509_);
  nor (_24721_, _24720_, _02510_);
  or (_24722_, _24721_, _24717_);
  and (_24723_, _03024_, _02532_);
  and (_24724_, _13516_, _13264_);
  nor (_24725_, _13516_, _13264_);
  nor (_24726_, _24725_, _24724_);
  not (_24727_, _24726_);
  not (_24728_, _14121_);
  and (_24730_, _24728_, _13804_);
  nor (_24731_, _24728_, _13804_);
  nor (_24732_, _24731_, _24730_);
  and (_24733_, _24732_, _24727_);
  nor (_24734_, _24732_, _24727_);
  nor (_24735_, _24734_, _24733_);
  not (_24736_, _15023_);
  nor (_24737_, _14724_, _14412_);
  and (_24738_, _14724_, _14412_);
  nor (_24739_, _24738_, _24737_);
  nor (_24741_, _24739_, _24736_);
  and (_24742_, _24739_, _24736_);
  nor (_24743_, _24742_, _24741_);
  nor (_24744_, _24743_, _24735_);
  and (_24745_, _24743_, _24735_);
  nor (_24746_, _24745_, _24744_);
  and (_24747_, _24746_, _07321_);
  nor (_24748_, _24746_, _07321_);
  or (_24749_, _24748_, _24747_);
  and (_24750_, _24749_, _05535_);
  or (_24752_, _24750_, _02841_);
  and (_24753_, _13573_, _13257_);
  nor (_24754_, _13573_, _13257_);
  or (_24755_, _24754_, _24753_);
  and (_24756_, _24755_, _13859_);
  nor (_24757_, _24755_, _13859_);
  or (_24758_, _24757_, _24756_);
  nand (_24759_, _24758_, _14179_);
  or (_24760_, _24758_, _14179_);
  and (_24761_, _24760_, _24759_);
  nor (_24763_, _14791_, _14473_);
  and (_24764_, _14791_, _14473_);
  nor (_24765_, _24764_, _24763_);
  not (_24766_, _15114_);
  and (_24767_, _24766_, _07493_);
  nor (_24768_, _24766_, _07493_);
  or (_24769_, _24768_, _24767_);
  or (_24770_, _24769_, _24765_);
  nand (_24771_, _24769_, _24765_);
  and (_24772_, _24771_, _24770_);
  nor (_24774_, _24772_, _24761_);
  and (_24775_, _24772_, _24761_);
  or (_24776_, _24775_, _24774_);
  and (_24777_, _24776_, _02877_);
  or (_24778_, _24717_, _02597_);
  or (_24779_, _24717_, _05361_);
  nor (_24780_, _24717_, _02601_);
  nor (_24781_, _24780_, _07433_);
  or (_24782_, _06168_, _06037_);
  nand (_24783_, _24782_, _10742_);
  or (_24785_, _24782_, _10742_);
  nand (_24786_, _24785_, _24783_);
  nor (_24787_, _06172_, _06129_);
  or (_24788_, _05855_, _05461_);
  or (_24789_, _06162_, _05810_);
  and (_24790_, _24789_, _24788_);
  nand (_24791_, _24790_, _24787_);
  or (_24792_, _24790_, _24787_);
  nand (_24793_, _24792_, _24791_);
  nand (_24794_, _24793_, _24786_);
  or (_24796_, _24793_, _24786_);
  and (_24797_, _24796_, _24794_);
  and (_24798_, _24797_, _07410_);
  nor (_24799_, _10559_, _05249_);
  and (_24800_, _10559_, _05249_);
  nor (_24801_, _24800_, _24799_);
  nor (_24802_, _05353_, _05251_);
  and (_24803_, _24802_, _04894_);
  nor (_24804_, _24802_, _04894_);
  or (_24805_, _24804_, _24803_);
  nand (_24807_, _24805_, _05260_);
  or (_24808_, _24805_, _05260_);
  and (_24809_, _24808_, _24807_);
  or (_24810_, _24809_, _24801_);
  nand (_24811_, _24809_, _24801_);
  and (_24812_, _24811_, _24810_);
  or (_24813_, _24812_, _07421_);
  or (_24814_, _24717_, _02602_);
  or (_24815_, _03382_, \oc8051_golden_model_1.PSW [0]);
  nand (_24816_, _24815_, _24814_);
  nand (_24818_, _24816_, _07421_);
  and (_24819_, _24818_, _07411_);
  and (_24820_, _24819_, _24813_);
  or (_24821_, _24820_, _02951_);
  or (_24822_, _24821_, _24798_);
  and (_24823_, _07638_, _07621_);
  nor (_24824_, _24823_, _07639_);
  and (_24825_, _24824_, _07566_);
  nor (_24826_, _24824_, _07566_);
  nor (_24827_, _24826_, _24825_);
  and (_24829_, _07596_, _07577_);
  and (_24830_, _07595_, _07578_);
  nor (_24831_, _24830_, _24829_);
  and (_24832_, _07607_, _07552_);
  nor (_24833_, _07607_, _07552_);
  or (_24834_, _24833_, _24832_);
  and (_24835_, _24834_, _24831_);
  nor (_24836_, _24834_, _24831_);
  or (_24837_, _24836_, _24835_);
  nor (_24838_, _24837_, _24827_);
  and (_24840_, _24837_, _24827_);
  nor (_24841_, _24840_, _24838_);
  nor (_24842_, _24841_, _05497_);
  and (_24843_, _24841_, _05497_);
  or (_24844_, _24843_, _24842_);
  or (_24845_, _24844_, _03401_);
  and (_24846_, _24845_, _19632_);
  and (_24847_, _24846_, _24822_);
  not (_24848_, xram_data_in_reg[5]);
  and (_24849_, xram_data_in_reg[1], xram_data_in_reg[0]);
  nor (_24851_, xram_data_in_reg[1], xram_data_in_reg[0]);
  nor (_24852_, _24851_, _24849_);
  nor (_24853_, _24852_, _24848_);
  and (_24854_, _24852_, _24848_);
  or (_24855_, _24854_, _24853_);
  and (_24856_, xram_data_in_reg[3], xram_data_in_reg[2]);
  nor (_24857_, xram_data_in_reg[3], xram_data_in_reg[2]);
  or (_24858_, _24857_, _24856_);
  and (_24859_, _24858_, xram_data_in_reg[4]);
  nor (_24860_, _24858_, xram_data_in_reg[4]);
  nor (_24862_, _24860_, _24859_);
  and (_24863_, xram_data_in_reg[6], xram_data_in_reg[7]);
  nor (_24864_, xram_data_in_reg[6], xram_data_in_reg[7]);
  or (_24865_, _24864_, _24863_);
  and (_24866_, _24865_, _24862_);
  nor (_24867_, _24865_, _24862_);
  or (_24868_, _24867_, _24866_);
  and (_24869_, _24868_, _24855_);
  nor (_24870_, _24868_, _24855_);
  or (_24871_, _24870_, _24869_);
  and (_24873_, _24871_, _07440_);
  or (_24874_, _24873_, _09169_);
  or (_24875_, _24874_, _24847_);
  and (_24876_, _24875_, _24781_);
  nand (_24877_, _24871_, _07433_);
  nand (_24878_, _24877_, _05361_);
  or (_24879_, _24878_, _24876_);
  and (_24880_, _24879_, _24779_);
  or (_24881_, _24880_, _03840_);
  nor (_24882_, _24708_, \oc8051_golden_model_1.ACC [6]);
  and (_24884_, _24708_, \oc8051_golden_model_1.ACC [6]);
  nor (_24885_, _24884_, _24882_);
  nor (_24886_, _24885_, _05364_);
  and (_24887_, _24885_, _05364_);
  nor (_24888_, _24887_, _24886_);
  and (_24889_, _24888_, _24786_);
  nor (_24890_, _24888_, _24786_);
  or (_24891_, _24890_, _05371_);
  or (_24892_, _24891_, _24889_);
  and (_24893_, _24892_, _24881_);
  or (_24895_, _24893_, _02948_);
  not (_24896_, _13294_);
  nor (_24897_, _13542_, _24896_);
  and (_24898_, _13542_, _24896_);
  nor (_24899_, _24898_, _24897_);
  and (_24900_, _24899_, _13827_);
  nor (_24901_, _24899_, _13827_);
  nor (_24902_, _24901_, _24900_);
  and (_24903_, _24902_, _14746_);
  nor (_24904_, _24902_, _14746_);
  or (_24906_, _24904_, _24903_);
  not (_24907_, _14426_);
  and (_24908_, _24907_, _14149_);
  nor (_24909_, _24907_, _14149_);
  nor (_24910_, _24909_, _24908_);
  and (_24911_, _24910_, _24906_);
  nor (_24912_, _24910_, _24906_);
  nor (_24913_, _24912_, _24911_);
  and (_24914_, _24913_, _15069_);
  nor (_24915_, _24913_, _15069_);
  or (_24917_, _24915_, _24914_);
  and (_24918_, _24917_, _07407_);
  nor (_24919_, _24917_, _07407_);
  or (_24920_, _24919_, _24918_);
  nor (_24921_, _24920_, _03006_);
  nor (_24922_, _24921_, _07405_);
  and (_24923_, _24922_, _24895_);
  and (_24924_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_24925_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_24926_, _24925_, _24924_);
  and (_24928_, _24926_, _13547_);
  nor (_24929_, _24926_, _13547_);
  nor (_24930_, _24929_, _24928_);
  and (_24931_, _14448_, _14156_);
  and (_24932_, _14447_, _14157_);
  nor (_24933_, _24932_, _24931_);
  nor (_24934_, _24933_, _24930_);
  and (_24935_, _24933_, _24930_);
  or (_24936_, _24935_, _24934_);
  nor (_24937_, _24936_, _14768_);
  and (_24939_, _24936_, _14768_);
  or (_24940_, _24939_, _24937_);
  not (_24941_, _24940_);
  nor (_24942_, _15092_, _07466_);
  and (_24943_, _15092_, _07466_);
  nor (_24944_, _24943_, _24942_);
  nand (_24945_, _24944_, _24941_);
  or (_24946_, _24944_, _24941_);
  and (_24947_, _24946_, _07405_);
  and (_24948_, _24947_, _24945_);
  or (_24950_, _24948_, _08996_);
  or (_24951_, _24950_, _24923_);
  not (_24952_, _08996_);
  or (_24953_, _24717_, _24952_);
  and (_24954_, _24953_, _02934_);
  and (_24955_, _24954_, _24951_);
  not (_24956_, _07472_);
  and (_24957_, _13555_, _13270_);
  nor (_24958_, _13555_, _13270_);
  or (_24959_, _24958_, _24957_);
  not (_24961_, _14161_);
  and (_24962_, _24961_, _13841_);
  nor (_24963_, _24961_, _13841_);
  nor (_24964_, _24963_, _24962_);
  and (_24965_, _24964_, _24959_);
  nor (_24966_, _24964_, _24959_);
  or (_24967_, _24966_, _24965_);
  nor (_24968_, _14772_, _14454_);
  and (_24969_, _14772_, _14454_);
  nor (_24970_, _24969_, _24968_);
  and (_24972_, _24970_, _15096_);
  nor (_24973_, _24970_, _15096_);
  nor (_24974_, _24973_, _24972_);
  nor (_24975_, _24974_, _24967_);
  and (_24976_, _24974_, _24967_);
  nor (_24977_, _24976_, _24975_);
  nand (_24978_, _24977_, _24956_);
  or (_24979_, _24977_, _24956_);
  and (_24980_, _24979_, _02884_);
  and (_24981_, _24980_, _24978_);
  or (_24983_, _24981_, _04225_);
  or (_24984_, _24983_, _24955_);
  and (_24985_, _24984_, _24778_);
  or (_24986_, _24985_, _02946_);
  or (_24987_, _24749_, _07474_);
  and (_24988_, _24987_, _07402_);
  and (_24989_, _24988_, _24986_);
  or (_24990_, _24812_, _03873_);
  and (_24991_, _24990_, _09187_);
  or (_24992_, _24991_, _24989_);
  or (_24993_, _24797_, _07481_);
  and (_24994_, _24993_, _02992_);
  and (_24995_, _24994_, _24992_);
  or (_24996_, _24844_, _09193_);
  and (_24997_, _24996_, _09194_);
  or (_24998_, _24997_, _24995_);
  or (_24999_, _24717_, _09200_);
  and (_25000_, _24999_, _02987_);
  and (_25001_, _25000_, _24998_);
  or (_25002_, _25001_, _24777_);
  and (_25005_, _09209_, _08986_);
  and (_25006_, _25005_, _22484_);
  and (_25007_, _25006_, _25002_);
  not (_25008_, _25006_);
  and (_25009_, _25008_, _24717_);
  or (_25010_, _25009_, _09252_);
  or (_25011_, _25010_, _25007_);
  or (_25012_, _24717_, _09251_);
  and (_25013_, _25012_, _06246_);
  and (_25014_, _25013_, _25011_);
  not (_25016_, _13864_);
  and (_25017_, _25016_, _13578_);
  nor (_25018_, _25016_, _13578_);
  nor (_25019_, _25018_, _25017_);
  and (_25020_, _25019_, _14743_);
  nor (_25021_, _25019_, _14743_);
  or (_25022_, _25021_, _25020_);
  nor (_25023_, _14126_, _24896_);
  and (_25024_, _14126_, _24896_);
  nor (_25025_, _25024_, _25023_);
  and (_25027_, _25025_, _14478_);
  nor (_25028_, _25025_, _14478_);
  nor (_25029_, _25028_, _25027_);
  nor (_25030_, _25029_, _25022_);
  and (_25031_, _25029_, _25022_);
  nor (_25032_, _25031_, _25030_);
  not (_25033_, _15065_);
  and (_25034_, _25033_, _07498_);
  nor (_25035_, _25033_, _07498_);
  nor (_25036_, _25035_, _25034_);
  or (_25037_, _25036_, _25032_);
  nand (_25038_, _25036_, _25032_);
  and (_25039_, _25038_, _02871_);
  and (_25040_, _25039_, _25037_);
  not (_25041_, _22918_);
  or (_25042_, _25041_, _09307_);
  or (_25043_, _25042_, _25040_);
  or (_25044_, _25043_, _25014_);
  not (_25045_, _25042_);
  or (_25046_, _25045_, _24717_);
  and (_25049_, _25046_, _06258_);
  and (_25050_, _25049_, _25044_);
  nor (_25051_, _13584_, _13319_);
  and (_25052_, _13584_, _13319_);
  or (_25053_, _25052_, _25051_);
  nor (_25054_, _25053_, _13869_);
  and (_25055_, _25053_, _13869_);
  nor (_25056_, _25055_, _25054_);
  nor (_25057_, _25056_, _14186_);
  and (_25058_, _25056_, _14186_);
  or (_25060_, _25058_, _25057_);
  nor (_25061_, _25060_, _14483_);
  and (_25062_, _25060_, _14483_);
  or (_25063_, _25062_, _25061_);
  nor (_25064_, _25063_, _14798_);
  and (_25065_, _25063_, _14798_);
  or (_25066_, _25065_, _25064_);
  nor (_25067_, _25066_, _15121_);
  and (_25068_, _25066_, _15121_);
  or (_25069_, _25068_, _25067_);
  or (_25070_, _25069_, _07503_);
  nand (_25071_, _25069_, _07503_);
  and (_25072_, _25071_, _06252_);
  nand (_25073_, _25072_, _25070_);
  and (_25074_, _07439_, _02939_);
  nor (_25075_, _25074_, _19627_);
  nand (_25076_, _25075_, _25073_);
  or (_25077_, _25076_, _25050_);
  or (_25078_, _25075_, _24717_);
  and (_25079_, _25078_, _10030_);
  and (_25082_, _25079_, _25077_);
  and (_25083_, _24717_, _02940_);
  or (_25084_, _25083_, _07400_);
  or (_25085_, _25084_, _25082_);
  not (_25086_, _07521_);
  and (_25087_, _13592_, _25086_);
  or (_25088_, _25087_, _07522_);
  nor (_25089_, _25088_, _13887_);
  and (_25090_, _25088_, _13887_);
  nor (_25091_, _25090_, _25089_);
  nand (_25093_, _25091_, _14201_);
  or (_25094_, _25091_, _14201_);
  and (_25095_, _25094_, _25093_);
  or (_25096_, _25095_, _14500_);
  nand (_25097_, _25095_, _14500_);
  and (_25098_, _25097_, _25096_);
  nor (_25099_, _25098_, _14814_);
  and (_25100_, _25098_, _14814_);
  or (_25101_, _25100_, _25099_);
  nor (_25102_, _25101_, _15060_);
  and (_25104_, _25101_, _15060_);
  nor (_25105_, _25104_, _25102_);
  or (_25106_, _25105_, _07535_);
  and (_25107_, _07534_, _07400_);
  nand (_25108_, _25107_, _25105_);
  nand (_25109_, _25108_, _25106_);
  and (_25110_, _07397_, _04138_);
  nor (_25111_, _25110_, _25109_);
  and (_25112_, _25111_, _25085_);
  nor (_25113_, _13600_, _07386_);
  and (_25115_, _13600_, _07386_);
  nor (_25116_, _25115_, _25113_);
  or (_25117_, _25116_, _14216_);
  nand (_25118_, _25116_, _14216_);
  and (_25119_, _25118_, _25117_);
  or (_25120_, _25119_, _13905_);
  nand (_25121_, _25119_, _13905_);
  and (_25122_, _25121_, _25120_);
  or (_25123_, _25122_, _14517_);
  nand (_25124_, _25122_, _14517_);
  and (_25125_, _25124_, _25123_);
  nor (_25126_, _25125_, _14830_);
  and (_25127_, _25125_, _14830_);
  or (_25128_, _25127_, _25126_);
  nor (_25129_, _25128_, _15047_);
  and (_25130_, _25128_, _15047_);
  or (_25131_, _25130_, _25129_);
  nor (_25132_, _25131_, _07396_);
  and (_25133_, _25131_, _07396_);
  or (_25134_, _25133_, _25132_);
  and (_25137_, _25134_, _25110_);
  or (_25138_, _25137_, _03451_);
  or (_25139_, _25138_, _25112_);
  not (_25140_, _03451_);
  or (_25141_, _25134_, _25140_);
  and (_25142_, _25141_, _02991_);
  and (_25143_, _25142_, _25139_);
  or (_25144_, _07707_, _07697_);
  and (_25145_, _25144_, _07708_);
  and (_25146_, _25145_, _13918_);
  nor (_25148_, _25145_, _13918_);
  or (_25149_, _25148_, _25146_);
  nor (_25150_, _25149_, _14228_);
  and (_25151_, _25149_, _14228_);
  or (_25152_, _25151_, _25150_);
  and (_25153_, _25152_, _14422_);
  nor (_25154_, _25152_, _14422_);
  or (_25155_, _25154_, _25153_);
  and (_25156_, _25155_, _14841_);
  nor (_25157_, _25155_, _14841_);
  or (_25159_, _25157_, _25156_);
  and (_25160_, _25159_, _15033_);
  nor (_25161_, _25159_, _15033_);
  or (_25162_, _25161_, _25160_);
  nor (_25163_, _25162_, _07717_);
  and (_25164_, _25162_, _07717_);
  or (_25165_, _25164_, _25163_);
  and (_25166_, _25165_, _02979_);
  or (_25167_, _25166_, _07540_);
  or (_25168_, _25167_, _25143_);
  or (_25170_, _07789_, _07780_);
  and (_25171_, _25170_, _07790_);
  nand (_25172_, _25171_, _13934_);
  or (_25173_, _25171_, _13934_);
  and (_25174_, _25173_, _25172_);
  nor (_25175_, _25174_, _14242_);
  and (_25176_, _25174_, _14242_);
  or (_25177_, _25176_, _25175_);
  and (_25178_, _14738_, _14533_);
  nor (_25179_, _14738_, _14533_);
  or (_25181_, _25179_, _25178_);
  and (_25182_, _25181_, _25177_);
  nor (_25183_, _25181_, _25177_);
  nor (_25184_, _25183_, _25182_);
  and (_25185_, _25184_, _15138_);
  nor (_25186_, _25184_, _15138_);
  nor (_25187_, _25186_, _25185_);
  nor (_25188_, _25187_, _07799_);
  and (_25189_, _25187_, _07799_);
  or (_25190_, _25189_, _25188_);
  or (_25192_, _25190_, _07541_);
  and (_25193_, _25192_, _25168_);
  or (_25194_, _25193_, _07721_);
  nor (_25195_, _04632_, _02925_);
  nor (_25196_, _04664_, _04658_);
  nor (_25197_, _04683_, _04652_);
  nor (_25198_, _04677_, _04645_);
  nor (_25199_, _25198_, _25197_);
  and (_25200_, _25198_, _25197_);
  nor (_25201_, _25200_, _25199_);
  nor (_25203_, _25201_, _25196_);
  and (_25204_, _25201_, _25196_);
  nor (_25205_, _25204_, _25203_);
  not (_25206_, _25205_);
  nor (_25207_, _25206_, _25195_);
  and (_25208_, _25206_, _25195_);
  or (_25209_, _25208_, _25207_);
  or (_25210_, _25209_, _02571_);
  and (_25211_, _25210_, _02986_);
  and (_25212_, _25211_, _25194_);
  not (_25214_, _07808_);
  nor (_25215_, _13614_, _13338_);
  and (_25216_, _13614_, _13338_);
  nor (_25217_, _25216_, _25215_);
  not (_25218_, _25217_);
  nor (_25219_, _14851_, _14541_);
  and (_25220_, _14851_, _14541_);
  nor (_25221_, _25220_, _25219_);
  and (_25222_, _25221_, _25218_);
  nor (_25223_, _25221_, _25218_);
  nor (_25225_, _25223_, _25222_);
  not (_25226_, _15146_);
  not (_25227_, _14250_);
  and (_25228_, _25227_, _13942_);
  nor (_25229_, _25227_, _13942_);
  nor (_25230_, _25229_, _25228_);
  nor (_25231_, _25230_, _25226_);
  and (_25232_, _25230_, _25226_);
  nor (_25233_, _25232_, _25231_);
  and (_25234_, _25233_, _25225_);
  nor (_25236_, _25233_, _25225_);
  nor (_25237_, _25236_, _25234_);
  nand (_25238_, _25237_, _25214_);
  or (_25239_, _25237_, _25214_);
  and (_25240_, _25239_, _02866_);
  and (_25241_, _25240_, _25238_);
  or (_25242_, _25241_, _22600_);
  or (_25243_, _25242_, _25212_);
  or (_25244_, _24717_, _22599_);
  and (_25245_, _25244_, _02859_);
  and (_25247_, _25245_, _25243_);
  or (_25248_, _25247_, _24752_);
  and (_25249_, _13621_, _13345_);
  nor (_25250_, _13621_, _13345_);
  nor (_25251_, _25250_, _25249_);
  not (_25252_, _14257_);
  and (_25253_, _25252_, _13949_);
  nor (_25254_, _25252_, _13949_);
  nor (_25255_, _25254_, _25253_);
  nor (_25256_, _25255_, _25251_);
  and (_25257_, _25255_, _25251_);
  or (_25258_, _25257_, _25256_);
  not (_25259_, _14858_);
  and (_25260_, _25259_, _14548_);
  nor (_25261_, _25259_, _14548_);
  nor (_25262_, _25261_, _25260_);
  nand (_25263_, _25262_, _15153_);
  or (_25264_, _25262_, _15153_);
  and (_25265_, _25264_, _25263_);
  nor (_25266_, _25265_, _25258_);
  and (_25269_, _25265_, _25258_);
  or (_25270_, _25269_, _25266_);
  nor (_25271_, _25270_, _07815_);
  and (_25272_, _25270_, _07815_);
  or (_25273_, _25272_, _02842_);
  or (_25274_, _25273_, _25271_);
  and (_25275_, _25274_, _02839_);
  and (_25276_, _25275_, _25248_);
  not (_25277_, _14553_);
  and (_25278_, _13626_, _13350_);
  nor (_25280_, _13626_, _13350_);
  nor (_25281_, _25280_, _25278_);
  not (_25282_, _25281_);
  not (_25283_, _14262_);
  and (_25284_, _25283_, _13954_);
  nor (_25285_, _25283_, _13954_);
  nor (_25286_, _25285_, _25284_);
  and (_25287_, _25286_, _25282_);
  nor (_25288_, _25286_, _25282_);
  or (_25289_, _25288_, _25287_);
  nor (_25291_, _25289_, _25277_);
  and (_25292_, _25289_, _25277_);
  or (_25293_, _25292_, _25291_);
  and (_25294_, _25293_, _14863_);
  nor (_25295_, _25293_, _14863_);
  or (_25296_, _25295_, _25294_);
  and (_25297_, _25296_, _15158_);
  nor (_25298_, _25296_, _15158_);
  or (_25299_, _25298_, _25297_);
  and (_25300_, _25299_, _07820_);
  nor (_25302_, _25299_, _07820_);
  or (_25303_, _25302_, _25300_);
  and (_25304_, _25303_, _02567_);
  or (_25305_, _25304_, _06786_);
  or (_25306_, _25305_, _25276_);
  and (_25307_, _06840_, _15163_);
  nor (_25308_, _06840_, _15163_);
  nor (_25309_, _25308_, _25307_);
  not (_25310_, _25309_);
  not (_25311_, _06872_);
  nor (_25313_, _06925_, _25311_);
  and (_25314_, _06925_, _25311_);
  nor (_25315_, _25314_, _25313_);
  not (_25316_, _25315_);
  and (_25317_, _25316_, _06978_);
  nor (_25318_, _25316_, _06978_);
  nor (_25319_, _25318_, _25317_);
  and (_25320_, _25319_, _25310_);
  nor (_25321_, _25319_, _25310_);
  nor (_25322_, _25321_, _25320_);
  and (_25324_, _07050_, _06805_);
  nor (_25325_, _07050_, _06805_);
  nor (_25326_, _25325_, _25324_);
  and (_25327_, _25326_, _25322_);
  nor (_25328_, _25326_, _25322_);
  nor (_25329_, _25328_, _25327_);
  and (_25330_, _25329_, _07133_);
  nor (_25331_, _25329_, _07133_);
  or (_25332_, _25331_, _06792_);
  or (_25333_, _25332_, _25330_);
  and (_25335_, _25333_, _02609_);
  and (_25336_, _25335_, _25306_);
  nand (_25337_, _25209_, _02542_);
  not (_25338_, _04075_);
  and (_25339_, _02968_, _02521_);
  nor (_25340_, _25339_, _03510_);
  and (_25341_, _25340_, _25338_);
  and (_25342_, _04393_, _03297_);
  nor (_25343_, _25342_, _05743_);
  and (_25344_, _25343_, _25341_);
  and (_25346_, _09366_, _09360_);
  and (_25347_, _25346_, _04080_);
  and (_25348_, _25347_, _25344_);
  nand (_25349_, _25348_, _25337_);
  or (_25350_, _25349_, _25336_);
  or (_25351_, _25348_, _24717_);
  and (_25352_, _25351_, _07140_);
  and (_25353_, _25352_, _25350_);
  nor (_25354_, _14273_, _13965_);
  and (_25355_, _14273_, _13965_);
  nor (_25357_, _25355_, _25354_);
  nor (_25358_, _13637_, _13361_);
  and (_25359_, _13637_, _13361_);
  or (_25360_, _25359_, _25358_);
  nor (_25361_, _25360_, _25357_);
  and (_25362_, _25360_, _25357_);
  nor (_25363_, _25362_, _25361_);
  not (_25364_, _15171_);
  nor (_25365_, _14874_, _14564_);
  and (_25366_, _14874_, _14564_);
  nor (_25368_, _25366_, _25365_);
  nor (_25369_, _25368_, _25364_);
  and (_25370_, _25368_, _25364_);
  nor (_25371_, _25370_, _25369_);
  nor (_25372_, _25371_, _25363_);
  and (_25373_, _25371_, _25363_);
  or (_25374_, _25373_, _25372_);
  or (_25375_, _25374_, _07833_);
  nand (_25376_, _25374_, _07833_);
  and (_25377_, _25376_, _02834_);
  and (_25379_, _25377_, _25375_);
  or (_25380_, _25379_, _25353_);
  and (_25381_, _25380_, _07831_);
  nand (_25382_, _25209_, _07830_);
  and (_25383_, _09415_, _19622_);
  and (_25384_, _25383_, _19621_);
  nand (_25385_, _25384_, _25382_);
  or (_25386_, _25385_, _25381_);
  or (_25387_, _25384_, _24717_);
  and (_25388_, _25387_, _07844_);
  and (_25390_, _25388_, _25386_);
  not (_25391_, _07844_);
  not (_25392_, _07195_);
  and (_25393_, _25392_, _07192_);
  nor (_25394_, _25392_, _07192_);
  nor (_25395_, _25394_, _25393_);
  and (_25396_, _13369_, _07211_);
  nor (_25397_, _25396_, _13880_);
  nor (_25398_, _14192_, _07207_);
  and (_25399_, _14192_, _07207_);
  nor (_25401_, _25399_, _25398_);
  nor (_25402_, _25401_, _25397_);
  and (_25403_, _25401_, _25397_);
  nor (_25404_, _25403_, _25402_);
  nor (_25405_, _07198_, _07202_);
  and (_25406_, _07198_, _07202_);
  nor (_25407_, _25406_, _25405_);
  nor (_25408_, _25407_, _25404_);
  and (_25409_, _25407_, _25404_);
  nor (_25410_, _25409_, _25408_);
  nor (_25412_, _25410_, _25395_);
  and (_25413_, _25410_, _25395_);
  or (_25414_, _25413_, _25412_);
  and (_25415_, _25414_, _25391_);
  or (_25416_, _25415_, _25390_);
  and (_25417_, _25416_, _07838_);
  not (_25418_, _07838_);
  and (_25419_, _25414_, _25418_);
  or (_25420_, _25419_, _07849_);
  or (_25421_, _25420_, _25417_);
  nor (_25423_, _14207_, _08046_);
  and (_25424_, _14207_, _08046_);
  nor (_25425_, _25424_, _25423_);
  and (_25426_, _13249_, _08050_);
  nor (_25427_, _25426_, _13898_);
  nor (_25428_, _25427_, _25425_);
  and (_25429_, _25427_, _25425_);
  nor (_25430_, _25429_, _25428_);
  nor (_25431_, _08041_, _08034_);
  and (_25432_, _08041_, _08034_);
  nor (_25433_, _25432_, _25431_);
  nor (_25434_, _25433_, _08037_);
  and (_25435_, _25433_, _08037_);
  nor (_25436_, _25435_, _25434_);
  nor (_25437_, _25436_, _25430_);
  and (_25438_, _25436_, _25430_);
  or (_25439_, _25438_, _25437_);
  and (_25440_, _25439_, _07856_);
  nor (_25441_, _25439_, _07856_);
  or (_25442_, _25441_, _25440_);
  or (_25445_, _25442_, _07850_);
  and (_25446_, _25445_, _03147_);
  and (_25447_, _25446_, _25421_);
  nor (_25448_, _10565_, _10369_);
  and (_25449_, _10565_, _10369_);
  nor (_25450_, _25449_, _25448_);
  nor (_25451_, _10964_, _10766_);
  and (_25452_, _10964_, _10766_);
  nor (_25453_, _25452_, _25451_);
  nor (_25454_, _25453_, _25450_);
  and (_25456_, _25453_, _25450_);
  nor (_25457_, _25456_, _25454_);
  nor (_25458_, _11356_, _11154_);
  and (_25459_, _11356_, _11154_);
  nor (_25460_, _25459_, _25458_);
  nor (_25461_, _11556_, _05772_);
  and (_25462_, _11556_, _05772_);
  nor (_25463_, _25462_, _25461_);
  not (_25464_, _25463_);
  and (_25465_, _25464_, _25460_);
  nor (_25467_, _25464_, _25460_);
  nor (_25468_, _25467_, _25465_);
  and (_25469_, _25468_, _25457_);
  nor (_25470_, _25468_, _25457_);
  or (_25471_, _25470_, _25469_);
  and (_25472_, _25471_, _03146_);
  or (_25473_, _25472_, _25447_);
  and (_25474_, _25473_, _07861_);
  and (_25475_, _09273_, _09272_);
  nor (_25476_, _25475_, _09274_);
  and (_25478_, _09269_, _08130_);
  nor (_25479_, _25478_, _09270_);
  and (_25480_, _25479_, _25476_);
  nor (_25481_, _25479_, _25476_);
  or (_25482_, _25481_, _25480_);
  not (_25483_, _08125_);
  and (_25484_, _25483_, _08120_);
  nor (_25485_, _25483_, _08120_);
  nor (_25486_, _25485_, _25484_);
  and (_25487_, _25486_, _09265_);
  nor (_25489_, _25486_, _09265_);
  nor (_25490_, _25489_, _25487_);
  nor (_25491_, _25490_, _25482_);
  and (_25492_, _25490_, _25482_);
  nor (_25493_, _25492_, _25491_);
  nand (_25494_, _25493_, _07867_);
  or (_25495_, _25493_, _07867_);
  and (_25496_, _25495_, _25494_);
  and (_25497_, _25496_, _07860_);
  or (_25498_, _25497_, _03051_);
  or (_25500_, _25498_, _25474_);
  not (_25501_, _14407_);
  nor (_25502_, _13513_, _13259_);
  and (_25503_, _13513_, _13259_);
  nor (_25504_, _25503_, _25502_);
  not (_25505_, _25504_);
  not (_25506_, _14117_);
  and (_25507_, _25506_, _13798_);
  nor (_25508_, _25506_, _13798_);
  nor (_25509_, _25508_, _25507_);
  and (_25511_, _25509_, _25505_);
  nor (_25512_, _25509_, _25505_);
  or (_25513_, _25512_, _25511_);
  nor (_25514_, _25513_, _25501_);
  and (_25515_, _25513_, _25501_);
  or (_25516_, _25515_, _25514_);
  and (_25517_, _25516_, _14719_);
  nor (_25518_, _25516_, _14719_);
  or (_25519_, _25518_, _25517_);
  and (_25520_, _25519_, _15019_);
  nor (_25522_, _25519_, _15019_);
  or (_25523_, _25522_, _25520_);
  and (_25524_, _25523_, _07317_);
  nor (_25525_, _25523_, _07317_);
  or (_25526_, _25525_, _25524_);
  or (_25527_, _25526_, _07139_);
  and (_25528_, _25527_, _07150_);
  and (_25529_, _25528_, _25500_);
  nand (_25530_, _24717_, _03148_);
  or (_25531_, _25530_, _04731_);
  nand (_25533_, _25531_, _23315_);
  or (_25534_, _25533_, _25529_);
  and (_25535_, _03298_, _02529_);
  nor (_25536_, _24717_, _23315_);
  nor (_25537_, _25536_, _25535_);
  and (_25538_, _25537_, _25534_);
  or (_25539_, _07212_, _07209_);
  nand (_25540_, _07212_, _07209_);
  and (_25541_, _25540_, _25539_);
  nand (_25542_, _25541_, _14001_);
  or (_25544_, _25541_, _14001_);
  and (_25545_, _25544_, _25542_);
  nor (_25546_, _25545_, _07203_);
  and (_25547_, _25545_, _07203_);
  or (_25548_, _25547_, _25546_);
  not (_25549_, _07196_);
  nor (_25550_, _07200_, _07193_);
  and (_25551_, _07200_, _07193_);
  nor (_25552_, _25551_, _25550_);
  nor (_25553_, _25552_, _25549_);
  and (_25555_, _25552_, _25549_);
  nor (_25556_, _25555_, _25553_);
  not (_25557_, _25556_);
  nor (_25558_, _25557_, _25548_);
  and (_25559_, _25557_, _25548_);
  nor (_25560_, _25559_, _25558_);
  nand (_25561_, _25560_, _07191_);
  or (_25562_, _25560_, _07191_);
  and (_25563_, _25562_, _25561_);
  and (_25564_, _25563_, _25535_);
  or (_25566_, _25564_, _03534_);
  or (_25567_, _25566_, _25538_);
  not (_25568_, _03534_);
  or (_25569_, _25563_, _25568_);
  and (_25570_, _25569_, _07881_);
  and (_25571_, _25570_, _25567_);
  and (_25572_, _25563_, _07880_);
  or (_25573_, _25572_, _07890_);
  or (_25574_, _25573_, _25571_);
  or (_25575_, _08051_, _08048_);
  nand (_25577_, _08051_, _08048_);
  and (_25578_, _25577_, _25575_);
  not (_25579_, _08042_);
  and (_25580_, _25579_, _08044_);
  nor (_25581_, _25579_, _08044_);
  nor (_25582_, _25581_, _25580_);
  not (_25583_, _25582_);
  and (_25584_, _25583_, _25578_);
  nor (_25585_, _25583_, _25578_);
  nor (_25586_, _25585_, _25584_);
  nor (_25588_, _08035_, _08039_);
  and (_25589_, _08035_, _08039_);
  nor (_25590_, _25589_, _25588_);
  and (_25591_, _08032_, _07855_);
  nor (_25592_, _25591_, _10161_);
  nor (_25593_, _25592_, _25590_);
  and (_25594_, _25592_, _25590_);
  nor (_25595_, _25594_, _25593_);
  or (_25596_, _25595_, _25586_);
  nand (_25597_, _25595_, _25586_);
  and (_25599_, _25597_, _25596_);
  or (_25600_, _25599_, _07891_);
  and (_25601_, _25600_, _03136_);
  and (_25602_, _25601_, _25574_);
  nor (_25603_, _10563_, _10368_);
  and (_25604_, _10563_, _10368_);
  nor (_25605_, _25604_, _25603_);
  not (_25606_, _25605_);
  not (_25607_, _10963_);
  and (_25608_, _25607_, _10764_);
  nor (_25610_, _25607_, _10764_);
  nor (_25611_, _25610_, _25608_);
  nor (_25612_, _25611_, _25606_);
  and (_25613_, _25611_, _25606_);
  nor (_25614_, _25613_, _25612_);
  not (_25615_, _11554_);
  nor (_25616_, _11354_, _11153_);
  and (_25617_, _11354_, _11153_);
  nor (_25618_, _25617_, _25616_);
  nor (_25619_, _25618_, _25615_);
  and (_25621_, _25618_, _25615_);
  nor (_25622_, _25621_, _25619_);
  not (_25623_, _25622_);
  nor (_25624_, _25623_, _25614_);
  and (_25625_, _25623_, _25614_);
  or (_25626_, _25625_, _25624_);
  not (_25627_, _25626_);
  nand (_25628_, _25627_, _05770_);
  or (_25629_, _25627_, _05770_);
  and (_25630_, _25629_, _03135_);
  and (_25631_, _25630_, _25628_);
  or (_25632_, _25631_, _07311_);
  or (_25633_, _25632_, _25602_);
  or (_25634_, _07781_, _08132_);
  nand (_25635_, _07781_, _08132_);
  and (_25636_, _25635_, _25634_);
  not (_25637_, _08126_);
  and (_25638_, _25637_, _08128_);
  nor (_25639_, _25637_, _08128_);
  nor (_25640_, _25639_, _25638_);
  and (_25643_, _25640_, _25636_);
  nor (_25644_, _25640_, _25636_);
  nor (_25645_, _25644_, _25643_);
  or (_25646_, _25645_, _08123_);
  nand (_25647_, _25645_, _08123_);
  and (_25648_, _25647_, _25646_);
  or (_25649_, _25648_, _08121_);
  nand (_25650_, _25648_, _08121_);
  and (_25651_, _25650_, _25649_);
  or (_25652_, _25651_, _08118_);
  nand (_25654_, _25651_, _08118_);
  and (_25655_, _25654_, _25652_);
  and (_25656_, _25655_, _07865_);
  nor (_25657_, _25655_, _07865_);
  or (_25658_, _25657_, _25656_);
  or (_25659_, _25658_, _07312_);
  and (_25660_, _25659_, _03023_);
  and (_25661_, _25660_, _25633_);
  and (_25662_, _08819_, _09470_);
  nor (_25663_, _14017_, _13417_);
  and (_25665_, _14017_, _13417_);
  nor (_25666_, _25665_, _25663_);
  nor (_25667_, _15209_, _14608_);
  and (_25668_, _15209_, _14608_);
  nor (_25669_, _25668_, _25667_);
  and (_25670_, _25669_, _25666_);
  nor (_25671_, _25669_, _25666_);
  nor (_25672_, _25671_, _25670_);
  nor (_25673_, _14916_, _14307_);
  and (_25674_, _14916_, _14307_);
  nor (_25676_, _25674_, _25673_);
  nor (_25677_, _13690_, _07901_);
  and (_25678_, _13690_, _07901_);
  nor (_25679_, _25678_, _25677_);
  and (_25680_, _25679_, _25676_);
  nor (_25681_, _25679_, _25676_);
  nor (_25682_, _25681_, _25680_);
  not (_25683_, _25682_);
  nand (_25684_, _25683_, _25672_);
  or (_25685_, _25683_, _25672_);
  and (_25687_, _25685_, _03022_);
  nand (_25688_, _25687_, _25684_);
  nand (_25689_, _25688_, _25662_);
  or (_25690_, _25689_, _25661_);
  and (_25691_, _02959_, _02532_);
  nor (_25692_, _13416_, _25691_);
  or (_25693_, _24717_, _25662_);
  and (_25694_, _25693_, _07913_);
  and (_25695_, _25694_, _25692_);
  and (_25696_, _25695_, _25690_);
  and (_25698_, _07915_, _04138_);
  nor (_25699_, _13368_, _07210_);
  and (_25700_, _13368_, _07210_);
  nor (_25701_, _25700_, _25699_);
  not (_25702_, _25701_);
  not (_25703_, _07204_);
  and (_25704_, _25703_, _07206_);
  nor (_25705_, _25703_, _07206_);
  nor (_25706_, _25705_, _25704_);
  nor (_25707_, _25706_, _25702_);
  and (_25709_, _25706_, _25702_);
  nor (_25710_, _25709_, _25707_);
  nor (_25711_, _07201_, _07194_);
  and (_25712_, _07201_, _07194_);
  nor (_25713_, _25712_, _25711_);
  nor (_25714_, _25713_, _14923_);
  and (_25715_, _25713_, _14923_);
  nor (_25716_, _25715_, _25714_);
  not (_25717_, _25716_);
  nor (_25718_, _25717_, _25710_);
  and (_25720_, _25717_, _25710_);
  nor (_25721_, _25720_, _25718_);
  or (_25722_, _25721_, _07190_);
  nand (_25723_, _25721_, _07190_);
  and (_25724_, _25723_, _14312_);
  and (_25725_, _25724_, _25722_);
  or (_25726_, _25725_, _25698_);
  or (_25727_, _25726_, _25696_);
  nand (_25728_, _03014_, _02532_);
  nor (_25729_, _13248_, _08049_);
  and (_25731_, _13248_, _08049_);
  nor (_25732_, _25731_, _25729_);
  not (_25733_, _08043_);
  and (_25734_, _25733_, _08045_);
  nor (_25735_, _25733_, _08045_);
  nor (_25736_, _25735_, _25734_);
  and (_25737_, _25736_, _25732_);
  nor (_25738_, _25736_, _25732_);
  nor (_25739_, _25738_, _25737_);
  nor (_25740_, _08040_, _08033_);
  and (_25742_, _08040_, _08033_);
  nor (_25743_, _25742_, _25740_);
  and (_25744_, _25743_, _08036_);
  nor (_25745_, _25743_, _08036_);
  nor (_25746_, _25745_, _25744_);
  and (_25747_, _25746_, _25739_);
  nor (_25748_, _25746_, _25739_);
  or (_25749_, _25748_, _25747_);
  nand (_25750_, _25749_, _07854_);
  or (_25751_, _25749_, _07854_);
  and (_25753_, _25751_, _25750_);
  or (_25754_, _25753_, _25728_);
  and (_25755_, _25754_, _25727_);
  or (_25756_, _25755_, _24723_);
  not (_25757_, _24723_);
  or (_25758_, _25753_, _25757_);
  and (_25759_, _25758_, _03142_);
  and (_25760_, _25759_, _25756_);
  nor (_25761_, _10564_, _10367_);
  and (_25762_, _10564_, _10367_);
  nor (_25764_, _25762_, _25761_);
  and (_25765_, _25764_, _10765_);
  nor (_25766_, _25764_, _10765_);
  or (_25767_, _25766_, _25765_);
  nand (_25768_, _25767_, _10962_);
  or (_25769_, _25767_, _10962_);
  and (_25770_, _25769_, _25768_);
  nor (_25771_, _11355_, _11152_);
  and (_25772_, _11355_, _11152_);
  nor (_25773_, _25772_, _25771_);
  nor (_25775_, _25773_, _11555_);
  and (_25776_, _25773_, _11555_);
  nor (_25777_, _25776_, _25775_);
  and (_25778_, _25777_, _25770_);
  nor (_25779_, _25777_, _25770_);
  nor (_25780_, _25779_, _25778_);
  and (_25781_, _25780_, _05771_);
  nor (_25782_, _25780_, _05771_);
  or (_25783_, _25782_, _25781_);
  and (_25784_, _25783_, _03141_);
  or (_25786_, _25784_, _07921_);
  or (_25787_, _25786_, _25760_);
  nor (_25788_, _07782_, _09271_);
  and (_25789_, _07782_, _09271_);
  nor (_25790_, _25789_, _25788_);
  not (_25791_, _08127_);
  and (_25792_, _25791_, _08129_);
  nor (_25793_, _25791_, _08129_);
  nor (_25794_, _25793_, _25792_);
  and (_25795_, _25794_, _25790_);
  nor (_25797_, _25794_, _25790_);
  nor (_25798_, _25797_, _25795_);
  not (_25799_, _08124_);
  nor (_25800_, _08122_, _08119_);
  and (_25801_, _08122_, _08119_);
  nor (_25802_, _25801_, _25800_);
  nor (_25803_, _25802_, _25799_);
  and (_25804_, _25802_, _25799_);
  nor (_25805_, _25804_, _25803_);
  and (_25806_, _25805_, _25798_);
  nor (_25808_, _25805_, _25798_);
  or (_25809_, _25808_, _25806_);
  and (_25810_, _25809_, _07866_);
  nor (_25811_, _25809_, _07866_);
  or (_25812_, _25811_, _25810_);
  or (_25813_, _25812_, _13434_);
  and (_25814_, _25813_, _03043_);
  and (_25815_, _25814_, _25787_);
  and (_25816_, _08809_, _19607_);
  nor (_25817_, _13711_, _13442_);
  and (_25819_, _13711_, _13442_);
  or (_25820_, _25819_, _25817_);
  not (_25821_, _14324_);
  and (_25822_, _25821_, _14039_);
  nor (_25823_, _25821_, _14039_);
  nor (_25824_, _25823_, _25822_);
  nor (_25825_, _25824_, _25820_);
  and (_25826_, _25824_, _25820_);
  or (_25827_, _25826_, _25825_);
  not (_25828_, _14943_);
  and (_25830_, _25828_, _14630_);
  nor (_25831_, _25828_, _14630_);
  nor (_25832_, _25831_, _25830_);
  not (_25833_, _15231_);
  and (_25834_, _25833_, _07929_);
  nor (_25835_, _25833_, _07929_);
  nor (_25836_, _25835_, _25834_);
  or (_25837_, _25836_, _25832_);
  nand (_25838_, _25836_, _25832_);
  and (_25839_, _25838_, _25837_);
  nor (_25841_, _25839_, _25827_);
  and (_25842_, _25839_, _25827_);
  or (_25843_, _25842_, _03043_);
  or (_25844_, _25843_, _25841_);
  nand (_25845_, _25844_, _25816_);
  or (_25846_, _25845_, _25815_);
  nor (_25847_, _24717_, _25816_);
  nor (_25848_, _25847_, _07230_);
  and (_25849_, _25848_, _25846_);
  not (_25850_, _14713_);
  not (_25852_, _14112_);
  nor (_25853_, _07521_, _07287_);
  nor (_25854_, _13716_, _25086_);
  nor (_25855_, _25854_, _25853_);
  nor (_25856_, _25855_, _14044_);
  and (_25857_, _25855_, _14044_);
  nor (_25858_, _25857_, _25856_);
  and (_25859_, _25858_, _25852_);
  nor (_25860_, _25858_, _25852_);
  nor (_25861_, _25860_, _25859_);
  nor (_25863_, _25861_, _14635_);
  and (_25864_, _25861_, _14635_);
  or (_25865_, _25864_, _25863_);
  nor (_25866_, _25865_, _25850_);
  and (_25867_, _25865_, _25850_);
  nor (_25868_, _25867_, _25866_);
  nor (_25869_, _25868_, _15236_);
  and (_25870_, _25868_, _15236_);
  or (_25871_, _25870_, _25869_);
  nand (_25872_, _25871_, _07307_);
  or (_25874_, _25871_, _07307_);
  and (_25875_, _25874_, _25872_);
  and (_25876_, _25875_, _07230_);
  or (_25877_, _25876_, _07233_);
  or (_25878_, _25877_, _25849_);
  or (_25879_, _25875_, _07232_);
  and (_25880_, _25879_, _07936_);
  and (_25881_, _25880_, _25878_);
  nor (_25882_, _13721_, _07386_);
  and (_25883_, _13721_, _07386_);
  or (_25885_, _25883_, _25882_);
  nor (_25886_, _25885_, _14049_);
  and (_25887_, _25885_, _14049_);
  nor (_25888_, _25887_, _25886_);
  nor (_25889_, _25888_, _14331_);
  and (_25890_, _25888_, _14331_);
  or (_25891_, _25890_, _25889_);
  and (_25892_, _25891_, _14640_);
  nor (_25893_, _25891_, _14640_);
  or (_25894_, _25893_, _25892_);
  nor (_25896_, _25894_, _14950_);
  and (_25897_, _25894_, _14950_);
  or (_25898_, _25897_, _25896_);
  nor (_25899_, _25898_, _15241_);
  and (_25900_, _25898_, _15241_);
  or (_25901_, _25900_, _25899_);
  nand (_25902_, _25901_, _07960_);
  or (_25903_, _25901_, _07960_);
  and (_25904_, _25903_, _07229_);
  and (_25905_, _25904_, _25902_);
  or (_25907_, _25905_, _25881_);
  and (_25908_, _25907_, _03134_);
  nor (_25909_, _13726_, _07697_);
  and (_25910_, _13726_, _07697_);
  or (_25911_, _25910_, _25909_);
  nor (_25912_, _25911_, _13792_);
  and (_25913_, _25911_, _13792_);
  nor (_25914_, _25913_, _25912_);
  nor (_25915_, _25914_, _14336_);
  and (_25916_, _25914_, _14336_);
  or (_25918_, _25916_, _25915_);
  nor (_25919_, _25918_, _14645_);
  and (_25920_, _25918_, _14645_);
  or (_25921_, _25920_, _25919_);
  nor (_25922_, _25921_, _14955_);
  and (_25923_, _25921_, _14955_);
  or (_25924_, _25923_, _25922_);
  and (_25925_, _25924_, _15246_);
  nor (_25926_, _25924_, _15246_);
  or (_25927_, _25926_, _25925_);
  nand (_25929_, _25927_, _07991_);
  or (_25930_, _25927_, _07991_);
  and (_25931_, _25930_, _03133_);
  and (_25932_, _25931_, _25929_);
  or (_25933_, _25932_, _07964_);
  or (_25934_, _25933_, _25908_);
  and (_25935_, _13731_, _07780_);
  nor (_25936_, _13731_, _07780_);
  nor (_25937_, _25936_, _25935_);
  nor (_25938_, _25937_, _14055_);
  and (_25940_, _25937_, _14055_);
  nor (_25941_, _25940_, _25938_);
  or (_25942_, _25941_, _14341_);
  nand (_25943_, _25941_, _14341_);
  and (_25944_, _25943_, _25942_);
  nor (_25945_, _25944_, _14650_);
  and (_25946_, _25944_, _14650_);
  nor (_25947_, _25946_, _25945_);
  or (_25948_, _25947_, _14960_);
  nand (_25949_, _25947_, _14960_);
  and (_25951_, _25949_, _25948_);
  nor (_25952_, _25951_, _15252_);
  and (_25953_, _25951_, _15252_);
  nor (_25954_, _25953_, _25952_);
  nor (_25955_, _25954_, _08022_);
  and (_25956_, _25954_, _08022_);
  or (_25957_, _25956_, _25955_);
  or (_25958_, _25957_, _07997_);
  and (_25959_, _25958_, _07996_);
  and (_25960_, _25959_, _25934_);
  nor (_25962_, _03155_, _02528_);
  and (_25963_, _25962_, _03223_);
  and (_25964_, _25963_, _07996_);
  nor (_25965_, _07702_, _07701_);
  nor (_25966_, _13833_, \oc8051_golden_model_1.ACC [3]);
  and (_25967_, _13833_, \oc8051_golden_model_1.ACC [3]);
  nor (_25968_, _25967_, _25966_);
  and (_25969_, _25968_, _24885_);
  nor (_25970_, _25968_, _24885_);
  nor (_25971_, _25970_, _25969_);
  nor (_25973_, _25971_, _25965_);
  and (_25974_, _25971_, _25965_);
  nor (_25975_, _25974_, _25973_);
  and (_25976_, _25975_, _25963_);
  nor (_25977_, _25976_, _25964_);
  or (_25978_, _25977_, _25960_);
  or (_25979_, _25963_, _24717_);
  and (_25980_, _25979_, _25978_);
  or (_25981_, _25980_, _10153_);
  not (_25982_, _13368_);
  and (_25983_, _25982_, _07211_);
  nor (_25984_, _25982_, _07211_);
  nor (_25985_, _25984_, _25983_);
  and (_25986_, _25985_, _14062_);
  nor (_25987_, _25985_, _14062_);
  nor (_25988_, _25987_, _25986_);
  and (_25989_, _25988_, _14349_);
  nor (_25990_, _25988_, _14349_);
  nor (_25991_, _25990_, _25989_);
  and (_25992_, _25991_, _14657_);
  nor (_25995_, _25991_, _14657_);
  nor (_25996_, _25995_, _25992_);
  nor (_25997_, _25996_, _14710_);
  and (_25998_, _25996_, _14710_);
  or (_25999_, _25998_, _25997_);
  and (_26000_, _25999_, _15261_);
  nor (_26001_, _25999_, _15261_);
  or (_26002_, _26001_, _26000_);
  nor (_26003_, _26002_, _07227_);
  and (_26004_, _26002_, _07227_);
  or (_26006_, _26004_, _26003_);
  or (_26007_, _26006_, _07189_);
  and (_26008_, _26007_, _25981_);
  or (_26009_, _26008_, _07185_);
  not (_26010_, _13248_);
  and (_26011_, _26010_, _08050_);
  nor (_26012_, _26010_, _08050_);
  nor (_26013_, _26012_, _26011_);
  and (_26014_, _26013_, _14067_);
  nor (_26015_, _26013_, _14067_);
  nor (_26017_, _26015_, _26014_);
  and (_26018_, _26017_, _14355_);
  nor (_26019_, _26017_, _14355_);
  nor (_26020_, _26019_, _26018_);
  and (_26021_, _26020_, _14662_);
  nor (_26022_, _26020_, _14662_);
  nor (_26023_, _26022_, _26021_);
  nor (_26024_, _26023_, _14970_);
  and (_26025_, _26023_, _14970_);
  or (_26026_, _26025_, _26024_);
  nor (_26028_, _26026_, _15266_);
  and (_26029_, _26026_, _15266_);
  or (_26030_, _26029_, _26028_);
  and (_26031_, _26030_, _08066_);
  nor (_26032_, _26030_, _08066_);
  or (_26033_, _26032_, _26031_);
  or (_26034_, _26033_, _08031_);
  and (_26035_, _26034_, _08789_);
  and (_26036_, _26035_, _26009_);
  nor (_26037_, _13754_, _09272_);
  nor (_26039_, _26037_, _25475_);
  nor (_26040_, _26039_, _14073_);
  and (_26041_, _26039_, _14073_);
  or (_26042_, _26041_, _26040_);
  nor (_26043_, _26042_, _14367_);
  and (_26044_, _26042_, _14367_);
  nor (_26045_, _26044_, _26043_);
  nor (_26046_, _26045_, _14670_);
  and (_26047_, _26045_, _14670_);
  or (_26048_, _26047_, _26046_);
  and (_26050_, _26048_, _14981_);
  nor (_26051_, _26048_, _14981_);
  nor (_26052_, _26051_, _26050_);
  nor (_26053_, _26052_, _15275_);
  and (_26054_, _26052_, _15275_);
  or (_26055_, _26054_, _26053_);
  not (_26056_, _26055_);
  nor (_26057_, _26056_, _08148_);
  and (_26058_, _26056_, _08148_);
  or (_26059_, _26058_, _26057_);
  nand (_26061_, _26059_, _08070_);
  nand (_26062_, _26061_, _24721_);
  not (_26063_, _14975_);
  nor (_26064_, _13749_, _09290_);
  and (_26065_, _13749_, _09290_);
  or (_26066_, _26065_, _26064_);
  nor (_26067_, _26066_, _13787_);
  and (_26068_, _26066_, _13787_);
  nor (_26069_, _26068_, _26067_);
  and (_26070_, _26069_, _14361_);
  nor (_26072_, _26069_, _14361_);
  nor (_26073_, _26072_, _26070_);
  nor (_26074_, _26073_, _14667_);
  and (_26075_, _26073_, _14667_);
  or (_26076_, _26075_, _26074_);
  and (_26077_, _26076_, _26063_);
  nor (_26078_, _26076_, _26063_);
  nor (_26079_, _26078_, _26077_);
  nor (_26080_, _26079_, _15272_);
  and (_26081_, _26079_, _15272_);
  or (_26083_, _26081_, _26080_);
  or (_26084_, _26083_, _08110_);
  nand (_26085_, _26083_, _08110_);
  and (_26086_, _26085_, _03359_);
  and (_26087_, _26086_, _26084_);
  or (_26088_, _26087_, _26062_);
  or (_26089_, _26088_, _26036_);
  nand (_26090_, _26089_, _24722_);
  not (_26091_, _03271_);
  nor (_26092_, _03761_, _02889_);
  and (_26093_, _26092_, _09718_);
  and (_26094_, _26093_, _26091_);
  nand (_26095_, _26094_, _26090_);
  or (_26096_, _26094_, _24717_);
  and (_26097_, _26096_, _04523_);
  and (_26098_, _26097_, _26095_);
  and (_26099_, _24717_, _04524_);
  or (_26100_, _26099_, _03927_);
  or (_26101_, _26100_, _26098_);
  or (_26102_, _24717_, _05809_);
  and (_26105_, _26102_, _03179_);
  and (_26106_, _26105_, _26101_);
  and (_26107_, _24920_, _03174_);
  or (_26108_, _26107_, _08155_);
  or (_26109_, _26108_, _26106_);
  not (_26110_, _08161_);
  and (_26111_, _13833_, _26110_);
  and (_26112_, _26111_, \oc8051_golden_model_1.ACC [3]);
  nor (_26113_, _26111_, \oc8051_golden_model_1.ACC [3]);
  nor (_26114_, _26113_, _26112_);
  and (_26116_, _26114_, _14684_);
  nor (_26117_, _26114_, _14684_);
  nor (_26118_, _26117_, _26116_);
  and (_26119_, _14991_, _06807_);
  nor (_26120_, _14991_, _06807_);
  nor (_26121_, _26120_, _26119_);
  nor (_26122_, _26121_, _26118_);
  and (_26123_, _26121_, _26118_);
  or (_26124_, _26123_, _26122_);
  nor (_26125_, _26124_, _08167_);
  and (_26127_, _26124_, _08167_);
  nor (_26128_, _26127_, _26125_);
  and (_26129_, _26128_, _08155_);
  nor (_26130_, _26129_, _08160_);
  and (_26131_, _26130_, _26109_);
  and (_26132_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_26133_, _26132_, _07462_);
  nand (_26134_, _26133_, _25971_);
  or (_26135_, _26133_, _25971_);
  and (_26136_, _26135_, _26134_);
  nand (_26138_, _26136_, _08160_);
  nand (_26139_, _26138_, _03936_);
  or (_26140_, _26139_, _26131_);
  and (_26141_, _26140_, _24719_);
  or (_26142_, _26141_, _02799_);
  nor (_26143_, _24776_, _03183_);
  and (_26144_, _03298_, _02498_);
  nor (_26145_, _26144_, _26143_);
  and (_26146_, _26145_, _26142_);
  and (_26147_, _26144_, _24717_);
  or (_26149_, _26147_, _03607_);
  or (_26150_, _26149_, _26146_);
  not (_26151_, _03607_);
  nor (_26152_, _24717_, _26151_);
  nor (_26153_, _26152_, _03608_);
  and (_26154_, _26153_, _26150_);
  and (_26155_, _24717_, _03608_);
  or (_26156_, _26155_, _03941_);
  or (_26157_, _26156_, _26154_);
  or (_26158_, _24717_, _06161_);
  and (_26160_, _26158_, _02888_);
  and (_26161_, _26160_, _26157_);
  not (_26162_, _14389_);
  nor (_26163_, _14695_, _26162_);
  and (_26164_, _14695_, _26162_);
  nor (_26165_, _26164_, _26163_);
  nor (_26166_, _26165_, _15300_);
  and (_26167_, _26165_, _15300_);
  nor (_26168_, _26167_, _26166_);
  not (_26169_, _26168_);
  nor (_26171_, _13773_, _13294_);
  and (_26172_, _13773_, _13294_);
  nor (_26173_, _26172_, _26171_);
  and (_26174_, _26173_, _14095_);
  nor (_26175_, _26173_, _14095_);
  nor (_26176_, _26175_, _26174_);
  and (_26177_, _26176_, _15003_);
  nor (_26178_, _26176_, _15003_);
  or (_26179_, _26178_, _26177_);
  and (_26180_, _26179_, _08180_);
  nor (_26182_, _26179_, _08180_);
  or (_26183_, _26182_, _26180_);
  nand (_26184_, _26183_, _26169_);
  or (_26185_, _26183_, _26169_);
  and (_26186_, _26185_, _02887_);
  and (_26187_, _26186_, _26184_);
  or (_26188_, _26187_, _26161_);
  and (_26189_, _26188_, _08178_);
  not (_26190_, _08185_);
  and (_26191_, _13833_, _26190_);
  and (_26193_, _26191_, _02625_);
  nor (_26194_, _26191_, _02625_);
  nor (_26195_, _26194_, _26193_);
  nor (_26196_, _26195_, _14700_);
  and (_26197_, _26195_, _14700_);
  or (_26198_, _26197_, _26196_);
  and (_26199_, _26198_, _15306_);
  nor (_26200_, _26198_, _15306_);
  nor (_26201_, _26200_, _26199_);
  not (_26202_, _26201_);
  nor (_26204_, _15008_, _08192_);
  and (_26205_, _15008_, _08192_);
  nor (_26206_, _26205_, _26204_);
  nand (_26207_, _26206_, _26202_);
  or (_26208_, _26206_, _26202_);
  and (_26209_, _26208_, _08177_);
  and (_26210_, _26209_, _26207_);
  or (_26211_, _26210_, _26189_);
  nor (_26212_, _08184_, _03036_);
  and (_26213_, _26212_, _22780_);
  and (_26215_, _26213_, _26211_);
  not (_26216_, _26213_);
  and (_26217_, _26216_, _24717_);
  or (_26218_, _26217_, _34659_);
  or (_26219_, _26218_, _26215_);
  or (_26220_, _34655_, \oc8051_golden_model_1.PSW [0]);
  and (_26221_, _26220_, _35796_);
  and (_35843_[0], _26221_, _26219_);
  or (_26222_, _10565_, _09779_);
  nor (_26223_, _04718_, \oc8051_golden_model_1.PSW [1]);
  nor (_26225_, _26223_, _07150_);
  and (_26226_, _26225_, _26222_);
  not (_26227_, _05316_);
  nor (_26228_, _10618_, _26227_);
  not (_26229_, \oc8051_golden_model_1.PSW [1]);
  nor (_26230_, _05316_, _26229_);
  or (_26231_, _26230_, _02986_);
  or (_26232_, _26231_, _26228_);
  and (_26233_, _10574_, _04718_);
  nor (_26234_, _26233_, _26223_);
  or (_26236_, _26234_, _03006_);
  and (_26237_, _04718_, _02543_);
  nor (_26238_, _26237_, _26223_);
  nand (_26239_, _26238_, _03845_);
  or (_26240_, _03845_, _26229_);
  and (_26241_, _26240_, _03006_);
  and (_26242_, _26241_, _26239_);
  nor (_26243_, _26242_, _02977_);
  and (_26244_, _26243_, _26236_);
  nor (_26245_, _04718_, _26229_);
  nor (_26247_, _09779_, _04020_);
  or (_26248_, _26247_, _26245_);
  and (_26249_, _26248_, _02946_);
  and (_26250_, _10569_, _05316_);
  or (_26251_, _26250_, _26230_);
  and (_26252_, _26251_, _02884_);
  or (_26253_, _26252_, _26249_);
  or (_26254_, _26253_, _02880_);
  or (_26255_, _26254_, _26244_);
  or (_26256_, _26238_, _02992_);
  and (_26258_, _26256_, _26255_);
  or (_26259_, _26258_, _02877_);
  and (_26260_, _10572_, _05316_);
  or (_26261_, _26260_, _26230_);
  or (_26262_, _26261_, _02987_);
  and (_26263_, _26262_, _06246_);
  and (_26264_, _26263_, _26259_);
  and (_26265_, _26250_, _10568_);
  or (_26266_, _26265_, _26230_);
  and (_26267_, _26266_, _02871_);
  or (_26269_, _26267_, _02866_);
  or (_26270_, _26269_, _26264_);
  and (_26271_, _26270_, _26232_);
  or (_26272_, _26271_, _05535_);
  or (_26273_, _26248_, _02859_);
  and (_26274_, _26273_, _26272_);
  or (_26275_, _26274_, _02841_);
  and (_26276_, _06163_, _04718_);
  or (_26277_, _26245_, _02842_);
  or (_26278_, _26277_, _26276_);
  and (_26280_, _26278_, _02839_);
  and (_26281_, _26280_, _26275_);
  and (_26282_, _10674_, _04718_);
  or (_26283_, _26282_, _26245_);
  and (_26284_, _26283_, _02567_);
  or (_26285_, _26284_, _26281_);
  and (_26286_, _26285_, _03052_);
  or (_26287_, _10689_, _09779_);
  and (_26288_, _26287_, _03051_);
  nand (_26289_, _04718_, _03720_);
  and (_26291_, _26289_, _02834_);
  nor (_26292_, _26291_, _26288_);
  nor (_26293_, _26292_, _26223_);
  or (_26294_, _26293_, _26286_);
  and (_26295_, _26294_, _07150_);
  or (_26296_, _26295_, _26226_);
  and (_26297_, _26296_, _03138_);
  or (_26298_, _26245_, _05038_);
  and (_26299_, _26238_, _03137_);
  and (_26300_, _26299_, _26298_);
  or (_26302_, _10688_, _09779_);
  nor (_26303_, _26223_, _03023_);
  and (_26304_, _26303_, _26302_);
  or (_26305_, _26304_, _26300_);
  or (_26306_, _26305_, _26297_);
  and (_26307_, _26306_, _03144_);
  nand (_26308_, _26237_, _05037_);
  nor (_26309_, _26223_, _07161_);
  and (_26310_, _26309_, _26308_);
  or (_26311_, _26310_, _03174_);
  or (_26313_, _26289_, _05038_);
  nor (_26314_, _26223_, _03043_);
  and (_26315_, _26314_, _26313_);
  or (_26316_, _26315_, _26311_);
  or (_26317_, _26316_, _26307_);
  or (_26318_, _26234_, _03179_);
  and (_26319_, _26318_, _03183_);
  and (_26320_, _26319_, _26317_);
  and (_26321_, _26261_, _02799_);
  or (_26322_, _26321_, _02887_);
  or (_26324_, _26322_, _26320_);
  or (_26325_, _26245_, _02888_);
  or (_26326_, _26325_, _26233_);
  and (_26327_, _26326_, _26324_);
  or (_26328_, _26327_, _34659_);
  or (_26329_, _34655_, \oc8051_golden_model_1.PSW [1]);
  and (_26330_, _26329_, _35796_);
  and (_35843_[1], _26330_, _26328_);
  not (_26331_, _07190_);
  nor (_26332_, _07224_, _26331_);
  and (_26334_, _07224_, _07191_);
  or (_26335_, _26334_, _26332_);
  and (_26336_, _26335_, _10153_);
  not (_26337_, \oc8051_golden_model_1.PSW [2]);
  nor (_26338_, _04718_, _26337_);
  not (_26339_, _26338_);
  and (_26340_, _26339_, _05134_);
  and (_26341_, _04718_, _05693_);
  nor (_26342_, _26341_, _26338_);
  or (_26343_, _26342_, _03023_);
  or (_26345_, _26343_, _26340_);
  or (_26346_, _09779_, _04449_);
  and (_26347_, _26346_, _26339_);
  and (_26348_, _26347_, _05535_);
  nor (_26349_, _07326_, _05810_);
  nor (_26350_, _26349_, \oc8051_golden_model_1.ACC [7]);
  and (_26351_, _26349_, \oc8051_golden_model_1.ACC [7]);
  nor (_26352_, _26351_, _26350_);
  not (_26353_, _26352_);
  or (_26354_, _26353_, _10058_);
  nand (_26356_, _26353_, _10058_);
  and (_26357_, _26356_, _26354_);
  nand (_26358_, _26357_, _07396_);
  or (_26359_, _26357_, _07396_);
  and (_26360_, _26359_, _26358_);
  and (_26361_, _26360_, _07397_);
  and (_26362_, _10043_, _07239_);
  nor (_26363_, _10043_, _07239_);
  or (_26364_, _26363_, _26362_);
  and (_26365_, _26364_, _07531_);
  nor (_26367_, _26364_, _07531_);
  or (_26368_, _26367_, _26365_);
  or (_26369_, _26368_, _07399_);
  nor (_26370_, _10788_, _09779_);
  nor (_26371_, _26370_, _26338_);
  and (_26372_, _26371_, _02948_);
  and (_26373_, _04718_, \oc8051_golden_model_1.ACC [2]);
  nor (_26374_, _26373_, _26338_);
  or (_26375_, _26374_, _04194_);
  or (_26376_, _03845_, _26337_);
  and (_26378_, _26376_, _03006_);
  and (_26379_, _26378_, _26375_);
  or (_26380_, _26379_, _02977_);
  or (_26381_, _26380_, _26372_);
  or (_26382_, _26347_, _07474_);
  nor (_26383_, _05316_, _26337_);
  not (_26384_, _26383_);
  nand (_26385_, _10792_, _05316_);
  and (_26386_, _26385_, _26384_);
  or (_26387_, _26386_, _02934_);
  and (_26389_, _26387_, _26382_);
  and (_26390_, _26389_, _02992_);
  and (_26391_, _26390_, _26381_);
  and (_26392_, _26374_, _02880_);
  or (_26393_, _26392_, _26391_);
  and (_26394_, _26393_, _02987_);
  and (_26395_, _10773_, _05316_);
  nor (_26396_, _26395_, _26383_);
  and (_26397_, _26396_, _02877_);
  or (_26398_, _26397_, _02871_);
  or (_26400_, _26398_, _26394_);
  and (_26401_, _26384_, _09939_);
  or (_26402_, _26401_, _06246_);
  or (_26403_, _26402_, _26386_);
  and (_26404_, _26403_, _06258_);
  and (_26405_, _26404_, _26400_);
  or (_26406_, _12609_, _12499_);
  or (_26407_, _26406_, _12717_);
  or (_26408_, _26407_, _12831_);
  or (_26409_, _26408_, _12946_);
  or (_26411_, _26409_, _13059_);
  or (_26412_, _26411_, _06769_);
  nor (_26413_, _26412_, _13174_);
  or (_26414_, _26413_, _07400_);
  or (_26415_, _26414_, _26405_);
  and (_26416_, _26415_, _07507_);
  and (_26417_, _26416_, _26369_);
  or (_26418_, _26417_, _02979_);
  or (_26419_, _26418_, _26361_);
  nor (_26420_, _07642_, \oc8051_golden_model_1.ACC [7]);
  and (_26422_, _07642_, \oc8051_golden_model_1.ACC [7]);
  or (_26423_, _26422_, _26420_);
  nor (_26424_, _26423_, _09795_);
  and (_26425_, _26423_, _09795_);
  or (_26426_, _26425_, _26424_);
  or (_26427_, _26426_, _07717_);
  nand (_26428_, _26426_, _07717_);
  and (_26429_, _26428_, _26427_);
  or (_26430_, _26429_, _02991_);
  and (_26431_, _26430_, _07541_);
  and (_26433_, _26431_, _26419_);
  nor (_26434_, _07725_, _10175_);
  nor (_26435_, _07726_, \oc8051_golden_model_1.ACC [7]);
  nor (_26436_, _26435_, _26434_);
  not (_26437_, _26436_);
  or (_26438_, _26437_, _10072_);
  nand (_26439_, _26437_, _10072_);
  and (_26440_, _26439_, _26438_);
  nand (_26441_, _26440_, _07799_);
  or (_26442_, _26440_, _07799_);
  and (_26444_, _26442_, _26441_);
  and (_26445_, _26444_, _07540_);
  or (_26446_, _26445_, _02866_);
  or (_26447_, _26446_, _26433_);
  or (_26448_, _10825_, _26227_);
  and (_26449_, _26448_, _26384_);
  or (_26450_, _26449_, _02986_);
  and (_26451_, _26450_, _02859_);
  and (_26452_, _26451_, _26447_);
  or (_26453_, _26452_, _26348_);
  and (_26455_, _26453_, _02842_);
  or (_26456_, _06036_, _09779_);
  nor (_26457_, _26338_, _02842_);
  and (_26458_, _26457_, _26456_);
  or (_26459_, _26458_, _02567_);
  or (_26460_, _26459_, _26455_);
  or (_26461_, _10881_, _09779_);
  and (_26462_, _26461_, _26339_);
  or (_26463_, _26462_, _02839_);
  and (_26464_, _26463_, _06792_);
  and (_26466_, _26464_, _26460_);
  nand (_26467_, _06804_, _06798_);
  and (_26468_, _26467_, _06786_);
  or (_26469_, _26468_, _26466_);
  and (_26470_, _26469_, _07140_);
  and (_26471_, _26342_, _02834_);
  or (_26472_, _26471_, _03051_);
  or (_26473_, _26472_, _26470_);
  nand (_26474_, _10770_, _04718_);
  nor (_26475_, _26338_, _03148_);
  and (_26477_, _26475_, _26474_);
  or (_26478_, _26477_, _03149_);
  and (_26479_, _26478_, _26473_);
  nand (_26480_, _10766_, _04718_);
  nor (_26481_, _26338_, _07150_);
  and (_26482_, _26481_, _26480_);
  or (_26483_, _26482_, _03022_);
  or (_26484_, _26483_, _26479_);
  and (_26485_, _26484_, _26345_);
  or (_26486_, _26485_, _03137_);
  or (_26488_, _26374_, _06213_);
  or (_26489_, _26488_, _26340_);
  and (_26490_, _26489_, _03043_);
  and (_26491_, _26490_, _26486_);
  or (_26492_, _10768_, _09779_);
  nor (_26493_, _26338_, _03043_);
  and (_26494_, _26493_, _26492_);
  or (_26495_, _26494_, _03143_);
  or (_26496_, _26495_, _26491_);
  or (_26497_, _10765_, _09779_);
  and (_26499_, _26497_, _26339_);
  or (_26500_, _26499_, _07161_);
  and (_26501_, _26500_, _07234_);
  and (_26502_, _26501_, _26496_);
  and (_26503_, _07238_, \oc8051_golden_model_1.ACC [7]);
  nor (_26504_, _07238_, \oc8051_golden_model_1.ACC [7]);
  nor (_26505_, _26504_, _10126_);
  nor (_26506_, _26505_, _26503_);
  nand (_26507_, _26506_, _07307_);
  and (_26508_, _26503_, _07304_);
  nor (_26510_, _26508_, _07234_);
  and (_26511_, _26510_, _26507_);
  or (_26512_, _26511_, _26502_);
  nand (_26513_, _26512_, _07936_);
  and (_26514_, _26352_, _10132_);
  nor (_26515_, _26514_, _26351_);
  and (_26516_, _26515_, _07960_);
  and (_26517_, _26351_, _07957_);
  or (_26518_, _26517_, _07936_);
  or (_26519_, _26518_, _26516_);
  and (_26521_, _26519_, _03134_);
  and (_26522_, _26521_, _26513_);
  and (_26523_, _26422_, _07988_);
  not (_26524_, _10138_);
  nor (_26525_, _26423_, _26524_);
  nor (_26526_, _26525_, _26422_);
  and (_26527_, _26526_, _07991_);
  or (_26528_, _26527_, _26523_);
  and (_26529_, _26528_, _03133_);
  or (_26530_, _26529_, _07964_);
  or (_26532_, _26530_, _26522_);
  and (_26533_, _26434_, _08019_);
  and (_26534_, _26436_, _10144_);
  nor (_26535_, _26534_, _26434_);
  or (_26536_, _26535_, _07997_);
  and (_26537_, _26536_, _08023_);
  or (_26538_, _26537_, _26533_);
  and (_26539_, _26538_, _07189_);
  and (_26540_, _26539_, _26532_);
  or (_26541_, _26540_, _26336_);
  and (_26542_, _26541_, _21293_);
  or (_26543_, _08063_, _07854_);
  not (_26544_, _10161_);
  or (_26545_, _26544_, _08062_);
  and (_26546_, _26545_, _07185_);
  and (_26547_, _26546_, _26543_);
  or (_26548_, _08107_, _08071_);
  and (_26549_, _26548_, _10171_);
  nand (_26550_, _08145_, _10175_);
  and (_26551_, _26550_, _10177_);
  or (_26554_, _26551_, _03174_);
  or (_26555_, _26554_, _26549_);
  or (_26556_, _26555_, _26547_);
  or (_26557_, _26556_, _26542_);
  nand (_26558_, _26371_, _03174_);
  and (_26559_, _26558_, _03183_);
  and (_26560_, _26559_, _26557_);
  nor (_26561_, _26396_, _03183_);
  or (_26562_, _26561_, _02887_);
  or (_26563_, _26562_, _26560_);
  and (_26565_, _10941_, _04718_);
  or (_26566_, _26565_, _26338_);
  or (_26567_, _26566_, _02888_);
  and (_26568_, _26567_, _26563_);
  or (_26569_, _26568_, _34659_);
  or (_26570_, _34655_, \oc8051_golden_model_1.PSW [2]);
  and (_26571_, _26570_, _35796_);
  and (_35843_[2], _26571_, _26569_);
  nor (_26572_, _04718_, _02974_);
  nor (_26573_, _09779_, _04275_);
  or (_26575_, _26573_, _26572_);
  or (_26576_, _26575_, _02859_);
  nor (_26577_, _10973_, _26227_);
  nor (_26578_, _05316_, _02974_);
  or (_26579_, _26578_, _02986_);
  or (_26580_, _26579_, _26577_);
  nor (_26581_, _10983_, _09779_);
  or (_26582_, _26581_, _26572_);
  or (_26583_, _26582_, _03006_);
  and (_26584_, _04718_, \oc8051_golden_model_1.ACC [3]);
  nor (_26586_, _26584_, _26572_);
  or (_26587_, _26586_, _04194_);
  or (_26588_, _03845_, _02974_);
  and (_26589_, _26588_, _03006_);
  and (_26590_, _26589_, _26587_);
  nor (_26591_, _26590_, _02977_);
  and (_26592_, _26591_, _26583_);
  and (_26593_, _26575_, _02946_);
  and (_26594_, _10976_, _05316_);
  or (_26595_, _26594_, _26578_);
  and (_26597_, _26595_, _02884_);
  or (_26598_, _26597_, _26593_);
  or (_26599_, _26598_, _02880_);
  or (_26600_, _26599_, _26592_);
  nand (_26601_, _26586_, _02880_);
  and (_26602_, _26601_, _26600_);
  or (_26603_, _26602_, _02877_);
  and (_26604_, _10979_, _05316_);
  or (_26605_, _26604_, _26578_);
  or (_26606_, _26605_, _02987_);
  and (_26608_, _26606_, _06246_);
  and (_26609_, _26608_, _26603_);
  or (_26610_, _26578_, _10975_);
  and (_26611_, _26610_, _02871_);
  and (_26612_, _26611_, _26595_);
  or (_26613_, _26612_, _02866_);
  or (_26614_, _26613_, _26609_);
  and (_26615_, _26614_, _26580_);
  or (_26616_, _26615_, _05535_);
  and (_26617_, _26616_, _26576_);
  or (_26619_, _26617_, _02841_);
  and (_26620_, _06166_, _04718_);
  or (_26621_, _26572_, _02842_);
  or (_26622_, _26621_, _26620_);
  and (_26623_, _26622_, _02839_);
  and (_26624_, _26623_, _26619_);
  nor (_26625_, _11076_, _09779_);
  or (_26626_, _26572_, _26625_);
  and (_26627_, _26626_, _02567_);
  or (_26628_, _26627_, _26624_);
  or (_26630_, _26628_, _08207_);
  and (_26631_, _10968_, _04718_);
  or (_26632_, _26572_, _07139_);
  or (_26633_, _26632_, _26631_);
  and (_26634_, _04718_, _05654_);
  or (_26635_, _26634_, _26572_);
  or (_26636_, _26635_, _07140_);
  and (_26637_, _26636_, _07150_);
  and (_26638_, _26637_, _26633_);
  and (_26639_, _26638_, _26630_);
  and (_26641_, _10964_, _04718_);
  or (_26642_, _26641_, _26572_);
  and (_26643_, _26642_, _03148_);
  or (_26644_, _26643_, _26639_);
  and (_26645_, _26644_, _03138_);
  or (_26646_, _26572_, _04993_);
  nor (_26647_, _26586_, _06213_);
  and (_26648_, _26635_, _03022_);
  or (_26649_, _26648_, _26647_);
  and (_26650_, _26649_, _26646_);
  or (_26652_, _26650_, _03042_);
  or (_26653_, _26652_, _26645_);
  nor (_26654_, _10967_, _09779_);
  or (_26655_, _26572_, _03043_);
  or (_26656_, _26655_, _26654_);
  and (_26657_, _26656_, _07161_);
  and (_26658_, _26657_, _26653_);
  nor (_26659_, _10962_, _09779_);
  or (_26660_, _26659_, _26572_);
  and (_26661_, _26660_, _03143_);
  or (_26663_, _26661_, _03174_);
  or (_26664_, _26663_, _26658_);
  or (_26665_, _26582_, _03179_);
  and (_26666_, _26665_, _03183_);
  and (_26667_, _26666_, _26664_);
  and (_26668_, _26605_, _02799_);
  or (_26669_, _26668_, _02887_);
  or (_26670_, _26669_, _26667_);
  and (_26671_, _11136_, _04718_);
  or (_26672_, _26572_, _02888_);
  or (_26674_, _26672_, _26671_);
  and (_26675_, _26674_, _26670_);
  or (_26676_, _26675_, _34659_);
  or (_26677_, _34655_, \oc8051_golden_model_1.PSW [3]);
  and (_26678_, _26677_, _35796_);
  and (_35843_[3], _26678_, _26676_);
  not (_26679_, \oc8051_golden_model_1.PSW [4]);
  nor (_26680_, _04718_, _26679_);
  nor (_26681_, _05192_, _09779_);
  or (_26682_, _26681_, _26680_);
  or (_26684_, _26682_, _02859_);
  nor (_26685_, _05316_, _26679_);
  and (_26686_, _11167_, _05316_);
  or (_26687_, _26686_, _26685_);
  or (_26688_, _26685_, _11201_);
  and (_26689_, _26688_, _02871_);
  and (_26690_, _26689_, _26687_);
  nor (_26691_, _11184_, _09779_);
  or (_26692_, _26691_, _26680_);
  or (_26693_, _26692_, _03006_);
  and (_26695_, _04718_, \oc8051_golden_model_1.ACC [4]);
  nor (_26696_, _26695_, _26680_);
  or (_26697_, _26696_, _04194_);
  or (_26698_, _03845_, _26679_);
  and (_26699_, _26698_, _03006_);
  and (_26700_, _26699_, _26697_);
  nor (_26701_, _26700_, _02977_);
  and (_26702_, _26701_, _26693_);
  and (_26703_, _26682_, _02946_);
  and (_26704_, _26687_, _02884_);
  or (_26707_, _26704_, _26703_);
  or (_26708_, _26707_, _02880_);
  or (_26709_, _26708_, _26702_);
  nand (_26710_, _26696_, _02880_);
  and (_26711_, _26710_, _26709_);
  or (_26712_, _26711_, _02877_);
  and (_26713_, _11165_, _05316_);
  or (_26714_, _26713_, _26685_);
  or (_26715_, _26714_, _02987_);
  and (_26716_, _26715_, _06246_);
  and (_26718_, _26716_, _26712_);
  or (_26719_, _26718_, _26690_);
  and (_26720_, _26719_, _02986_);
  nor (_26721_, _11163_, _26227_);
  or (_26722_, _26721_, _26685_);
  and (_26723_, _26722_, _02866_);
  or (_26724_, _26723_, _05535_);
  or (_26725_, _26724_, _26720_);
  and (_26726_, _26725_, _26684_);
  or (_26727_, _26726_, _02841_);
  and (_26729_, _06171_, _04718_);
  or (_26730_, _26680_, _02842_);
  or (_26731_, _26730_, _26729_);
  and (_26732_, _26731_, _02839_);
  and (_26733_, _26732_, _26727_);
  nor (_26734_, _11271_, _09779_);
  or (_26735_, _26734_, _26680_);
  and (_26736_, _26735_, _02567_);
  or (_26737_, _26736_, _26733_);
  or (_26738_, _26737_, _08207_);
  and (_26740_, _11158_, _04718_);
  or (_26741_, _26680_, _07139_);
  or (_26742_, _26741_, _26740_);
  and (_26743_, _05618_, _04718_);
  or (_26744_, _26743_, _26680_);
  or (_26745_, _26744_, _07140_);
  and (_26746_, _26745_, _07150_);
  and (_26747_, _26746_, _26742_);
  and (_26748_, _26747_, _26738_);
  and (_26749_, _11154_, _04718_);
  or (_26751_, _26749_, _26680_);
  and (_26752_, _26751_, _03148_);
  or (_26753_, _26752_, _26748_);
  and (_26754_, _26753_, _03138_);
  or (_26755_, _26680_, _05240_);
  nor (_26756_, _26696_, _06213_);
  and (_26757_, _26744_, _03022_);
  or (_26758_, _26757_, _26756_);
  and (_26759_, _26758_, _26755_);
  or (_26760_, _26759_, _03042_);
  or (_26762_, _26760_, _26754_);
  nor (_26763_, _11157_, _09779_);
  or (_26764_, _26680_, _03043_);
  or (_26765_, _26764_, _26763_);
  and (_26766_, _26765_, _07161_);
  and (_26767_, _26766_, _26762_);
  nor (_26768_, _11152_, _09779_);
  or (_26769_, _26768_, _26680_);
  and (_26770_, _26769_, _03143_);
  or (_26771_, _26770_, _03174_);
  or (_26773_, _26771_, _26767_);
  or (_26774_, _26692_, _03179_);
  and (_26775_, _26774_, _03183_);
  and (_26776_, _26775_, _26773_);
  and (_26777_, _26714_, _02799_);
  or (_26778_, _26777_, _02887_);
  or (_26779_, _26778_, _26776_);
  and (_26780_, _11338_, _04718_);
  or (_26781_, _26680_, _02888_);
  or (_26782_, _26781_, _26780_);
  and (_26784_, _26782_, _26779_);
  or (_26785_, _26784_, _34659_);
  or (_26786_, _34655_, \oc8051_golden_model_1.PSW [4]);
  and (_26787_, _26786_, _35796_);
  and (_35843_[4], _26787_, _26785_);
  not (_26788_, \oc8051_golden_model_1.PSW [5]);
  nor (_26789_, _04718_, _26788_);
  nor (_26790_, _11380_, _09779_);
  or (_26791_, _26790_, _26789_);
  or (_26792_, _26791_, _03006_);
  and (_26794_, _04718_, \oc8051_golden_model_1.ACC [5]);
  nor (_26795_, _26794_, _26789_);
  or (_26796_, _26795_, _04194_);
  or (_26797_, _03845_, _26788_);
  and (_26798_, _26797_, _03006_);
  and (_26799_, _26798_, _26796_);
  nor (_26800_, _26799_, _02977_);
  and (_26801_, _26800_, _26792_);
  nor (_26802_, _04894_, _09779_);
  or (_26803_, _26802_, _26789_);
  and (_26805_, _26803_, _02946_);
  nor (_26806_, _05316_, _26788_);
  and (_26807_, _11365_, _05316_);
  or (_26808_, _26807_, _26806_);
  and (_26809_, _26808_, _02884_);
  or (_26810_, _26809_, _26805_);
  or (_26811_, _26810_, _02880_);
  or (_26812_, _26811_, _26801_);
  nand (_26813_, _26795_, _02880_);
  and (_26814_, _26813_, _26812_);
  or (_26816_, _26814_, _02877_);
  and (_26817_, _11363_, _05316_);
  or (_26818_, _26817_, _26806_);
  or (_26819_, _26818_, _02987_);
  and (_26820_, _26819_, _06246_);
  and (_26821_, _26820_, _26816_);
  and (_26822_, _11398_, _05316_);
  or (_26823_, _26822_, _26806_);
  and (_26824_, _26823_, _02871_);
  or (_26825_, _26824_, _26821_);
  and (_26827_, _26825_, _02986_);
  nor (_26828_, _11361_, _26227_);
  or (_26829_, _26828_, _26806_);
  and (_26830_, _26829_, _02866_);
  or (_26831_, _26830_, _05535_);
  or (_26832_, _26831_, _26827_);
  or (_26833_, _26803_, _02859_);
  and (_26834_, _26833_, _26832_);
  or (_26835_, _26834_, _02841_);
  and (_26836_, _06170_, _04718_);
  or (_26837_, _26789_, _02842_);
  or (_26838_, _26837_, _26836_);
  and (_26839_, _26838_, _02839_);
  and (_26840_, _26839_, _26835_);
  nor (_26841_, _11467_, _09779_);
  or (_26842_, _26841_, _26789_);
  and (_26843_, _26842_, _02567_);
  or (_26844_, _26843_, _08207_);
  or (_26845_, _26844_, _26840_);
  and (_26846_, _11482_, _04718_);
  or (_26849_, _26789_, _07139_);
  or (_26850_, _26849_, _26846_);
  and (_26851_, _05671_, _04718_);
  or (_26852_, _26851_, _26789_);
  or (_26853_, _26852_, _07140_);
  and (_26854_, _26853_, _07150_);
  and (_26855_, _26854_, _26850_);
  and (_26856_, _26855_, _26845_);
  and (_26857_, _11356_, _04718_);
  or (_26858_, _26857_, _26789_);
  and (_26860_, _26858_, _03148_);
  or (_26861_, _26860_, _26856_);
  and (_26862_, _26861_, _03138_);
  or (_26863_, _26789_, _04945_);
  nor (_26864_, _26795_, _06213_);
  and (_26865_, _26852_, _03022_);
  or (_26866_, _26865_, _26864_);
  and (_26867_, _26866_, _26863_);
  or (_26868_, _26867_, _03042_);
  or (_26869_, _26868_, _26862_);
  nor (_26871_, _11480_, _09779_);
  or (_26872_, _26789_, _03043_);
  or (_26873_, _26872_, _26871_);
  and (_26874_, _26873_, _07161_);
  and (_26875_, _26874_, _26869_);
  nor (_26876_, _11355_, _09779_);
  or (_26877_, _26876_, _26789_);
  and (_26878_, _26877_, _03143_);
  or (_26879_, _26878_, _03174_);
  or (_26880_, _26879_, _26875_);
  or (_26882_, _26791_, _03179_);
  and (_26883_, _26882_, _03183_);
  and (_26884_, _26883_, _26880_);
  and (_26885_, _26818_, _02799_);
  or (_26886_, _26885_, _02887_);
  or (_26887_, _26886_, _26884_);
  and (_26888_, _11541_, _04718_);
  or (_26889_, _26789_, _02888_);
  or (_26890_, _26889_, _26888_);
  and (_26891_, _26890_, _26887_);
  or (_26893_, _26891_, _34659_);
  or (_26894_, _34655_, \oc8051_golden_model_1.PSW [5]);
  and (_26895_, _26894_, _35796_);
  and (_35843_[5], _26895_, _26893_);
  or (_26896_, _08101_, _03166_);
  and (_26897_, _26896_, _08117_);
  nor (_26898_, _04718_, _14153_);
  nor (_26899_, _04790_, _09779_);
  or (_26900_, _26899_, _26898_);
  or (_26901_, _26900_, _02859_);
  or (_26903_, _07389_, _07344_);
  or (_26904_, _26903_, _07507_);
  nor (_26905_, _11567_, _09779_);
  or (_26906_, _26905_, _26898_);
  or (_26907_, _26906_, _03006_);
  and (_26908_, _04718_, \oc8051_golden_model_1.ACC [6]);
  nor (_26909_, _26908_, _26898_);
  or (_26910_, _26909_, _04194_);
  or (_26911_, _03845_, _14153_);
  and (_26912_, _26911_, _03006_);
  and (_26914_, _26912_, _26910_);
  nor (_26915_, _26914_, _02977_);
  and (_26916_, _26915_, _26907_);
  and (_26917_, _26900_, _02946_);
  nor (_26918_, _05316_, _14153_);
  and (_26919_, _11564_, _05316_);
  or (_26920_, _26919_, _26918_);
  and (_26921_, _26920_, _02884_);
  or (_26922_, _26921_, _26917_);
  or (_26923_, _26922_, _02880_);
  or (_26925_, _26923_, _26916_);
  nand (_26926_, _26909_, _02880_);
  and (_26927_, _26926_, _26925_);
  or (_26928_, _26927_, _02877_);
  and (_26929_, _11562_, _05316_);
  or (_26930_, _26929_, _26918_);
  or (_26931_, _26930_, _02987_);
  and (_26932_, _26931_, _06246_);
  and (_26933_, _26932_, _26928_);
  or (_26934_, _26918_, _11596_);
  and (_26936_, _26934_, _02871_);
  and (_26937_, _26936_, _26920_);
  or (_26938_, _26937_, _07400_);
  or (_26939_, _26938_, _26933_);
  or (_26940_, _07259_, _07399_);
  or (_26941_, _26940_, _07524_);
  and (_26942_, _26941_, _26939_);
  or (_26943_, _26942_, _07397_);
  and (_26944_, _26943_, _02991_);
  and (_26945_, _26944_, _26904_);
  or (_26946_, _07611_, _07540_);
  or (_26947_, _26946_, _07710_);
  and (_26948_, _26947_, _09325_);
  or (_26949_, _26948_, _26945_);
  or (_26950_, _07723_, _07541_);
  or (_26951_, _26950_, _07792_);
  and (_26952_, _26951_, _02986_);
  and (_26953_, _26952_, _26949_);
  nor (_26954_, _11614_, _26227_);
  or (_26955_, _26954_, _26918_);
  and (_26958_, _26955_, _02866_);
  or (_26959_, _26958_, _05535_);
  or (_26960_, _26959_, _26953_);
  and (_26961_, _26960_, _26901_);
  or (_26962_, _26961_, _02841_);
  and (_26963_, _06162_, _04718_);
  or (_26964_, _26898_, _02842_);
  or (_26965_, _26964_, _26963_);
  and (_26966_, _26965_, _02839_);
  and (_26967_, _26966_, _26962_);
  nor (_26969_, _11671_, _09779_);
  or (_26970_, _26969_, _26898_);
  and (_26971_, _26970_, _02567_);
  or (_26972_, _26971_, _08207_);
  or (_26973_, _26972_, _26967_);
  and (_26974_, _11560_, _04718_);
  or (_26975_, _26898_, _07139_);
  or (_26976_, _26975_, _26974_);
  and (_26977_, _11678_, _04718_);
  or (_26978_, _26977_, _26898_);
  or (_26980_, _26978_, _07140_);
  and (_26981_, _26980_, _07150_);
  and (_26982_, _26981_, _26976_);
  and (_26983_, _26982_, _26973_);
  and (_26984_, _11556_, _04718_);
  or (_26985_, _26984_, _26898_);
  and (_26986_, _26985_, _03148_);
  or (_26987_, _26986_, _26983_);
  and (_26988_, _26987_, _03138_);
  or (_26989_, _26898_, _04838_);
  nor (_26991_, _26909_, _06213_);
  and (_26992_, _26978_, _03022_);
  or (_26993_, _26992_, _26991_);
  and (_26994_, _26993_, _26989_);
  or (_26995_, _26994_, _03042_);
  or (_26996_, _26995_, _26988_);
  nor (_26997_, _11558_, _09779_);
  or (_26998_, _26997_, _26898_);
  or (_26999_, _26998_, _03043_);
  and (_27000_, _26999_, _26996_);
  or (_27002_, _27000_, _03143_);
  nor (_27003_, _11555_, _09779_);
  or (_27004_, _26898_, _07161_);
  nor (_27005_, _27004_, _27003_);
  nor (_27006_, _27005_, _03282_);
  and (_27007_, _27006_, _27002_);
  not (_27008_, _07259_);
  nand (_27009_, _07298_, _27008_);
  and (_27010_, _27009_, _03282_);
  or (_27011_, _27010_, _27007_);
  and (_27013_, _27011_, _03280_);
  and (_27014_, _27009_, _03279_);
  nor (_27015_, _27014_, _27013_);
  nor (_27016_, _27015_, _03277_);
  and (_27017_, _27009_, _03277_);
  nor (_27018_, _27017_, _27016_);
  or (_27019_, _27018_, _03730_);
  nand (_27020_, _27009_, _03730_);
  nand (_27021_, _27020_, _27019_);
  or (_27022_, _27021_, _03734_);
  and (_27024_, _02845_, _02527_);
  not (_27025_, _03734_);
  nor (_27026_, _27009_, _27025_);
  nor (_27027_, _27026_, _27024_);
  and (_27028_, _27027_, _27022_);
  and (_27029_, _03014_, _02527_);
  and (_27030_, _27009_, _27024_);
  or (_27031_, _27030_, _27029_);
  or (_27032_, _27031_, _27028_);
  not (_27033_, _27029_);
  not (_27035_, _07344_);
  nand (_27036_, _07951_, _27035_);
  or (_27037_, _27036_, _27033_);
  nand (_27038_, _27037_, _27032_);
  nor (_27039_, _27038_, _03556_);
  and (_27040_, _27036_, _03556_);
  or (_27041_, _27040_, _03133_);
  or (_27042_, _27041_, _27039_);
  nor (_27043_, _07611_, _03134_);
  nand (_27044_, _27043_, _07982_);
  and (_27046_, _27044_, _07997_);
  and (_27047_, _27046_, _27042_);
  not (_27048_, _07723_);
  nand (_27049_, _08013_, _27048_);
  and (_27050_, _27049_, _07964_);
  or (_27051_, _27050_, _10153_);
  or (_27052_, _27051_, _27047_);
  or (_27053_, _07218_, _07189_);
  and (_27054_, _27053_, _08031_);
  and (_27055_, _27054_, _27052_);
  and (_27057_, _08057_, _07185_);
  or (_27058_, _27057_, _03359_);
  or (_27059_, _27058_, _27055_);
  and (_27060_, _27059_, _26897_);
  and (_27061_, _08139_, _08070_);
  or (_27062_, _27061_, _03174_);
  or (_27063_, _27062_, _27060_);
  or (_27064_, _26906_, _03179_);
  and (_27065_, _27064_, _03183_);
  and (_27066_, _27065_, _27063_);
  and (_27068_, _26930_, _02799_);
  or (_27069_, _27068_, _02887_);
  or (_27070_, _27069_, _27066_);
  and (_27071_, _11744_, _04718_);
  or (_27072_, _26898_, _02888_);
  or (_27073_, _27072_, _27071_);
  and (_27074_, _27073_, _27070_);
  or (_27075_, _27074_, _34659_);
  or (_27076_, _34655_, \oc8051_golden_model_1.PSW [6]);
  and (_27077_, _27076_, _35796_);
  and (_35843_[6], _27077_, _27075_);
  and (_35841_[0], \oc8051_golden_model_1.PCON [0], _35796_);
  and (_35841_[1], \oc8051_golden_model_1.PCON [1], _35796_);
  and (_35841_[2], \oc8051_golden_model_1.PCON [2], _35796_);
  and (_35841_[3], \oc8051_golden_model_1.PCON [3], _35796_);
  and (_35841_[4], \oc8051_golden_model_1.PCON [4], _35796_);
  and (_35841_[5], \oc8051_golden_model_1.PCON [5], _35796_);
  and (_35841_[6], \oc8051_golden_model_1.PCON [6], _35796_);
  and (_35844_[0], \oc8051_golden_model_1.SBUF [0], _35796_);
  and (_35844_[1], \oc8051_golden_model_1.SBUF [1], _35796_);
  and (_35844_[2], \oc8051_golden_model_1.SBUF [2], _35796_);
  and (_35844_[3], \oc8051_golden_model_1.SBUF [3], _35796_);
  and (_35844_[4], \oc8051_golden_model_1.SBUF [4], _35796_);
  and (_35844_[5], \oc8051_golden_model_1.SBUF [5], _35796_);
  and (_35844_[6], \oc8051_golden_model_1.SBUF [6], _35796_);
  and (_35845_[0], \oc8051_golden_model_1.SCON [0], _35796_);
  and (_35845_[1], \oc8051_golden_model_1.SCON [1], _35796_);
  and (_35845_[2], \oc8051_golden_model_1.SCON [2], _35796_);
  and (_35845_[3], \oc8051_golden_model_1.SCON [3], _35796_);
  and (_35845_[4], \oc8051_golden_model_1.SCON [4], _35796_);
  and (_35845_[5], \oc8051_golden_model_1.SCON [5], _35796_);
  and (_35845_[6], \oc8051_golden_model_1.SCON [6], _35796_);
  nor (_27081_, _04638_, _02868_);
  nor (_27082_, _05085_, _10206_);
  or (_27083_, _27082_, _27081_);
  or (_27084_, _27083_, _03360_);
  or (_27085_, _10369_, _10206_);
  nor (_27086_, _04638_, \oc8051_golden_model_1.SP [0]);
  nor (_27087_, _27086_, _07150_);
  and (_27088_, _27087_, _27085_);
  or (_27090_, _10372_, _10206_);
  nor (_27091_, _27086_, _07139_);
  and (_27092_, _27091_, _27090_);
  and (_27093_, _06164_, _04638_);
  or (_27094_, _27081_, _02842_);
  or (_27095_, _27094_, _27093_);
  and (_27096_, _04638_, _03838_);
  or (_27097_, _27081_, _02859_);
  or (_27098_, _27097_, _27096_);
  and (_27099_, _27083_, _02948_);
  not (_27101_, _27086_);
  nand (_27102_, _04638_, _02696_);
  and (_27103_, _27102_, _27101_);
  and (_27104_, _27103_, _03845_);
  nor (_27105_, _03845_, _02868_);
  or (_27106_, _27105_, _27104_);
  and (_27107_, _27106_, _03006_);
  or (_27108_, _27107_, _02946_);
  or (_27109_, _27108_, _27099_);
  or (_27110_, _27086_, _07474_);
  or (_27112_, _27110_, _27096_);
  and (_27113_, _27112_, _27109_);
  or (_27114_, _27113_, _02880_);
  or (_27115_, _27103_, _02992_);
  and (_27116_, _27115_, _03962_);
  and (_27117_, _27116_, _27114_);
  nand (_27118_, _02859_, _03881_);
  or (_27119_, _27118_, _27117_);
  and (_27120_, _27119_, _27098_);
  or (_27121_, _27120_, _02841_);
  and (_27123_, _27121_, _02839_);
  and (_27124_, _27123_, _27095_);
  nand (_27125_, _10475_, _04638_);
  nor (_27126_, _27086_, _02839_);
  and (_27127_, _27126_, _27125_);
  or (_27128_, _27127_, _02834_);
  or (_27129_, _27128_, _27124_);
  nand (_27130_, _04638_, _03505_);
  and (_27131_, _27130_, _27101_);
  or (_27132_, _27131_, _07140_);
  and (_27134_, _27132_, _07139_);
  and (_27135_, _27134_, _27129_);
  or (_27136_, _27135_, _27092_);
  and (_27137_, _27136_, _07150_);
  or (_27138_, _27137_, _27088_);
  and (_27139_, _27138_, _03138_);
  nand (_27140_, _27103_, _03137_);
  nor (_27141_, _27140_, _27082_);
  nand (_27142_, _27131_, _03022_);
  nor (_27143_, _27142_, _27082_);
  or (_27144_, _27143_, _27141_);
  or (_27145_, _27144_, _27139_);
  and (_27146_, _27145_, _03144_);
  or (_27147_, _27102_, _05085_);
  nor (_27148_, _27086_, _07161_);
  and (_27149_, _27148_, _27147_);
  or (_27150_, _27130_, _05085_);
  nor (_27151_, _27086_, _03043_);
  and (_27152_, _27151_, _27150_);
  or (_27153_, _27152_, _03361_);
  or (_27156_, _27153_, _27149_);
  or (_27157_, _27156_, _27146_);
  and (_27158_, _27157_, _27084_);
  and (_27159_, _27158_, _34655_);
  nor (_27160_, \oc8051_golden_model_1.SP [0], rst);
  nor (_27161_, _27160_, _00000_);
  or (_35846_[0], _27161_, _27159_);
  nor (_27162_, _04638_, _03741_);
  and (_27163_, _10574_, _04638_);
  nor (_27164_, _27163_, _27162_);
  nor (_27166_, _27164_, _02888_);
  not (_27167_, _25962_);
  and (_27168_, _04638_, _02543_);
  nand (_27169_, _27168_, _05037_);
  nor (_27170_, _04638_, \oc8051_golden_model_1.SP [1]);
  nor (_27171_, _27170_, _07161_);
  and (_27172_, _27171_, _27169_);
  and (_27173_, _02530_, _03741_);
  and (_27174_, _02522_, _03741_);
  nor (_27175_, _10206_, _04020_);
  or (_27177_, _27162_, _02841_);
  nor (_27178_, _27177_, _27175_);
  nor (_27179_, _27178_, _02860_);
  nor (_27180_, _27170_, _27163_);
  nor (_27181_, _27180_, _03006_);
  nor (_27182_, _27168_, _27170_);
  and (_27183_, _27182_, _03845_);
  nor (_27184_, _03845_, _03741_);
  or (_27185_, _27184_, _27183_);
  and (_27186_, _27185_, _02603_);
  nor (_27188_, _02603_, \oc8051_golden_model_1.SP [1]);
  or (_27189_, _27188_, _27186_);
  nor (_27190_, _27189_, _02948_);
  nor (_27191_, _27190_, _27181_);
  and (_27192_, _27191_, _22534_);
  nor (_27193_, _02597_, \oc8051_golden_model_1.SP [1]);
  nor (_27194_, _27193_, _27192_);
  nor (_27195_, _04638_, _03957_);
  nor (_27196_, _27195_, _27175_);
  nor (_27197_, _27196_, _07474_);
  nor (_27199_, _27197_, _02880_);
  and (_27200_, _27199_, _27194_);
  nor (_27201_, _27182_, _02992_);
  nor (_27202_, _27201_, _02876_);
  not (_27203_, _27202_);
  nor (_27204_, _27203_, _27200_);
  or (_27205_, _27204_, _10219_);
  nor (_27206_, _27205_, _03961_);
  nor (_27207_, _04135_, _03741_);
  nor (_27208_, _27207_, _05535_);
  not (_27210_, _27208_);
  nor (_27211_, _27210_, _27206_);
  nor (_27212_, _27211_, _27179_);
  and (_27213_, _06163_, _04638_);
  nor (_27214_, _27162_, _02842_);
  not (_27215_, _27214_);
  nor (_27216_, _27215_, _27213_);
  nor (_27217_, _27216_, _02567_);
  not (_27218_, _27217_);
  nor (_27219_, _27218_, _27212_);
  and (_27221_, _10674_, _04638_);
  nor (_27222_, _27221_, _27162_);
  nor (_27223_, _27222_, _02839_);
  nor (_27224_, _27223_, _27219_);
  nor (_27225_, _27224_, _02834_);
  and (_27226_, _04638_, _03720_);
  not (_27227_, _27226_);
  nor (_27228_, _27170_, _07140_);
  and (_27229_, _27228_, _27227_);
  or (_27230_, _27229_, _27225_);
  and (_27232_, _27230_, _04131_);
  or (_27233_, _27232_, _27174_);
  and (_27234_, _27233_, _07139_);
  not (_27235_, _27170_);
  nor (_27236_, _10689_, _10206_);
  nor (_27237_, _27236_, _07139_);
  and (_27238_, _27237_, _27235_);
  nor (_27239_, _27238_, _27234_);
  nor (_27240_, _27239_, _03148_);
  nor (_27241_, _10565_, _10206_);
  nor (_27243_, _27241_, _07150_);
  and (_27244_, _27243_, _27235_);
  nor (_27245_, _27244_, _27240_);
  nor (_27246_, _27245_, _03022_);
  nor (_27247_, _10688_, _10206_);
  nor (_27248_, _27247_, _03023_);
  and (_27249_, _27248_, _27235_);
  nor (_27250_, _27249_, _27246_);
  nor (_27251_, _27250_, _09463_);
  nor (_27252_, _27162_, _05038_);
  nor (_27254_, _27252_, _06213_);
  and (_27255_, _27254_, _27182_);
  or (_27256_, _27255_, _27251_);
  nor (_27257_, _27256_, _27173_);
  nor (_27258_, _27257_, _03042_);
  and (_27259_, _27226_, _05037_);
  nor (_27260_, _27259_, _03043_);
  and (_27261_, _27260_, _27235_);
  or (_27262_, _27261_, _27258_);
  and (_27263_, _27262_, _07161_);
  nor (_27265_, _27263_, _27172_);
  nor (_27266_, _27265_, _27167_);
  nor (_27267_, _25962_, \oc8051_golden_model_1.SP [1]);
  nor (_27268_, _27267_, _02890_);
  not (_27269_, _27268_);
  nor (_27270_, _27269_, _27266_);
  nor (_27271_, _03722_, _03174_);
  not (_27272_, _27271_);
  nor (_27273_, _27272_, _27270_);
  and (_27274_, _03936_, _03179_);
  nor (_27276_, _27180_, _04150_);
  nor (_27277_, _27276_, _27274_);
  nor (_27278_, _27277_, _27273_);
  nor (_27279_, _03936_, _03741_);
  nor (_27280_, _27279_, _02887_);
  not (_27281_, _27280_);
  nor (_27282_, _27281_, _27278_);
  nor (_27283_, _27282_, _27166_);
  nor (_27284_, _27283_, _34659_);
  nor (_27285_, \oc8051_golden_model_1.SP [1], rst);
  nor (_27287_, _27285_, _00000_);
  or (_35846_[1], _27287_, _27284_);
  and (_27288_, _04548_, _02528_);
  nor (_27289_, _04638_, _03264_);
  and (_27290_, _10766_, _04638_);
  nor (_27291_, _27290_, _27289_);
  nor (_27292_, _27291_, _07150_);
  and (_27293_, _12112_, _02522_);
  nor (_27294_, _10206_, _04449_);
  or (_27295_, _27289_, _02859_);
  nor (_27297_, _27295_, _27294_);
  nor (_27298_, _10788_, _10206_);
  nor (_27299_, _27298_, _27289_);
  nor (_27300_, _27299_, _03006_);
  nor (_27301_, _12112_, _02603_);
  nor (_27302_, _03845_, _03264_);
  and (_27303_, _04638_, \oc8051_golden_model_1.ACC [2]);
  nor (_27304_, _27303_, _27289_);
  nor (_27305_, _27304_, _04194_);
  or (_27306_, _27305_, _27302_);
  and (_27308_, _27306_, _02603_);
  nor (_27309_, _27308_, _27301_);
  nor (_27310_, _27309_, _02948_);
  or (_27311_, _27310_, _04225_);
  nor (_27312_, _27311_, _27300_);
  nor (_27313_, _04548_, _02597_);
  nor (_27314_, _27313_, _27312_);
  and (_27315_, _27314_, _07474_);
  nor (_27316_, _05376_, _04638_);
  nor (_27317_, _27316_, _27294_);
  nor (_27319_, _27317_, _07474_);
  or (_27320_, _27319_, _27315_);
  and (_27321_, _27320_, _02992_);
  nor (_27322_, _27304_, _02992_);
  or (_27323_, _27322_, _27321_);
  and (_27324_, _27323_, _03962_);
  nor (_27325_, _27324_, _04394_);
  nor (_27326_, _27325_, _10219_);
  nor (_27327_, _12112_, _04135_);
  nor (_27328_, _27327_, _05535_);
  not (_27330_, _27328_);
  nor (_27331_, _27330_, _27326_);
  nor (_27332_, _27331_, _27297_);
  nor (_27333_, _27332_, _02841_);
  and (_27334_, _06167_, _04638_);
  nor (_27335_, _27289_, _02842_);
  not (_27336_, _27335_);
  nor (_27337_, _27336_, _27334_);
  or (_27338_, _27337_, _02567_);
  nor (_27339_, _27338_, _27333_);
  nor (_27341_, _10881_, _10206_);
  nor (_27342_, _27341_, _27289_);
  nor (_27343_, _27342_, _02839_);
  or (_27344_, _27343_, _02834_);
  or (_27345_, _27344_, _27339_);
  and (_27346_, _04638_, _05693_);
  nor (_27347_, _27346_, _27289_);
  nand (_27348_, _27347_, _02834_);
  and (_27349_, _27348_, _27345_);
  nor (_27350_, _27349_, _02522_);
  nor (_27352_, _27350_, _27293_);
  and (_27353_, _27352_, _07139_);
  and (_27354_, _10770_, _04638_);
  nor (_27355_, _27354_, _27289_);
  nor (_27356_, _27355_, _07139_);
  or (_27357_, _27356_, _27353_);
  and (_27358_, _27357_, _07150_);
  nor (_27359_, _27358_, _27292_);
  nor (_27360_, _27359_, _03022_);
  nor (_27361_, _27289_, _05135_);
  not (_27363_, _27361_);
  nor (_27364_, _27347_, _03023_);
  and (_27365_, _27364_, _27363_);
  nor (_27366_, _27365_, _27360_);
  nor (_27367_, _27366_, _09463_);
  and (_27368_, _04548_, _02530_);
  or (_27369_, _27361_, _06213_);
  nor (_27370_, _27369_, _27304_);
  or (_27371_, _27370_, _27368_);
  or (_27372_, _27371_, _03042_);
  nor (_27374_, _27372_, _27367_);
  nor (_27375_, _10768_, _10206_);
  nor (_27376_, _27375_, _27289_);
  and (_27377_, _27376_, _03042_);
  nor (_27378_, _27377_, _27374_);
  nor (_27379_, _27378_, _03143_);
  nor (_27380_, _10765_, _10206_);
  or (_27381_, _27289_, _07161_);
  nor (_27382_, _27381_, _27380_);
  or (_27383_, _27382_, _03155_);
  nor (_27385_, _27383_, _27379_);
  and (_27386_, _12112_, _03155_);
  or (_27387_, _27386_, _27385_);
  and (_27388_, _27387_, _05790_);
  or (_27389_, _27388_, _27288_);
  and (_27390_, _27389_, _02891_);
  and (_27391_, _12112_, _02890_);
  or (_27392_, _27391_, _03174_);
  nor (_27393_, _27392_, _27390_);
  and (_27394_, _27299_, _03174_);
  nor (_27396_, _27394_, _04150_);
  not (_27397_, _27396_);
  nor (_27398_, _27397_, _27393_);
  nor (_27399_, _12112_, _03936_);
  nor (_27400_, _27399_, _02887_);
  not (_27401_, _27400_);
  nor (_27402_, _27401_, _27398_);
  and (_27403_, _10941_, _04638_);
  nor (_27404_, _27403_, _27289_);
  and (_27405_, _27404_, _02887_);
  nor (_27406_, _27405_, _27402_);
  and (_27407_, _27406_, _34655_);
  nor (_27408_, \oc8051_golden_model_1.SP [2], rst);
  nor (_27409_, _27408_, _00000_);
  or (_35846_[2], _27409_, _27407_);
  nor (_27410_, _04638_, _05412_);
  and (_27411_, _11136_, _04638_);
  nor (_27412_, _27411_, _27410_);
  nor (_27413_, _27412_, _02888_);
  and (_27414_, _10964_, _04638_);
  nor (_27417_, _27414_, _27410_);
  nor (_27418_, _27417_, _07150_);
  and (_27419_, _11922_, _02522_);
  nor (_27420_, _10206_, _04275_);
  or (_27421_, _27410_, _02841_);
  nor (_27422_, _27421_, _27420_);
  nor (_27423_, _27422_, _02860_);
  and (_27424_, _04638_, \oc8051_golden_model_1.ACC [3]);
  nor (_27425_, _27424_, _27410_);
  nor (_27426_, _27425_, _04194_);
  nor (_27428_, _03845_, _05412_);
  or (_27429_, _27428_, _03849_);
  nor (_27430_, _27429_, _27426_);
  nor (_27431_, _04551_, _02603_);
  nor (_27432_, _27431_, _27430_);
  and (_27433_, _27432_, _03006_);
  nor (_27434_, _10983_, _10206_);
  nor (_27435_, _27434_, _27410_);
  nor (_27436_, _27435_, _03006_);
  or (_27437_, _27436_, _27433_);
  and (_27439_, _27437_, _02597_);
  nor (_27440_, _11922_, _02597_);
  or (_27441_, _27440_, _27439_);
  and (_27442_, _27441_, _07474_);
  nor (_27443_, _05417_, _04638_);
  nor (_27444_, _27443_, _27420_);
  nor (_27445_, _27444_, _07474_);
  or (_27446_, _27445_, _27442_);
  and (_27447_, _27446_, _02992_);
  nor (_27448_, _27425_, _02992_);
  or (_27450_, _27448_, _27447_);
  and (_27451_, _27450_, _03962_);
  or (_27452_, _27451_, _10219_);
  nor (_27453_, _27452_, _04313_);
  nor (_27454_, _04551_, _04135_);
  nor (_27455_, _27454_, _05535_);
  not (_27456_, _27455_);
  nor (_27457_, _27456_, _27453_);
  nor (_27458_, _27457_, _27423_);
  and (_27459_, _06166_, _04638_);
  nor (_27461_, _27410_, _02842_);
  not (_27462_, _27461_);
  nor (_27463_, _27462_, _27459_);
  or (_27464_, _27463_, _02567_);
  nor (_27465_, _27464_, _27458_);
  nor (_27466_, _11076_, _10206_);
  nor (_27467_, _27466_, _27410_);
  nor (_27468_, _27467_, _02839_);
  or (_27469_, _27468_, _02834_);
  or (_27470_, _27469_, _27465_);
  and (_27472_, _04638_, _05654_);
  nor (_27473_, _27472_, _27410_);
  nand (_27474_, _27473_, _02834_);
  and (_27475_, _27474_, _27470_);
  nor (_27476_, _27475_, _02522_);
  nor (_27477_, _27476_, _27419_);
  and (_27478_, _27477_, _07139_);
  and (_27479_, _10968_, _04638_);
  nor (_27480_, _27479_, _27410_);
  nor (_27481_, _27480_, _07139_);
  or (_27483_, _27481_, _27478_);
  and (_27484_, _27483_, _07150_);
  nor (_27485_, _27484_, _27418_);
  nor (_27486_, _27485_, _03022_);
  nor (_27487_, _27410_, _04993_);
  not (_27488_, _27487_);
  nor (_27489_, _27473_, _03023_);
  and (_27490_, _27489_, _27488_);
  nor (_27491_, _27490_, _27486_);
  nor (_27492_, _27491_, _09463_);
  and (_27494_, _04551_, _02530_);
  or (_27495_, _27487_, _06213_);
  nor (_27496_, _27495_, _27425_);
  or (_27497_, _27496_, _27494_);
  or (_27498_, _27497_, _03042_);
  nor (_27499_, _27498_, _27492_);
  nor (_27500_, _10967_, _10206_);
  nor (_27501_, _27500_, _27410_);
  and (_27502_, _27501_, _03042_);
  nor (_27503_, _27502_, _27499_);
  and (_27505_, _27503_, _07161_);
  nor (_27506_, _10962_, _10206_);
  nor (_27507_, _27506_, _27410_);
  nor (_27508_, _27507_, _07161_);
  or (_27509_, _27508_, _27505_);
  and (_27510_, _27509_, _20557_);
  nor (_27511_, _05414_, _05412_);
  nor (_27512_, _27511_, _05415_);
  nor (_27513_, _27512_, _20557_);
  or (_27514_, _27513_, _02528_);
  nor (_27516_, _27514_, _27510_);
  and (_27517_, _11922_, _02528_);
  nor (_27518_, _27517_, _27516_);
  and (_27519_, _27518_, _02891_);
  nor (_27520_, _27512_, _02891_);
  or (_27521_, _27520_, _27519_);
  and (_27522_, _27521_, _03179_);
  nor (_27523_, _27435_, _03179_);
  or (_27524_, _27523_, _04150_);
  nor (_27525_, _27524_, _27522_);
  nor (_27527_, _04551_, _03936_);
  nor (_27528_, _27527_, _02887_);
  not (_27529_, _27528_);
  nor (_27530_, _27529_, _27525_);
  nor (_27531_, _27530_, _27413_);
  nand (_27532_, _27531_, _34655_);
  or (_27533_, _34655_, \oc8051_golden_model_1.SP [3]);
  and (_27534_, _27533_, _35796_);
  and (_35846_[3], _27534_, _27532_);
  nor (_27535_, _04638_, _10243_);
  and (_27537_, _11338_, _04638_);
  nor (_27538_, _27537_, _27535_);
  nor (_27539_, _27538_, _02888_);
  and (_27540_, _11154_, _04638_);
  nor (_27541_, _27540_, _27535_);
  nor (_27542_, _27541_, _07150_);
  nor (_27543_, _05192_, _10206_);
  or (_27544_, _27535_, _02841_);
  nor (_27545_, _27544_, _27543_);
  nor (_27546_, _27545_, _02860_);
  nor (_27548_, _03845_, _10243_);
  and (_27549_, _04638_, \oc8051_golden_model_1.ACC [4]);
  nor (_27550_, _27549_, _27535_);
  nor (_27551_, _27550_, _04194_);
  or (_27552_, _27551_, _27548_);
  and (_27553_, _27552_, _02603_);
  nor (_27554_, _04219_, \oc8051_golden_model_1.SP [4]);
  nor (_27555_, _27554_, _10211_);
  not (_27556_, _27555_);
  nor (_27557_, _27556_, _02603_);
  nor (_27559_, _27557_, _27553_);
  nor (_27560_, _27559_, _02948_);
  nor (_27561_, _11184_, _10206_);
  nor (_27562_, _27561_, _27535_);
  nor (_27563_, _27562_, _03006_);
  or (_27564_, _27563_, _27560_);
  and (_27565_, _27564_, _02597_);
  nor (_27566_, _27556_, _02597_);
  or (_27567_, _27566_, _27565_);
  and (_27568_, _27567_, _07474_);
  and (_27570_, _10244_, _02868_);
  nor (_27571_, _05416_, _10243_);
  nor (_27572_, _27571_, _27570_);
  nor (_27573_, _27572_, _04638_);
  nor (_27574_, _27573_, _27543_);
  nor (_27575_, _27574_, _07474_);
  or (_27576_, _27575_, _27568_);
  and (_27577_, _27576_, _02992_);
  nor (_27578_, _27550_, _02992_);
  or (_27579_, _27578_, _27577_);
  and (_27581_, _27579_, _03962_);
  nor (_27582_, _04220_, _10243_);
  and (_27583_, _04220_, _10243_);
  nor (_27584_, _27583_, _27582_);
  and (_27585_, _27584_, _02876_);
  nor (_27586_, _27585_, _10219_);
  not (_27587_, _27586_);
  nor (_27588_, _27587_, _27581_);
  nor (_27589_, _27555_, _04135_);
  nor (_27590_, _27589_, _05535_);
  not (_27592_, _27590_);
  nor (_27593_, _27592_, _27588_);
  nor (_27594_, _27593_, _27546_);
  and (_27595_, _06171_, _04638_);
  nor (_27596_, _27535_, _02842_);
  not (_27597_, _27596_);
  nor (_27598_, _27597_, _27595_);
  or (_27599_, _27598_, _02567_);
  nor (_27600_, _27599_, _27594_);
  nor (_27601_, _11271_, _10206_);
  nor (_27603_, _27601_, _27535_);
  nor (_27604_, _27603_, _02839_);
  or (_27605_, _27604_, _02834_);
  or (_27606_, _27605_, _27600_);
  and (_27607_, _05618_, _04638_);
  nor (_27608_, _27607_, _27535_);
  nand (_27609_, _27608_, _02834_);
  and (_27610_, _27609_, _27606_);
  nor (_27611_, _27610_, _02522_);
  and (_27612_, _27556_, _02522_);
  nor (_27614_, _27612_, _27611_);
  and (_27615_, _27614_, _07139_);
  and (_27616_, _11158_, _04638_);
  nor (_27617_, _27616_, _27535_);
  nor (_27618_, _27617_, _07139_);
  or (_27619_, _27618_, _27615_);
  and (_27620_, _27619_, _07150_);
  nor (_27621_, _27620_, _27542_);
  nor (_27622_, _27621_, _03022_);
  not (_27623_, _27535_);
  and (_27625_, _27623_, _05239_);
  or (_27626_, _27625_, _03023_);
  nor (_27627_, _27626_, _27608_);
  nor (_27628_, _27627_, _27622_);
  nor (_27629_, _27628_, _09463_);
  and (_27630_, _27555_, _02530_);
  nor (_27631_, _27630_, _03042_);
  or (_27632_, _27550_, _06213_);
  or (_27633_, _27632_, _27625_);
  nand (_27634_, _27633_, _27631_);
  nor (_27636_, _27634_, _27629_);
  nor (_27637_, _11157_, _10206_);
  nor (_27638_, _27637_, _27535_);
  and (_27639_, _27638_, _03042_);
  nor (_27640_, _27639_, _27636_);
  nor (_27641_, _27640_, _03143_);
  nor (_27642_, _11152_, _10206_);
  or (_27643_, _27535_, _07161_);
  nor (_27644_, _27643_, _27642_);
  or (_27645_, _27644_, _03155_);
  nor (_27647_, _27645_, _27641_);
  nor (_27648_, _05415_, _10243_);
  nor (_27649_, _27648_, _10244_);
  nor (_27650_, _27649_, _20557_);
  or (_27651_, _27650_, _02528_);
  nor (_27652_, _27651_, _27647_);
  and (_27653_, _27556_, _02528_);
  nor (_27654_, _27653_, _27652_);
  and (_27655_, _27654_, _02891_);
  nor (_27656_, _27649_, _02891_);
  or (_27658_, _27656_, _27655_);
  and (_27659_, _27658_, _03179_);
  nor (_27660_, _27562_, _03179_);
  or (_27661_, _27660_, _04150_);
  nor (_27662_, _27661_, _27659_);
  nor (_27663_, _27555_, _03936_);
  nor (_27664_, _27663_, _02887_);
  not (_27665_, _27664_);
  nor (_27666_, _27665_, _27662_);
  nor (_27667_, _27666_, _27539_);
  nand (_27669_, _27667_, _34655_);
  or (_27670_, _34655_, \oc8051_golden_model_1.SP [4]);
  and (_27671_, _27670_, _35796_);
  and (_35846_[4], _27671_, _27669_);
  nor (_27672_, _04638_, _10242_);
  and (_27673_, _11541_, _04638_);
  nor (_27674_, _27673_, _27672_);
  nor (_27675_, _27674_, _02888_);
  and (_27676_, _10212_, \oc8051_golden_model_1.SP [0]);
  nor (_27677_, _27582_, \oc8051_golden_model_1.SP [5]);
  nor (_27679_, _27677_, _27676_);
  and (_27680_, _27679_, _02876_);
  nor (_27681_, _03845_, _10242_);
  and (_27682_, _04638_, \oc8051_golden_model_1.ACC [5]);
  nor (_27683_, _27682_, _27672_);
  nor (_27684_, _27683_, _04194_);
  or (_27685_, _27684_, _27681_);
  and (_27686_, _27685_, _02603_);
  nor (_27687_, _10211_, \oc8051_golden_model_1.SP [5]);
  nor (_27688_, _27687_, _10212_);
  not (_27689_, _27688_);
  nor (_27690_, _27689_, _02603_);
  nor (_27691_, _27690_, _27686_);
  nor (_27692_, _27691_, _02948_);
  nor (_27693_, _11380_, _10206_);
  nor (_27694_, _27693_, _27672_);
  nor (_27695_, _27694_, _03006_);
  or (_27696_, _27695_, _27692_);
  and (_27697_, _27696_, _02597_);
  nor (_27698_, _27689_, _02597_);
  or (_27701_, _27698_, _27697_);
  and (_27702_, _27701_, _07474_);
  nor (_27703_, _04894_, _10206_);
  and (_27704_, _10245_, _02868_);
  nor (_27705_, _27570_, _10242_);
  nor (_27706_, _27705_, _27704_);
  nor (_27707_, _27706_, _04638_);
  nor (_27708_, _27707_, _27703_);
  nor (_27709_, _27708_, _07474_);
  or (_27710_, _27709_, _27702_);
  and (_27712_, _27710_, _02992_);
  nor (_27713_, _27683_, _02992_);
  or (_27714_, _27713_, _27712_);
  and (_27715_, _27714_, _03962_);
  or (_27716_, _27715_, _10219_);
  nor (_27717_, _27716_, _27680_);
  nor (_27718_, _27688_, _04135_);
  or (_27719_, _27718_, _27717_);
  and (_27720_, _27719_, _02859_);
  nor (_27721_, _27672_, _02859_);
  not (_27723_, _27721_);
  nor (_27724_, _27723_, _27703_);
  nor (_27725_, _27724_, _27720_);
  nor (_27726_, _27725_, _02841_);
  and (_27727_, _06170_, _04638_);
  nor (_27728_, _27672_, _02842_);
  not (_27729_, _27728_);
  nor (_27730_, _27729_, _27727_);
  nor (_27731_, _27730_, _27726_);
  nor (_27732_, _27731_, _02567_);
  nor (_27734_, _11467_, _10206_);
  nor (_27735_, _27734_, _27672_);
  and (_27736_, _27735_, _02567_);
  nor (_27737_, _27736_, _27732_);
  and (_27738_, _27737_, _07140_);
  and (_27739_, _05671_, _04638_);
  nor (_27740_, _27739_, _27672_);
  nor (_27741_, _27740_, _07140_);
  or (_27742_, _27741_, _27738_);
  and (_27743_, _27742_, _04131_);
  and (_27745_, _27688_, _02522_);
  or (_27746_, _27745_, _27743_);
  and (_27747_, _27746_, _07139_);
  and (_27748_, _11482_, _04638_);
  nor (_27749_, _27748_, _27672_);
  nor (_27750_, _27749_, _07139_);
  or (_27751_, _27750_, _27747_);
  and (_27752_, _27751_, _07150_);
  and (_27753_, _11356_, _04638_);
  nor (_27754_, _27753_, _27672_);
  nor (_27756_, _27754_, _07150_);
  or (_27757_, _27756_, _27752_);
  and (_27758_, _27757_, _03023_);
  nor (_27759_, _27672_, _04945_);
  not (_27760_, _27759_);
  nor (_27761_, _27740_, _03023_);
  and (_27762_, _27761_, _27760_);
  nor (_27763_, _27762_, _27758_);
  nor (_27764_, _27763_, _09463_);
  nor (_27765_, _27683_, _06213_);
  and (_27767_, _27765_, _27760_);
  and (_27768_, _27688_, _02530_);
  nor (_27769_, _27768_, _27767_);
  and (_27770_, _27769_, _03043_);
  not (_27771_, _27770_);
  nor (_27772_, _27771_, _27764_);
  nor (_27773_, _11480_, _10206_);
  nor (_27774_, _27773_, _27672_);
  and (_27775_, _27774_, _03042_);
  nor (_27776_, _27775_, _27772_);
  nor (_27778_, _27776_, _03143_);
  nor (_27779_, _11355_, _10206_);
  or (_27780_, _27672_, _07161_);
  nor (_27781_, _27780_, _27779_);
  or (_27782_, _27781_, _03155_);
  nor (_27783_, _27782_, _27778_);
  nor (_27784_, _10244_, _10242_);
  nor (_27785_, _27784_, _10245_);
  nor (_27786_, _27785_, _20557_);
  or (_27787_, _27786_, _02528_);
  nor (_27789_, _27787_, _27783_);
  and (_27790_, _27689_, _02528_);
  nor (_27791_, _27790_, _27789_);
  and (_27792_, _27791_, _02891_);
  nor (_27793_, _27785_, _02891_);
  or (_27794_, _27793_, _27792_);
  and (_27795_, _27794_, _03179_);
  nor (_27796_, _27694_, _03179_);
  or (_27797_, _27796_, _04150_);
  nor (_27798_, _27797_, _27795_);
  nor (_27800_, _27688_, _03936_);
  nor (_27801_, _27800_, _02887_);
  not (_27802_, _27801_);
  nor (_27803_, _27802_, _27798_);
  nor (_27804_, _27803_, _27675_);
  nand (_27805_, _27804_, _34655_);
  or (_27806_, _34655_, \oc8051_golden_model_1.SP [5]);
  and (_27807_, _27806_, _35796_);
  and (_35846_[5], _27807_, _27805_);
  nor (_27808_, _04790_, _10206_);
  nor (_27810_, _04638_, _10241_);
  nor (_27811_, _27810_, _02859_);
  not (_27812_, _27811_);
  nor (_27813_, _27812_, _27808_);
  nor (_27814_, _03845_, _10241_);
  and (_27815_, _04638_, \oc8051_golden_model_1.ACC [6]);
  nor (_27816_, _27815_, _27810_);
  nor (_27817_, _27816_, _04194_);
  or (_27818_, _27817_, _27814_);
  and (_27819_, _27818_, _02603_);
  nor (_27821_, _10212_, \oc8051_golden_model_1.SP [6]);
  nor (_27822_, _27821_, _10213_);
  not (_27823_, _27822_);
  nor (_27824_, _27823_, _02603_);
  nor (_27825_, _27824_, _27819_);
  nor (_27826_, _27825_, _02948_);
  nor (_27827_, _11567_, _10206_);
  nor (_27828_, _27827_, _27810_);
  nor (_27829_, _27828_, _03006_);
  or (_27830_, _27829_, _27826_);
  and (_27832_, _27830_, _02597_);
  nor (_27833_, _27823_, _02597_);
  or (_27834_, _27833_, _27832_);
  and (_27835_, _27834_, _07474_);
  nor (_27836_, _27704_, _10241_);
  nor (_27837_, _27836_, _10247_);
  nor (_27838_, _27837_, _04638_);
  nor (_27839_, _27838_, _27808_);
  nor (_27840_, _27839_, _07474_);
  or (_27841_, _27840_, _27835_);
  and (_27843_, _27841_, _02992_);
  nor (_27844_, _27816_, _02992_);
  or (_27845_, _27844_, _27843_);
  and (_27846_, _27845_, _03962_);
  nor (_27847_, _27676_, \oc8051_golden_model_1.SP [6]);
  nor (_27848_, _27847_, _10214_);
  and (_27849_, _27848_, _02876_);
  nor (_27850_, _27849_, _27846_);
  nor (_27851_, _27850_, _10219_);
  nor (_27852_, _27823_, _04135_);
  nor (_27854_, _27852_, _05535_);
  not (_27855_, _27854_);
  nor (_27856_, _27855_, _27851_);
  nor (_27857_, _27856_, _27813_);
  nor (_27858_, _27857_, _02841_);
  and (_27859_, _06162_, _04638_);
  nor (_27860_, _27810_, _02842_);
  not (_27861_, _27860_);
  nor (_27862_, _27861_, _27859_);
  nor (_27863_, _27862_, _27858_);
  nor (_27865_, _27863_, _02567_);
  nor (_27866_, _11671_, _10206_);
  nor (_27867_, _27866_, _27810_);
  and (_27868_, _27867_, _02567_);
  nor (_27869_, _27868_, _27865_);
  and (_27870_, _27869_, _07140_);
  and (_27871_, _11678_, _04638_);
  nor (_27872_, _27871_, _27810_);
  nor (_27873_, _27872_, _07140_);
  or (_27874_, _27873_, _27870_);
  and (_27876_, _27874_, _04131_);
  and (_27877_, _27822_, _02522_);
  or (_27878_, _27877_, _27876_);
  and (_27879_, _27878_, _07139_);
  and (_27880_, _11560_, _04638_);
  nor (_27881_, _27880_, _27810_);
  nor (_27882_, _27881_, _07139_);
  or (_27883_, _27882_, _27879_);
  and (_27884_, _27883_, _07150_);
  and (_27885_, _11556_, _04638_);
  nor (_27887_, _27885_, _27810_);
  nor (_27888_, _27887_, _07150_);
  or (_27889_, _27888_, _27884_);
  and (_27890_, _27889_, _03023_);
  nor (_27891_, _27810_, _04838_);
  not (_27892_, _27891_);
  nor (_27893_, _27872_, _03023_);
  and (_27894_, _27893_, _27892_);
  nor (_27895_, _27894_, _27890_);
  nor (_27896_, _27895_, _09463_);
  and (_27898_, _27822_, _02530_);
  or (_27899_, _27891_, _06213_);
  nor (_27900_, _27899_, _27816_);
  or (_27901_, _27900_, _27898_);
  or (_27902_, _27901_, _03042_);
  nor (_27903_, _27902_, _27896_);
  nor (_27904_, _11558_, _10206_);
  nor (_27905_, _27904_, _27810_);
  and (_27906_, _27905_, _03042_);
  nor (_27907_, _27906_, _27903_);
  nor (_27909_, _27907_, _03143_);
  nor (_27910_, _11555_, _10206_);
  or (_27911_, _27810_, _07161_);
  nor (_27912_, _27911_, _27910_);
  or (_27913_, _27912_, _03155_);
  nor (_27914_, _27913_, _27909_);
  nor (_27915_, _10245_, _10241_);
  nor (_27916_, _27915_, _10246_);
  not (_27917_, _27916_);
  and (_27918_, _27917_, _03155_);
  or (_27920_, _27918_, _02528_);
  nor (_27921_, _27920_, _27914_);
  and (_27922_, _27823_, _02528_);
  or (_27923_, _27922_, _02890_);
  nor (_27924_, _27923_, _27921_);
  and (_27925_, _27917_, _02890_);
  or (_27926_, _27925_, _03174_);
  nor (_27927_, _27926_, _27924_);
  and (_27928_, _27828_, _03174_);
  nor (_27929_, _27928_, _04150_);
  not (_27931_, _27929_);
  nor (_27932_, _27931_, _27927_);
  nor (_27933_, _27823_, _03936_);
  nor (_27934_, _27933_, _02887_);
  not (_27935_, _27934_);
  nor (_27936_, _27935_, _27932_);
  and (_27937_, _11744_, _04638_);
  nor (_27938_, _27937_, _27810_);
  and (_27939_, _27938_, _02887_);
  nor (_27940_, _27939_, _27936_);
  or (_27942_, _27940_, _34659_);
  or (_27943_, _34655_, \oc8051_golden_model_1.SP [6]);
  and (_27944_, _27943_, _35796_);
  and (_35846_[6], _27944_, _27942_);
  and (_35847_[0], \oc8051_golden_model_1.TCON [0], _35796_);
  and (_35847_[1], \oc8051_golden_model_1.TCON [1], _35796_);
  and (_35847_[2], \oc8051_golden_model_1.TCON [2], _35796_);
  and (_35847_[3], \oc8051_golden_model_1.TCON [3], _35796_);
  and (_35847_[4], \oc8051_golden_model_1.TCON [4], _35796_);
  and (_35847_[5], \oc8051_golden_model_1.TCON [5], _35796_);
  and (_35847_[6], \oc8051_golden_model_1.TCON [6], _35796_);
  and (_35848_[0], \oc8051_golden_model_1.TH0 [0], _35796_);
  and (_35848_[1], \oc8051_golden_model_1.TH0 [1], _35796_);
  and (_35848_[2], \oc8051_golden_model_1.TH0 [2], _35796_);
  and (_35848_[3], \oc8051_golden_model_1.TH0 [3], _35796_);
  and (_35848_[4], \oc8051_golden_model_1.TH0 [4], _35796_);
  and (_35848_[5], \oc8051_golden_model_1.TH0 [5], _35796_);
  and (_35848_[6], \oc8051_golden_model_1.TH0 [6], _35796_);
  and (_35849_[0], \oc8051_golden_model_1.TH1 [0], _35796_);
  and (_35849_[1], \oc8051_golden_model_1.TH1 [1], _35796_);
  and (_35849_[2], \oc8051_golden_model_1.TH1 [2], _35796_);
  and (_35849_[3], \oc8051_golden_model_1.TH1 [3], _35796_);
  and (_35849_[4], \oc8051_golden_model_1.TH1 [4], _35796_);
  and (_35849_[5], \oc8051_golden_model_1.TH1 [5], _35796_);
  and (_35849_[6], \oc8051_golden_model_1.TH1 [6], _35796_);
  and (_35850_[0], \oc8051_golden_model_1.TL0 [0], _35796_);
  and (_35850_[1], \oc8051_golden_model_1.TL0 [1], _35796_);
  and (_35850_[2], \oc8051_golden_model_1.TL0 [2], _35796_);
  and (_35850_[3], \oc8051_golden_model_1.TL0 [3], _35796_);
  and (_35850_[4], \oc8051_golden_model_1.TL0 [4], _35796_);
  and (_35850_[5], \oc8051_golden_model_1.TL0 [5], _35796_);
  and (_35850_[6], \oc8051_golden_model_1.TL0 [6], _35796_);
  and (_35851_[0], \oc8051_golden_model_1.TL1 [0], _35796_);
  and (_35851_[1], \oc8051_golden_model_1.TL1 [1], _35796_);
  and (_35851_[2], \oc8051_golden_model_1.TL1 [2], _35796_);
  and (_35851_[3], \oc8051_golden_model_1.TL1 [3], _35796_);
  and (_35851_[4], \oc8051_golden_model_1.TL1 [4], _35796_);
  and (_35851_[5], \oc8051_golden_model_1.TL1 [5], _35796_);
  and (_35851_[6], \oc8051_golden_model_1.TL1 [6], _35796_);
  and (_35852_[0], \oc8051_golden_model_1.TMOD [0], _35796_);
  and (_35852_[1], \oc8051_golden_model_1.TMOD [1], _35796_);
  and (_35852_[2], \oc8051_golden_model_1.TMOD [2], _35796_);
  and (_35852_[3], \oc8051_golden_model_1.TMOD [3], _35796_);
  and (_35852_[4], \oc8051_golden_model_1.TMOD [4], _35796_);
  and (_35852_[5], \oc8051_golden_model_1.TMOD [5], _35796_);
  and (_35852_[6], \oc8051_golden_model_1.TMOD [6], _35796_);
  and (_27949_, _21260_, _07965_);
  and (_27950_, _03144_, _02534_);
  and (_27951_, _21747_, _08812_);
  and (_27952_, _27951_, _27950_);
  and (_27954_, _27952_, _27949_);
  not (_27955_, _03591_);
  not (_27956_, _07187_);
  not (_27957_, _03570_);
  and (_27958_, _03002_, _02509_);
  nor (_27959_, _03728_, _27958_);
  and (_27960_, _27959_, _27957_);
  and (_27961_, _27960_, _27956_);
  not (_27962_, _24720_);
  nor (_27963_, _03276_, _03358_);
  and (_27965_, _27963_, _27962_);
  and (_27966_, _27965_, _27961_);
  nor (_27967_, _23075_, _09719_);
  and (_27968_, _27967_, _27966_);
  and (_27969_, _27968_, _20609_);
  and (_27970_, _27969_, _27955_);
  and (_27971_, _27970_, _27954_);
  and (_27972_, _09345_, _09336_);
  and (_27973_, _03138_, _19615_);
  and (_27974_, _09437_, _07139_);
  and (_27976_, _21214_, _09455_);
  and (_27977_, _27976_, _27974_);
  and (_27978_, _27977_, _27973_);
  and (_27979_, _27978_, _27972_);
  and (_27980_, _09186_, _07474_);
  and (_27981_, _08993_, _03006_);
  and (_27982_, _27981_, _08997_);
  and (_27983_, _27982_, _27980_);
  and (_27984_, _09134_, \oc8051_golden_model_1.ACC [0]);
  nor (_27985_, _02798_, _02370_);
  and (_27987_, _27985_, _03382_);
  not (_27988_, _27987_);
  and (_27989_, _27988_, \oc8051_golden_model_1.XRAM_DATA_OUT [0]);
  nor (_27990_, _27989_, _27984_);
  nor (_27991_, _09150_, _03849_);
  not (_27992_, _27991_);
  nor (_27993_, _27992_, _27990_);
  and (_27994_, _09150_, \oc8051_golden_model_1.ACC [0]);
  nor (_27995_, _27994_, _27993_);
  not (_27996_, _27995_);
  and (_27998_, _09195_, _08990_);
  and (_27999_, _25005_, _03962_);
  and (_28000_, _27999_, _27998_);
  not (_28001_, _04029_);
  and (_28002_, _05360_, _28001_);
  and (_28003_, _09133_, _28002_);
  and (_28004_, _28003_, _28000_);
  and (_28005_, _28004_, _27996_);
  and (_28006_, _28005_, _27983_);
  and (_28007_, _09366_, _05748_);
  and (_28009_, _09360_, _09353_);
  and (_28010_, _28009_, _28007_);
  and (_28011_, _28010_, _07140_);
  nor (_28012_, _02967_, _02960_);
  nor (_28013_, _08786_, _02957_);
  and (_28014_, _28013_, _28012_);
  nor (_28015_, _03927_, _03587_);
  and (_28016_, _28015_, _02601_);
  and (_28017_, _28016_, _24424_);
  and (_28018_, _28017_, _28014_);
  and (_28020_, _07421_, _07411_);
  and (_28021_, _09260_, _09258_);
  nor (_28022_, _03840_, _04028_);
  and (_28023_, _28022_, _09251_);
  and (_28024_, _28023_, _28021_);
  and (_28025_, _28024_, _28020_);
  and (_28026_, _09732_, _27274_);
  and (_28027_, _19862_, _20617_);
  and (_28028_, _28027_, _28026_);
  not (_28029_, _02963_);
  nor (_28031_, _25074_, _03889_);
  and (_28032_, _28031_, _28029_);
  and (_28033_, _28032_, _09308_);
  and (_28034_, _02864_, _02565_);
  nor (_28035_, _28034_, _03448_);
  and (_28036_, _28035_, _10027_);
  and (_28037_, _28036_, _22802_);
  and (_28038_, _28037_, _28033_);
  and (_28039_, _28038_, _28028_);
  and (_28040_, _28039_, _28025_);
  and (_28042_, _28040_, _28018_);
  and (_28043_, _25964_, _03270_);
  and (_28044_, _05797_, _09718_);
  and (_28045_, _28044_, _28043_);
  and (_28046_, _25384_, _07831_);
  and (_28047_, _28046_, _08822_);
  and (_28048_, _28047_, _08823_);
  and (_28049_, _28048_, _28045_);
  and (_28050_, _28049_, _28042_);
  and (_28051_, _28050_, _28011_);
  and (_28053_, _28051_, _28006_);
  and (_28054_, _28053_, _27979_);
  and (_28055_, _28054_, _27971_);
  or (_28056_, _28055_, _34659_);
  or (_28057_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [0]);
  and (_28058_, _28057_, _35796_);
  and (_35854_[0], _28058_, _28056_);
  and (_28059_, _28020_, _24424_);
  and (_28060_, _28059_, _02601_);
  and (_28061_, _28060_, _27972_);
  and (_28063_, _11570_, _09133_);
  and (_28064_, _28063_, _27983_);
  and (_28065_, _09134_, \oc8051_golden_model_1.ACC [1]);
  and (_28066_, _27988_, \oc8051_golden_model_1.XRAM_DATA_OUT [1]);
  nor (_28067_, _28066_, _28065_);
  nor (_28068_, _28067_, _27992_);
  and (_28069_, _09150_, \oc8051_golden_model_1.ACC [1]);
  nor (_28070_, _28069_, _28068_);
  not (_28071_, _28070_);
  and (_28072_, _09324_, _08787_);
  and (_28074_, _28072_, _28015_);
  and (_28075_, _28074_, _28028_);
  and (_28076_, _28075_, _28045_);
  and (_28077_, _28076_, _28071_);
  and (_28078_, _28077_, _28064_);
  and (_28079_, _28078_, _28061_);
  and (_28080_, _28079_, _27971_);
  and (_28081_, _09316_, _09309_);
  and (_28082_, _28081_, _09263_);
  and (_28083_, _27999_, _09251_);
  and (_28084_, _28083_, _28082_);
  and (_28085_, _28084_, _09320_);
  and (_28086_, _28085_, _27998_);
  and (_28087_, _28048_, _07140_);
  and (_28088_, _28087_, _27978_);
  and (_28089_, _28088_, _28010_);
  and (_28090_, _28089_, _28086_);
  and (_28091_, _28090_, _28080_);
  or (_28092_, _28091_, _34659_);
  or (_28093_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [1]);
  and (_28096_, _28093_, _35796_);
  and (_35854_[1], _28096_, _28092_);
  and (_28097_, _28072_, _27955_);
  and (_28098_, _28097_, _28026_);
  and (_28099_, _28098_, _27969_);
  and (_28100_, _09134_, \oc8051_golden_model_1.ACC [2]);
  and (_28101_, _27988_, \oc8051_golden_model_1.XRAM_DATA_OUT [2]);
  nor (_28102_, _28101_, _28100_);
  nor (_28103_, _28102_, _27992_);
  and (_28104_, _09150_, \oc8051_golden_model_1.ACC [2]);
  nor (_28106_, _28104_, _28103_);
  and (_28107_, _04105_, _05809_);
  and (_28108_, _04130_, _09718_);
  and (_28109_, _28108_, _28107_);
  and (_28110_, _28109_, _28043_);
  and (_28111_, _28027_, _27998_);
  and (_28112_, _28111_, _28110_);
  not (_28113_, _28112_);
  nor (_28114_, _28113_, _28106_);
  and (_28115_, _28114_, _28087_);
  and (_28117_, _28115_, _28099_);
  and (_28118_, _28117_, _28085_);
  and (_28119_, _28064_, _27978_);
  and (_28120_, _28119_, _28010_);
  and (_28121_, _28061_, _27954_);
  and (_28122_, _28121_, _28120_);
  and (_28123_, _28122_, _28118_);
  or (_28124_, _28123_, _34659_);
  or (_28125_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [2]);
  and (_28126_, _28125_, _35796_);
  and (_35854_[2], _28126_, _28124_);
  or (_28128_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [3]);
  and (_28129_, _28128_, _35796_);
  and (_28130_, _09134_, \oc8051_golden_model_1.ACC [3]);
  and (_28131_, _27988_, \oc8051_golden_model_1.XRAM_DATA_OUT [3]);
  nor (_28132_, _28131_, _28130_);
  nor (_28133_, _28132_, _27992_);
  and (_28134_, _09150_, \oc8051_golden_model_1.ACC [3]);
  nor (_28135_, _28134_, _28133_);
  not (_28136_, _28135_);
  and (_28138_, _28112_, _28087_);
  and (_28139_, _28138_, _28136_);
  and (_28140_, _28098_, _09320_);
  and (_28141_, _28140_, _27969_);
  and (_28142_, _28141_, _28084_);
  and (_28143_, _28142_, _28139_);
  and (_28144_, _28143_, _28121_);
  and (_28145_, _28144_, _28120_);
  or (_28146_, _28145_, _34659_);
  and (_35854_[3], _28146_, _28129_);
  and (_28148_, _27970_, _28026_);
  and (_28149_, _28148_, _28110_);
  and (_28150_, _28048_, _09345_);
  and (_28151_, _28009_, _09336_);
  and (_28152_, _28151_, _28072_);
  and (_28153_, _28152_, _28027_);
  and (_28154_, _28153_, _28060_);
  and (_28155_, _28154_, _28150_);
  and (_28156_, _28155_, _07140_);
  and (_28157_, _28156_, _28149_);
  and (_28159_, _09134_, \oc8051_golden_model_1.ACC [4]);
  and (_28160_, _27988_, \oc8051_golden_model_1.XRAM_DATA_OUT [4]);
  nor (_28161_, _28160_, _28159_);
  nor (_28162_, _28161_, _27992_);
  and (_28163_, _09150_, \oc8051_golden_model_1.ACC [4]);
  nor (_28164_, _28163_, _28162_);
  nand (_28165_, _28064_, _28007_);
  nor (_28166_, _28165_, _28164_);
  and (_28167_, _28166_, _28157_);
  and (_28168_, _27954_, _27978_);
  and (_28170_, _28168_, _28086_);
  and (_28171_, _28170_, _28167_);
  or (_28172_, _28171_, _34659_);
  or (_28173_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [4]);
  and (_28174_, _28173_, _35796_);
  and (_35854_[4], _28174_, _28172_);
  and (_28175_, _27983_, _02600_);
  and (_28176_, _09134_, \oc8051_golden_model_1.ACC [5]);
  and (_28177_, _27988_, \oc8051_golden_model_1.XRAM_DATA_OUT [5]);
  nor (_28178_, _28177_, _28176_);
  nor (_28180_, _28178_, _27992_);
  and (_28181_, _09150_, \oc8051_golden_model_1.ACC [5]);
  nor (_28182_, _28181_, _28180_);
  not (_28183_, _28182_);
  and (_28184_, _28083_, _28021_);
  and (_28185_, _28184_, _28183_);
  and (_28186_, _28185_, _28175_);
  and (_28187_, _27950_, _09336_);
  and (_28188_, _28187_, _11570_);
  and (_28189_, _28188_, _28014_);
  and (_28191_, _28111_, _28038_);
  and (_28192_, _28191_, _28189_);
  and (_28193_, _28192_, _27949_);
  and (_28194_, _27951_, _09345_);
  and (_28195_, _28194_, _28193_);
  and (_28196_, _28195_, _28186_);
  and (_28197_, _28196_, _28089_);
  and (_28198_, _28197_, _28149_);
  or (_28199_, _28198_, _34659_);
  or (_28200_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [5]);
  and (_28202_, _28200_, _35796_);
  and (_35854_[5], _28202_, _28199_);
  and (_28203_, _28027_, _08787_);
  and (_28204_, _20609_, _28026_);
  and (_28205_, _28204_, _28015_);
  and (_28206_, _28205_, _28203_);
  and (_28207_, _09134_, \oc8051_golden_model_1.ACC [6]);
  and (_28208_, _27988_, \oc8051_golden_model_1.XRAM_DATA_OUT [6]);
  nor (_28209_, _28208_, _28207_);
  nor (_28210_, _28209_, _27992_);
  and (_28212_, _09150_, \oc8051_golden_model_1.ACC [6]);
  nor (_28213_, _28212_, _28210_);
  not (_28214_, _28213_);
  and (_28215_, _23074_, _11503_);
  and (_28216_, _28215_, _27966_);
  and (_28217_, _28036_, _28081_);
  and (_28218_, _28063_, _09259_);
  and (_28219_, _28218_, _28217_);
  and (_28220_, _28219_, _28216_);
  and (_28221_, _28220_, _28214_);
  and (_28223_, _28221_, _27952_);
  and (_28224_, _28223_, _28061_);
  and (_28225_, _28224_, _28206_);
  and (_28226_, _28043_, _27949_);
  and (_28227_, _28184_, _27998_);
  and (_28228_, _27983_, _04063_);
  and (_28229_, _28228_, _28227_);
  and (_28230_, _28229_, _28226_);
  and (_28231_, _28230_, _28089_);
  and (_28232_, _28231_, _28225_);
  or (_28234_, _28232_, _34659_);
  or (_28235_, _34655_, \oc8051_golden_model_1.XRAM_DATA_OUT [6]);
  and (_28236_, _28235_, _35796_);
  and (_35854_[6], _28236_, _28234_);
  and (_28237_, _07433_, \oc8051_golden_model_1.DPL [0]);
  nor (_28238_, _07433_, _09169_);
  not (_28239_, _28238_);
  nor (_28240_, _09134_, _07440_);
  or (_28241_, _28240_, _03872_);
  and (_28242_, _09150_, \oc8051_golden_model_1.DPL [0]);
  nand (_28244_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [0]);
  nor (_28245_, _28244_, _27987_);
  or (_28246_, _28245_, _28242_);
  nand (_28247_, _28246_, _28059_);
  and (_28248_, _28247_, _28241_);
  nor (_28249_, _28248_, _28239_);
  nor (_28250_, _28249_, _28237_);
  and (_28251_, _28228_, _11570_);
  and (_28252_, _28251_, _28227_);
  and (_28253_, _28252_, _09259_);
  and (_28255_, _28217_, _27972_);
  and (_28256_, _28255_, _28011_);
  and (_28257_, _28256_, _28253_);
  and (_28258_, _28048_, _27978_);
  and (_28259_, _28226_, _27952_);
  and (_28260_, _28259_, _28258_);
  and (_28261_, _28260_, _28257_);
  and (_28262_, _28216_, _28206_);
  and (_28263_, _28262_, _28261_);
  not (_28264_, _28263_);
  nor (_28265_, _28264_, _28250_);
  or (_28266_, _28265_, _34659_);
  or (_28267_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [0]);
  and (_28268_, _28267_, _35796_);
  and (_35853_[0], _28268_, _28266_);
  and (_28269_, _07433_, \oc8051_golden_model_1.DPL [1]);
  or (_28270_, _28240_, _04020_);
  and (_28271_, _09150_, \oc8051_golden_model_1.DPL [1]);
  nand (_28272_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [1]);
  nor (_28273_, _28272_, _27987_);
  or (_28276_, _28273_, _28271_);
  nand (_28277_, _28276_, _28059_);
  and (_28278_, _28277_, _28270_);
  nor (_28279_, _28278_, _28239_);
  nor (_28280_, _28279_, _28269_);
  nor (_28281_, _28280_, _28264_);
  or (_28282_, _28281_, _34659_);
  or (_28283_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [1]);
  and (_28284_, _28283_, _35796_);
  and (_35853_[1], _28284_, _28282_);
  and (_28286_, _07433_, \oc8051_golden_model_1.DPL [2]);
  or (_28287_, _28240_, _04449_);
  and (_28288_, _09150_, \oc8051_golden_model_1.DPL [2]);
  nand (_28289_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [2]);
  nor (_28290_, _28289_, _27987_);
  or (_28291_, _28290_, _28288_);
  nand (_28292_, _28291_, _28059_);
  and (_28293_, _28292_, _28287_);
  nor (_28294_, _28293_, _28239_);
  nor (_28295_, _28294_, _28286_);
  nor (_28297_, _28295_, _28264_);
  or (_28298_, _28297_, _34659_);
  or (_28299_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [2]);
  and (_28300_, _28299_, _35796_);
  and (_35853_[2], _28300_, _28298_);
  and (_28301_, _07433_, \oc8051_golden_model_1.DPL [3]);
  or (_28302_, _28240_, _04275_);
  and (_28303_, _09150_, \oc8051_golden_model_1.DPL [3]);
  nand (_28304_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [3]);
  nor (_28305_, _28304_, _27987_);
  or (_28307_, _28305_, _28303_);
  nand (_28308_, _28307_, _28059_);
  and (_28309_, _28308_, _28302_);
  nor (_28310_, _28309_, _28239_);
  nor (_28311_, _28310_, _28301_);
  nor (_28312_, _28311_, _28264_);
  or (_28313_, _28312_, _34659_);
  or (_28314_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [3]);
  and (_28315_, _28314_, _35796_);
  and (_35853_[3], _28315_, _28313_);
  and (_28317_, _07433_, \oc8051_golden_model_1.DPL [4]);
  or (_28318_, _28240_, _05192_);
  and (_28319_, _09150_, \oc8051_golden_model_1.DPL [4]);
  nand (_28320_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [4]);
  nor (_28321_, _28320_, _27987_);
  or (_28322_, _28321_, _28319_);
  nand (_28323_, _28322_, _28059_);
  and (_28324_, _28323_, _28318_);
  nor (_28325_, _28324_, _28239_);
  nor (_28326_, _28325_, _28317_);
  nor (_28328_, _28326_, _28264_);
  or (_28329_, _28328_, _34659_);
  or (_28330_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [4]);
  and (_28331_, _28330_, _35796_);
  and (_35853_[4], _28331_, _28329_);
  and (_28332_, _07433_, \oc8051_golden_model_1.DPL [5]);
  or (_28333_, _28240_, _04894_);
  and (_28334_, _09150_, \oc8051_golden_model_1.DPL [5]);
  nand (_28335_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [5]);
  nor (_28336_, _28335_, _27987_);
  or (_28338_, _28336_, _28334_);
  nand (_28339_, _28338_, _28059_);
  and (_28340_, _28339_, _28333_);
  nor (_28341_, _28340_, _28239_);
  nor (_28342_, _28341_, _28332_);
  nor (_28343_, _28342_, _28264_);
  or (_28344_, _28343_, _34659_);
  or (_28345_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [5]);
  and (_28346_, _28345_, _35796_);
  and (_35853_[5], _28346_, _28344_);
  and (_28348_, _07433_, \oc8051_golden_model_1.DPL [6]);
  or (_28349_, _28240_, _04790_);
  and (_28350_, _09150_, \oc8051_golden_model_1.DPL [6]);
  nand (_28351_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [6]);
  nor (_28352_, _28351_, _27987_);
  or (_28353_, _28352_, _28350_);
  nand (_28354_, _28353_, _28059_);
  and (_28355_, _28354_, _28349_);
  nor (_28356_, _28355_, _28239_);
  nor (_28357_, _28356_, _28348_);
  nor (_28359_, _28357_, _28264_);
  or (_28360_, _28359_, _34659_);
  or (_28361_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [6]);
  and (_28362_, _28361_, _35796_);
  and (_35853_[6], _28362_, _28360_);
  and (_28363_, _07433_, \oc8051_golden_model_1.DPL [7]);
  or (_28364_, _28240_, _04630_);
  and (_28365_, _09150_, \oc8051_golden_model_1.DPL [7]);
  nand (_28366_, _27991_, \oc8051_golden_model_1.XRAM_ADDR [7]);
  nor (_28367_, _28366_, _27987_);
  or (_28369_, _28367_, _28365_);
  nand (_28370_, _28369_, _28059_);
  and (_28371_, _28370_, _28364_);
  nor (_28372_, _28371_, _28239_);
  nor (_28373_, _28372_, _28363_);
  nor (_28374_, _28373_, _28264_);
  or (_28375_, _28374_, _34659_);
  or (_28376_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [7]);
  and (_28377_, _28376_, _35796_);
  and (_35853_[7], _28377_, _28375_);
  or (_28379_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [8]);
  and (_28380_, _28379_, _35796_);
  nor (_28381_, _10345_, _09380_);
  or (_28382_, _28381_, _34659_);
  and (_35853_[8], _28382_, _28380_);
  and (_28383_, _27962_, _07188_);
  and (_28384_, _28383_, _21293_);
  and (_28385_, _28384_, _28215_);
  and (_28386_, _28385_, _27952_);
  and (_28387_, _28386_, _28088_);
  and (_28389_, _28387_, _28253_);
  and (_28390_, _02602_, \oc8051_golden_model_1.XRAM_ADDR [9]);
  and (_28391_, _09150_, \oc8051_golden_model_1.DPH [1]);
  nor (_28392_, _28391_, _28390_);
  nor (_28393_, _28392_, _02949_);
  and (_28394_, _07433_, \oc8051_golden_model_1.DPH [1]);
  nor (_28395_, _28394_, _28393_);
  not (_28396_, _28395_);
  and (_28397_, _28010_, _27972_);
  and (_28398_, _25964_, _07186_);
  and (_28400_, _28398_, _27949_);
  and (_28401_, _28217_, _28206_);
  and (_28402_, _28401_, _28400_);
  and (_28403_, _28402_, _28397_);
  and (_28404_, _28403_, _28396_);
  and (_28405_, _28404_, _28389_);
  or (_28406_, _28405_, _34659_);
  or (_28407_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [9]);
  and (_28408_, _28407_, _35796_);
  and (_35853_[9], _28408_, _28406_);
  or (_28409_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [10]);
  and (_28410_, _28409_, _35796_);
  and (_28411_, _27972_, _27977_);
  and (_28412_, _28036_, _10030_);
  and (_28413_, _28412_, _28033_);
  nor (_28414_, _02960_, _19627_);
  and (_28415_, _28414_, _02958_);
  and (_28416_, _28415_, _28413_);
  and (_28417_, _28416_, _28385_);
  and (_28418_, _28417_, _28010_);
  and (_28420_, _28418_, _28087_);
  and (_28421_, _28420_, _28411_);
  and (_28422_, _02602_, \oc8051_golden_model_1.XRAM_ADDR [10]);
  and (_28423_, _09150_, \oc8051_golden_model_1.DPH [2]);
  nor (_28424_, _28423_, _28422_);
  nor (_28425_, _28424_, _02949_);
  and (_28426_, _07433_, \oc8051_golden_model_1.DPH [2]);
  nor (_28427_, _28426_, _28425_);
  not (_28428_, _28427_);
  and (_28429_, _28428_, _28206_);
  and (_28431_, _28429_, _28421_);
  and (_28432_, _27952_, _27973_);
  and (_28433_, _28432_, _28400_);
  and (_28434_, _28433_, _28252_);
  and (_28435_, _28434_, _28431_);
  or (_28436_, _28435_, _34659_);
  and (_35853_[10], _28436_, _28410_);
  or (_28437_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [11]);
  and (_28438_, _28437_, _35796_);
  and (_28439_, _28398_, _28203_);
  and (_28441_, _28439_, _28217_);
  and (_28442_, _28441_, _28397_);
  and (_28443_, _02602_, \oc8051_golden_model_1.XRAM_ADDR [11]);
  and (_28444_, _09150_, \oc8051_golden_model_1.DPH [3]);
  nor (_28445_, _28444_, _28443_);
  nor (_28446_, _28445_, _02949_);
  and (_28447_, _07433_, \oc8051_golden_model_1.DPH [3]);
  nor (_28448_, _28447_, _28446_);
  not (_28449_, _28448_);
  and (_28450_, _28205_, _27949_);
  and (_28452_, _28450_, _28449_);
  and (_28453_, _28452_, _28442_);
  and (_28454_, _28453_, _28389_);
  or (_28455_, _28454_, _34659_);
  and (_35853_[11], _28455_, _28438_);
  or (_28456_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [12]);
  and (_28457_, _28456_, _35796_);
  and (_28458_, _28397_, _28252_);
  and (_28459_, _02602_, \oc8051_golden_model_1.XRAM_ADDR [12]);
  and (_28460_, _09150_, \oc8051_golden_model_1.DPH [4]);
  nor (_28462_, _28460_, _28459_);
  nor (_28463_, _28462_, _02949_);
  and (_28464_, _07433_, \oc8051_golden_model_1.DPH [4]);
  nor (_28465_, _28464_, _28463_);
  not (_28466_, _28465_);
  and (_28467_, _28046_, _13645_);
  and (_28468_, _28467_, _28385_);
  and (_28469_, _08822_, _07850_);
  and (_28470_, _28469_, _13654_);
  nor (_28471_, _08786_, _02834_);
  and (_28473_, _28471_, _02958_);
  and (_28474_, _28473_, _28414_);
  and (_28475_, _28474_, _28027_);
  and (_28476_, _28475_, _28470_);
  and (_28477_, _28476_, _28413_);
  and (_28478_, _28477_, _27977_);
  and (_28479_, _28478_, _28468_);
  and (_28480_, _28479_, _28205_);
  and (_28481_, _28480_, _28466_);
  and (_28482_, _28481_, _28433_);
  and (_28484_, _28482_, _28458_);
  or (_28485_, _28484_, _34659_);
  and (_35853_[12], _28485_, _28457_);
  or (_28486_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [13]);
  and (_28487_, _28486_, _35796_);
  and (_28488_, _02602_, \oc8051_golden_model_1.XRAM_ADDR [13]);
  and (_28489_, _09150_, \oc8051_golden_model_1.DPH [5]);
  nor (_28490_, _28489_, _28488_);
  nor (_28491_, _28490_, _02949_);
  and (_28492_, _07433_, \oc8051_golden_model_1.DPH [5]);
  nor (_28494_, _28492_, _28491_);
  nor (_28495_, _28494_, _28264_);
  or (_28496_, _28495_, _34659_);
  and (_35853_[13], _28496_, _28487_);
  or (_28497_, _34655_, \oc8051_golden_model_1.XRAM_ADDR [14]);
  and (_28498_, _28497_, _35796_);
  and (_28499_, _27976_, _27973_);
  and (_28500_, _03298_, _02864_);
  not (_28501_, _28500_);
  and (_28502_, _22802_, _28501_);
  and (_28504_, _28502_, _02958_);
  and (_28505_, _28035_, _28033_);
  nor (_28506_, _03767_, _03456_);
  and (_28507_, _09437_, _08822_);
  nor (_28508_, _02960_, _02834_);
  and (_28509_, _28508_, _28507_);
  and (_28510_, _28509_, _28506_);
  and (_28511_, _28510_, _28505_);
  and (_28512_, _28511_, _28504_);
  and (_28513_, _28512_, _28046_);
  and (_28515_, _28513_, _28499_);
  and (_28516_, _28515_, _19619_);
  and (_28517_, _28516_, _28400_);
  and (_28518_, _28517_, _28206_);
  and (_28519_, _02602_, \oc8051_golden_model_1.XRAM_ADDR [14]);
  and (_28520_, _09150_, \oc8051_golden_model_1.DPH [6]);
  nor (_28521_, _28520_, _28519_);
  nor (_28522_, _28521_, _02949_);
  and (_28523_, _07433_, \oc8051_golden_model_1.DPH [6]);
  nor (_28524_, _28523_, _28522_);
  not (_28526_, _28524_);
  and (_28527_, _28526_, _28386_);
  and (_28528_, _28527_, _28518_);
  and (_28529_, _28528_, _28458_);
  or (_28530_, _28529_, _34659_);
  and (_35853_[14], _28530_, _28498_);
  and (_28531_, _34659_, \oc8051_golden_model_1.P0INREG [0]);
  or (_28532_, _28531_, _00500_);
  and (_35833_[0], _28532_, _35796_);
  and (_28533_, _34659_, \oc8051_golden_model_1.P0INREG [1]);
  or (_28535_, _28533_, _00532_);
  and (_35833_[1], _28535_, _35796_);
  and (_28536_, _34659_, \oc8051_golden_model_1.P0INREG [2]);
  or (_28537_, _28536_, _00516_);
  and (_35833_[2], _28537_, _35796_);
  and (_28538_, _34659_, \oc8051_golden_model_1.P0INREG [3]);
  or (_28539_, _28538_, _00485_);
  and (_35833_[3], _28539_, _35796_);
  and (_28540_, _34659_, \oc8051_golden_model_1.P0INREG [4]);
  or (_28541_, _28540_, _00493_);
  and (_35833_[4], _28541_, _35796_);
  and (_28543_, _34659_, \oc8051_golden_model_1.P0INREG [5]);
  or (_28544_, _28543_, _00525_);
  and (_35833_[5], _28544_, _35796_);
  and (_28545_, _34659_, \oc8051_golden_model_1.P0INREG [6]);
  or (_28546_, _28545_, _00509_);
  and (_35833_[6], _28546_, _35796_);
  and (_28547_, _34659_, \oc8051_golden_model_1.P1INREG [0]);
  or (_28548_, _28547_, _00568_);
  and (_35835_[0], _28548_, _35796_);
  and (_28550_, _34659_, \oc8051_golden_model_1.P1INREG [1]);
  or (_28551_, _28550_, _00601_);
  and (_35835_[1], _28551_, _35796_);
  and (_28552_, _34659_, \oc8051_golden_model_1.P1INREG [2]);
  or (_28553_, _28552_, _00584_);
  and (_35835_[2], _28553_, _35796_);
  and (_28554_, _34659_, \oc8051_golden_model_1.P1INREG [3]);
  or (_28555_, _28554_, _00546_);
  and (_35835_[3], _28555_, _35796_);
  and (_28556_, _34659_, \oc8051_golden_model_1.P1INREG [4]);
  or (_28558_, _28556_, _00561_);
  and (_35835_[4], _28558_, _35796_);
  and (_28559_, _34659_, \oc8051_golden_model_1.P1INREG [5]);
  or (_28560_, _28559_, _00594_);
  and (_35835_[5], _28560_, _35796_);
  and (_28561_, _34659_, \oc8051_golden_model_1.P1INREG [6]);
  or (_28562_, _28561_, _00577_);
  and (_35835_[6], _28562_, _35796_);
  and (_28563_, _34659_, \oc8051_golden_model_1.P2INREG [0]);
  or (_28564_, _28563_, _00697_);
  and (_35837_[0], _28564_, _35796_);
  and (_28566_, _34659_, \oc8051_golden_model_1.P2INREG [1]);
  or (_28567_, _28566_, _00738_);
  and (_35837_[1], _28567_, _35796_);
  and (_28568_, _34659_, \oc8051_golden_model_1.P2INREG [2]);
  or (_28569_, _28568_, _00722_);
  and (_35837_[2], _28569_, _35796_);
  and (_28570_, _34659_, \oc8051_golden_model_1.P2INREG [3]);
  or (_28571_, _28570_, _00706_);
  and (_35837_[3], _28571_, _35796_);
  and (_28573_, _34659_, \oc8051_golden_model_1.P2INREG [4]);
  or (_28574_, _28573_, _00690_);
  and (_35837_[4], _28574_, _35796_);
  and (_28575_, _34659_, \oc8051_golden_model_1.P2INREG [5]);
  or (_28576_, _28575_, _00731_);
  and (_35837_[5], _28576_, _35796_);
  and (_28577_, _34659_, \oc8051_golden_model_1.P2INREG [6]);
  or (_28578_, _28577_, _00715_);
  and (_35837_[6], _28578_, _35796_);
  and (_28579_, _34659_, \oc8051_golden_model_1.P3INREG [0]);
  or (_28581_, _28579_, _00630_);
  and (_35839_[0], _28581_, _35796_);
  and (_28582_, _34659_, \oc8051_golden_model_1.P3INREG [1]);
  or (_28583_, _28582_, _00671_);
  and (_35839_[1], _28583_, _35796_);
  and (_28584_, _34659_, \oc8051_golden_model_1.P3INREG [2]);
  or (_28585_, _28584_, _00655_);
  and (_35839_[2], _28585_, _35796_);
  and (_28586_, _34659_, \oc8051_golden_model_1.P3INREG [3]);
  or (_28587_, _28586_, _00639_);
  and (_35839_[3], _28587_, _35796_);
  and (_28589_, _34659_, \oc8051_golden_model_1.P3INREG [4]);
  or (_28590_, _28589_, _00623_);
  and (_35839_[4], _28590_, _35796_);
  and (_28591_, _34659_, \oc8051_golden_model_1.P3INREG [5]);
  or (_28592_, _28591_, _00664_);
  and (_35839_[5], _28592_, _35796_);
  and (_28593_, _34659_, \oc8051_golden_model_1.P3INREG [6]);
  or (_28594_, _28593_, _00648_);
  and (_35839_[6], _28594_, _35796_);
  and (_00005_[6], _00649_, _35796_);
  and (_00005_[5], _00665_, _35796_);
  and (_00005_[4], _00624_, _35796_);
  and (_00005_[3], _00640_, _35796_);
  and (_00005_[2], _00656_, _35796_);
  and (_00005_[1], _00672_, _35796_);
  and (_00005_[0], _00631_, _35796_);
  and (_00004_[6], _00716_, _35796_);
  and (_00004_[5], _00732_, _35796_);
  and (_00004_[4], _00691_, _35796_);
  and (_00004_[3], _00707_, _35796_);
  and (_00004_[2], _00723_, _35796_);
  and (_00004_[1], _00739_, _35796_);
  and (_00004_[0], _00698_, _35796_);
  and (_00003_[6], _00578_, _35796_);
  and (_00003_[5], _00595_, _35796_);
  and (_00003_[4], _00562_, _35796_);
  and (_00003_[3], _00547_, _35796_);
  and (_00003_[2], _00585_, _35796_);
  and (_00003_[1], _00602_, _35796_);
  and (_00003_[0], _00569_, _35796_);
  and (_00002_[6], _00510_, _35796_);
  and (_00002_[5], _00526_, _35796_);
  and (_00002_[4], _00494_, _35796_);
  and (_00002_[3], _00486_, _35796_);
  and (_00002_[2], _00517_, _35796_);
  and (_00002_[1], _00533_, _35796_);
  and (_00002_[0], _00501_, _35796_);
  and (_28598_, _34659_, xram_data_in_reg[6]);
  and (_28599_, _34655_, xram_data_in[6]);
  or (_28601_, _28599_, _28598_);
  and (_00008_[6], _28601_, _35796_);
  nor (_28602_, _34655_, _24848_);
  and (_28603_, _34655_, xram_data_in[5]);
  or (_28604_, _28603_, _28602_);
  and (_00008_[5], _28604_, _35796_);
  and (_28605_, _34659_, xram_data_in_reg[4]);
  and (_28606_, _34655_, xram_data_in[4]);
  or (_28607_, _28606_, _28605_);
  and (_00008_[4], _28607_, _35796_);
  and (_28609_, _34659_, xram_data_in_reg[3]);
  and (_28610_, _34655_, xram_data_in[3]);
  or (_28611_, _28610_, _28609_);
  and (_00008_[3], _28611_, _35796_);
  and (_28612_, _34659_, xram_data_in_reg[2]);
  and (_28613_, _34655_, xram_data_in[2]);
  or (_28614_, _28613_, _28612_);
  and (_00008_[2], _28614_, _35796_);
  and (_28615_, _34659_, xram_data_in_reg[1]);
  and (_28616_, _34655_, xram_data_in[1]);
  or (_28618_, _28616_, _28615_);
  and (_00008_[1], _28618_, _35796_);
  and (_28619_, _34659_, xram_data_in_reg[0]);
  and (_28620_, _34655_, xram_data_in[0]);
  or (_28621_, _28620_, _28619_);
  and (_00008_[0], _28621_, _35796_);
  and (_28622_, _02976_, _02938_);
  and (_28623_, _28622_, _08997_);
  and (_28624_, _02986_, op0_cnst);
  and (_28625_, _09879_, _09250_);
  and (_28627_, _28625_, _28624_);
  and (_28628_, _02942_, _03041_);
  and (_28629_, _28628_, _28627_);
  and (_28630_, _28629_, _03224_);
  and (_28631_, _28630_, _28623_);
  and (_28632_, _28631_, _34655_);
  and (_28633_, _28632_, _35796_);
  and (_28634_, _27940_, _31024_);
  nor (_28635_, _27940_, _31024_);
  or (_28636_, _28635_, _28634_);
  and (_28638_, _10334_, _32130_);
  nor (_28639_, _10334_, _32130_);
  or (_28640_, _28639_, _28638_);
  or (_28641_, _28640_, _28636_);
  and (_28642_, _27804_, _32282_);
  nor (_28643_, _27804_, _32282_);
  and (_28644_, _27531_, _32176_);
  or (_28645_, _27158_, _32228_);
  nand (_28646_, _27158_, _32228_);
  and (_28647_, _28646_, _28645_);
  and (_28649_, _27283_, _32417_);
  nor (_28650_, _27283_, _32417_);
  or (_28651_, _28650_, _28649_);
  or (_28652_, _28651_, _28647_);
  nor (_28653_, _27531_, _32176_);
  or (_28654_, _28653_, _28652_);
  or (_28655_, _28654_, _28644_);
  nor (_28656_, _27406_, _31000_);
  and (_28657_, _27406_, _31000_);
  or (_28658_, _28657_, _28656_);
  nor (_28660_, _27667_, _32385_);
  and (_28661_, _27667_, _32385_);
  or (_28662_, _28661_, _28660_);
  or (_28663_, _28662_, _28658_);
  or (_28664_, _28663_, _28655_);
  or (_28665_, _28664_, _28643_);
  or (_28666_, _28665_, _28642_);
  or (_28667_, _28666_, _28641_);
  and (_00007_, _28667_, _28633_);
  nor (_28668_, _27074_, _30224_);
  and (_28670_, _27074_, _30224_);
  or (_28671_, _28670_, _28668_);
  nor (_28672_, _26568_, _31427_);
  and (_28673_, _26568_, _31427_);
  and (_28674_, _26675_, _32046_);
  nor (_28675_, _26675_, _32046_);
  not (_28676_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_28677_, _26891_, _28676_);
  or (_28678_, _28677_, _28675_);
  or (_28679_, _28678_, _28674_);
  and (_28681_, _26784_, _32405_);
  nor (_28682_, _26784_, _32405_);
  nor (_28683_, _26327_, _31392_);
  and (_28684_, _26327_, _31392_);
  or (_28685_, _28684_, _28683_);
  nor (_28686_, _26891_, _28676_);
  or (_28687_, _28686_, _28685_);
  or (_28688_, _28687_, _28682_);
  or (_28689_, _28688_, _28681_);
  or (_28690_, _28689_, _28679_);
  or (_28692_, _28690_, _28673_);
  or (_28693_, _28692_, _28672_);
  or (_28694_, _28693_, _28671_);
  and (_28695_, _10194_, _31375_);
  nor (_28696_, _10194_, _31375_);
  or (_28697_, _28696_, _28695_);
  or (_28698_, _28697_, _28694_);
  and (_00006_, _28698_, _28633_);
  or (_00001_, _28631_, rst);
  and (_00005_[7], _00617_, _35796_);
  and (_00004_[7], _00684_, _35796_);
  and (_00003_[7], _00554_, _35796_);
  and (_00002_[7], _00479_, _35796_);
  and (_28700_, _34659_, xram_data_in_reg[7]);
  and (_28701_, _34655_, xram_data_in[7]);
  or (_28702_, _28701_, _28700_);
  and (_00008_[7], _28702_, _35796_);
  and (_28703_, _02833_, _32243_);
  nor (_28704_, _02833_, _32243_);
  or (_28705_, _28704_, _28703_);
  not (_28707_, _32456_);
  nor (_28708_, _03687_, _28707_);
  and (_28709_, _03687_, _28707_);
  or (_28710_, _28709_, _28708_);
  or (_28711_, _28710_, _28705_);
  not (_28712_, _32295_);
  nor (_28713_, _03220_, _28712_);
  and (_28714_, _03220_, _28712_);
  or (_28715_, _28714_, _28713_);
  not (_28716_, _32398_);
  nor (_28717_, _03647_, _28716_);
  and (_28718_, _03647_, _28716_);
  or (_28719_, _28718_, _28717_);
  or (_28720_, _28719_, _28715_);
  or (_28721_, _28720_, _28711_);
  and (_28722_, _02794_, _32195_);
  nor (_28723_, _02794_, _32195_);
  or (_28724_, _28723_, _28722_);
  not (_28725_, _32347_);
  nor (_28726_, _03356_, _28725_);
  and (_28729_, _03356_, _28725_);
  or (_28730_, _28729_, _28726_);
  or (_28731_, _28730_, _28724_);
  and (_28732_, _02838_, _32122_);
  nor (_28733_, _02838_, _32122_);
  or (_28734_, _28733_, _28732_);
  nand (_28735_, _02924_, _32512_);
  or (_28736_, _02924_, _32512_);
  and (_28737_, _28736_, _28735_);
  or (_28738_, _28737_, _28734_);
  or (_28740_, _28738_, _28731_);
  or (_28741_, _28740_, _28721_);
  nor (_28742_, _35685_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_28743_, _28742_, _34815_);
  nor (_28744_, _09036_, _03056_);
  and (_28745_, _23122_, _03056_);
  nor (_28746_, _28745_, _28744_);
  not (_28747_, _28746_);
  nand (_28748_, _28747_, _28743_);
  and (_28749_, _34810_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_28751_, _28749_, _35264_);
  nor (_28752_, _28749_, _35264_);
  or (_28753_, _28752_, _28751_);
  or (_28754_, _09062_, _03056_);
  nand (_28755_, _21356_, _03056_);
  and (_28756_, _28755_, _28754_);
  or (_28757_, _28756_, _28753_);
  and (_28758_, _28757_, _28748_);
  not (_28759_, _35724_);
  and (_28760_, _23791_, _03056_);
  nor (_28762_, _09026_, _03056_);
  nor (_28763_, _28762_, _28760_);
  nand (_28764_, _28763_, _28759_);
  nor (_28765_, _34810_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_28766_, _28765_, _28749_);
  nor (_28767_, _09067_, _03056_);
  and (_28768_, _20994_, _03056_);
  nor (_28769_, _28768_, _28767_);
  or (_28770_, _28769_, _28766_);
  and (_28771_, _28770_, _28764_);
  and (_28773_, _28771_, _28758_);
  and (_28774_, _28749_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_28775_, _28774_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_28776_, _28774_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_28777_, _28776_, _28775_);
  nor (_28778_, _09054_, _03056_);
  and (_28779_, _21741_, _03056_);
  or (_28780_, _28779_, _28778_);
  or (_28781_, _28780_, _28777_);
  and (_28782_, _23445_, _03056_);
  nor (_28784_, _09031_, _03056_);
  nor (_28785_, _28784_, _28782_);
  nand (_28786_, _28785_, _35689_);
  and (_28787_, _28786_, _28781_);
  nor (_28788_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_28789_, _28788_, _34809_);
  or (_28790_, _28789_, _03060_);
  nand (_28791_, _28789_, _03060_);
  and (_28792_, _28791_, _28790_);
  and (_28793_, _28792_, _28787_);
  and (_28795_, _28793_, _28773_);
  nor (_28796_, _35684_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_28797_, _28796_, _35685_);
  nor (_28798_, _09044_, _03056_);
  and (_28799_, _22791_, _03056_);
  nor (_28800_, _28799_, _28798_);
  nand (_28801_, _28800_, _28797_);
  or (_28802_, _28800_, _28797_);
  and (_28803_, _28802_, _28801_);
  or (_28804_, _28747_, _28743_);
  or (_28806_, _28763_, _28759_);
  and (_28807_, _28806_, _28804_);
  and (_28808_, _28807_, _28803_);
  nand (_28809_, _28769_, _28766_);
  nand (_28810_, _03067_, _35245_);
  and (_28811_, _28810_, _28809_);
  or (_28812_, _28785_, _35689_);
  or (_28813_, _03067_, _35245_);
  and (_28814_, _28813_, _28812_);
  and (_28815_, _28814_, _28811_);
  and (_28817_, _28815_, _28808_);
  and (_28818_, _28817_, _28795_);
  or (_28819_, _35256_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_28820_, _34809_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_28821_, _28820_, _34810_);
  nand (_28822_, _28821_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_28823_, _28822_, _28819_);
  nand (_28824_, _28823_, _02663_);
  nor (_28825_, _08988_, _03056_);
  and (_28826_, _08802_, _03056_);
  nor (_28828_, _28826_, _28825_);
  nand (_28829_, _28828_, _34822_);
  or (_28830_, _28828_, _34822_);
  and (_28831_, _28830_, _28829_);
  and (_28832_, _28831_, _28824_);
  nor (_28833_, _09022_, _03056_);
  and (_28834_, _24077_, _03056_);
  nor (_28835_, _28834_, _28833_);
  nand (_28836_, _28835_, _35749_);
  or (_28837_, _28835_, _35749_);
  and (_28839_, _28837_, _28836_);
  nand (_28840_, _28821_, _03063_);
  or (_28841_, _28821_, _03063_);
  and (_28842_, _28841_, _28840_);
  and (_28843_, _28842_, _28839_);
  and (_28844_, _28843_, _28832_);
  and (_28845_, _34810_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_28846_, _28845_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_28847_, _28845_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_28848_, _28847_, _28846_);
  not (_28850_, _28848_);
  not (_28851_, _02537_);
  and (_28852_, _20994_, \oc8051_golden_model_1.ACC [4]);
  nor (_28853_, _20994_, \oc8051_golden_model_1.ACC [4]);
  nor (_28854_, _28853_, _28852_);
  nor (_28855_, _02630_, _02624_);
  nor (_28856_, _28855_, _02629_);
  nor (_28857_, _28856_, _28854_);
  and (_28858_, _28856_, _28854_);
  or (_28859_, _28858_, _28857_);
  or (_28861_, _28859_, _02609_);
  nand (_28862_, _02570_, _02609_);
  or (_28863_, _21182_, _02571_);
  nand (_28864_, _20996_, _02571_);
  or (_28865_, _28864_, _02605_);
  and (_28866_, _28865_, _28863_);
  or (_28867_, _28866_, _28862_);
  and (_28868_, _28867_, _28861_);
  or (_28869_, _28868_, _28851_);
  and (_28870_, _02611_, _02537_);
  or (_28872_, _09066_, _28870_);
  and (_28873_, _28872_, _28869_);
  nand (_28874_, _28873_, _28850_);
  nor (_28875_, \oc8051_golden_model_1.PC [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_28876_, \oc8051_golden_model_1.PC [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_28877_, _28876_, _28875_);
  or (_28878_, _28877_, _03065_);
  nor (_28879_, _02304_, _30692_);
  and (_28880_, _02304_, _30692_);
  or (_28881_, _28880_, _28879_);
  nor (_28883_, _02273_, _30669_);
  and (_28884_, _02273_, _30669_);
  or (_28885_, _28884_, _28883_);
  or (_28886_, _28885_, _28881_);
  or (_28887_, _02506_, _30590_);
  nand (_28888_, _02506_, _30590_);
  and (_28889_, _28888_, _28887_);
  or (_28890_, _02501_, _30520_);
  or (_28891_, _02464_, _35181_);
  and (_28892_, _28891_, _28890_);
  or (_28893_, _28892_, _28889_);
  or (_28894_, _28893_, _28886_);
  and (_28895_, _02367_, _30643_);
  nor (_28896_, _02367_, _30643_);
  or (_28897_, _28896_, _28895_);
  nand (_28898_, _02336_, _30617_);
  or (_28899_, _02336_, _30617_);
  and (_28900_, _28899_, _28898_);
  or (_28901_, _28900_, _28897_);
  and (_28902_, _02513_, _30567_);
  nor (_28904_, _02513_, _30567_);
  or (_28905_, _28904_, _28902_);
  not (_28906_, _02432_);
  nor (_28907_, _28906_, _30545_);
  and (_28908_, _28906_, _30545_);
  or (_28909_, _28908_, _28907_);
  or (_28910_, _28909_, _28905_);
  or (_28911_, _28910_, _28901_);
  or (_28912_, _28911_, _28894_);
  nor (_28913_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_28915_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_28916_, _28915_, _28913_);
  nor (_28917_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_28918_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_28919_, _28918_, _28917_);
  and (_28920_, _28919_, _28916_);
  or (_28921_, \oc8051_golden_model_1.PC [12], _31059_);
  or (_28922_, _23794_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_28923_, _28922_, _28921_);
  nand (_28924_, \oc8051_golden_model_1.PC [13], _31034_);
  or (_28926_, \oc8051_golden_model_1.PC [13], _31034_);
  and (_28927_, _28926_, _28924_);
  and (_28928_, _28927_, _28923_);
  and (_28929_, _28928_, _28920_);
  and (_28930_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_28931_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_28932_, _28931_, _28930_);
  nor (_28933_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_28934_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_28935_, _28934_, _28933_);
  and (_28937_, _28935_, _28932_);
  and (_28938_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_28939_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_28940_, _28939_, _28938_);
  nor (_28941_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_28942_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_28943_, _28942_, _28941_);
  and (_28944_, _28943_, _28940_);
  and (_28945_, _28944_, _28937_);
  and (_28946_, _28945_, _28929_);
  or (_28948_, \oc8051_golden_model_1.PC [0], _35245_);
  or (_28949_, _02247_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_28950_, _28949_, _28948_);
  nor (_28951_, _28950_, _28877_);
  and (_28952_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_28953_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_28954_, _28953_, _28952_);
  or (_28955_, \oc8051_golden_model_1.PC [3], _35256_);
  or (_28956_, _02216_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_28957_, _28956_, _28955_);
  and (_28959_, _28957_, _28954_);
  and (_28960_, _28959_, _28951_);
  or (_28961_, \oc8051_golden_model_1.PC [4], _35260_);
  or (_28962_, _20991_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_28963_, _28962_, _28961_);
  nand (_28964_, \oc8051_golden_model_1.PC [5], _35264_);
  or (_28965_, \oc8051_golden_model_1.PC [5], _35264_);
  and (_28966_, _28965_, _28964_);
  and (_28967_, _28966_, _28963_);
  or (_28968_, \oc8051_golden_model_1.PC [6], _35268_);
  or (_28970_, _21757_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_28971_, _28970_, _28968_);
  and (_28972_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_28973_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_28974_, _28973_, _28972_);
  and (_28975_, _28974_, _28971_);
  and (_28976_, _28975_, _28967_);
  and (_28977_, _28976_, _28960_);
  and (_28978_, _28977_, _28946_);
  and (_28979_, _28978_, _34655_);
  and (_28981_, _28979_, _28912_);
  and (_28982_, _28981_, _28878_);
  and (_28983_, _28982_, _28874_);
  or (_28984_, _28873_, _28850_);
  or (_28985_, _28823_, _02663_);
  and (_28986_, _28985_, _28984_);
  and (_28987_, _28986_, _28983_);
  and (_28988_, _28987_, _28844_);
  and (_28989_, _28988_, _28818_);
  and (_28990_, _28845_, _34813_);
  and (_28992_, _28990_, _34930_);
  and (_28993_, _28992_, _31059_);
  nor (_28994_, _28992_, _31059_);
  or (_28995_, _28994_, _28993_);
  nor (_28996_, _23922_, _02571_);
  not (_28997_, _02570_);
  and (_28998_, _23791_, _02610_);
  and (_28999_, _09027_, _02605_);
  nor (_29000_, _28999_, _28998_);
  nor (_29001_, _29000_, _07721_);
  nor (_29003_, _29001_, _28997_);
  not (_29004_, _29003_);
  nor (_29005_, _29004_, _28996_);
  nor (_29006_, _09027_, _02570_);
  or (_29007_, _29006_, _02542_);
  nor (_29008_, _29007_, _29005_);
  and (_29009_, _22093_, \oc8051_golden_model_1.ACC [7]);
  nor (_29010_, _22093_, \oc8051_golden_model_1.ACC [7]);
  nor (_29011_, _29010_, _29009_);
  and (_29012_, _21738_, \oc8051_golden_model_1.ACC [6]);
  nor (_29014_, _21738_, \oc8051_golden_model_1.ACC [6]);
  nor (_29015_, _29014_, _29012_);
  and (_29016_, _21356_, \oc8051_golden_model_1.ACC [5]);
  nor (_29017_, _21356_, \oc8051_golden_model_1.ACC [5]);
  nor (_29018_, _29017_, _29016_);
  and (_29019_, _29018_, _28852_);
  nor (_29020_, _29019_, _29016_);
  not (_29021_, _28856_);
  and (_29022_, _29018_, _28854_);
  nand (_29023_, _29022_, _29021_);
  nand (_29025_, _29023_, _29020_);
  and (_29026_, _29025_, _29015_);
  or (_29027_, _29026_, _29012_);
  and (_29028_, _29027_, _29011_);
  nor (_29029_, _29028_, _29009_);
  and (_29030_, _22791_, _22468_);
  and (_29031_, _23445_, _23119_);
  and (_29032_, _29031_, _29030_);
  not (_29033_, _29032_);
  nor (_29034_, _29033_, _29029_);
  and (_29036_, _29034_, _23776_);
  nor (_29037_, _29034_, _23776_);
  nor (_29038_, _29037_, _29036_);
  nor (_29039_, _29038_, _02609_);
  or (_29040_, _29039_, _28851_);
  nor (_29041_, _29040_, _29008_);
  nor (_29042_, _09027_, _02537_);
  or (_29043_, _29042_, _29041_);
  and (_29044_, _29043_, _28995_);
  nor (_29045_, _29043_, _28995_);
  or (_29047_, _29045_, _29044_);
  or (_29048_, _03505_, _34547_);
  nand (_29049_, _03505_, _34547_);
  and (_29050_, _29049_, _29048_);
  or (_29051_, _03720_, _34564_);
  nand (_29052_, _03720_, _34564_);
  and (_29053_, _29052_, _29051_);
  or (_29054_, _29053_, _29050_);
  or (_29055_, _05649_, _34632_);
  nand (_29056_, _05649_, _34632_);
  and (_29058_, _29056_, _29055_);
  not (_29059_, _34615_);
  nor (_29060_, _05617_, _29059_);
  and (_29061_, _05617_, _29059_);
  or (_29062_, _29061_, _29060_);
  or (_29063_, _29062_, _29058_);
  or (_29064_, _29063_, _29054_);
  not (_29065_, _34598_);
  nor (_29066_, _03128_, _29065_);
  and (_29067_, _03128_, _29065_);
  or (_29069_, _29067_, _29066_);
  nand (_29070_, _03262_, _34581_);
  or (_29071_, _03262_, _34581_);
  and (_29072_, _29071_, _29070_);
  or (_29073_, _29072_, _29069_);
  or (_29074_, _05302_, _34530_);
  nand (_29075_, _05302_, _34530_);
  and (_29076_, _29075_, _29074_);
  nand (_29077_, _05585_, _34649_);
  or (_29078_, _05585_, _34649_);
  and (_29080_, _29078_, _29077_);
  or (_29081_, _29080_, _29076_);
  or (_29082_, _29081_, _29073_);
  or (_29083_, _29082_, _29064_);
  and (_29084_, _29083_, _29047_);
  and (_29085_, _28992_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_29086_, _29085_, _31034_);
  nor (_29087_, _29085_, _31034_);
  or (_29088_, _29087_, _29086_);
  not (_29089_, _29088_);
  and (_29091_, _24240_, _07721_);
  and (_29092_, _24077_, _02610_);
  and (_29093_, _09021_, _02605_);
  nor (_29094_, _29093_, _29092_);
  nor (_29095_, _29094_, _07721_);
  or (_29096_, _29095_, _28997_);
  nor (_29097_, _29096_, _29091_);
  nor (_29098_, _09021_, _02570_);
  nor (_29099_, _29098_, _02542_);
  not (_29100_, _29099_);
  nor (_29102_, _29100_, _29097_);
  and (_29103_, _29036_, _24129_);
  nor (_29104_, _29036_, _24129_);
  or (_29105_, _29104_, _29103_);
  and (_29106_, _29105_, _02542_);
  nor (_29107_, _29106_, _29102_);
  nor (_29108_, _29107_, _28851_);
  nor (_29109_, _09022_, _02537_);
  or (_29110_, _29109_, _29108_);
  nand (_29111_, _29110_, _29089_);
  or (_29113_, _29110_, _29089_);
  and (_29114_, _29113_, _29111_);
  and (_29115_, _29114_, _29084_);
  and (_29116_, _29115_, _28989_);
  and (property_invalid_rom_pc, _29116_, _28741_);
  nor (_29117_, _30980_, \oc8051_golden_model_1.SP [7]);
  and (_29118_, _30980_, \oc8051_golden_model_1.SP [7]);
  or (_29119_, _29118_, _29117_);
  nor (_29120_, _31024_, \oc8051_golden_model_1.SP [6]);
  and (_29121_, _31024_, \oc8051_golden_model_1.SP [6]);
  or (_29123_, _29121_, _29120_);
  and (_29124_, _31018_, \oc8051_golden_model_1.SP [5]);
  nor (_29125_, _31018_, \oc8051_golden_model_1.SP [5]);
  or (_29126_, _29125_, _29124_);
  and (_29127_, _31006_, \oc8051_golden_model_1.SP [3]);
  nor (_29128_, _31006_, \oc8051_golden_model_1.SP [3]);
  or (_29129_, _29128_, _29127_);
  and (_29130_, _31000_, \oc8051_golden_model_1.SP [2]);
  or (_29131_, _30988_, _02868_);
  nand (_29132_, _30988_, _02868_);
  and (_29134_, _29132_, _29131_);
  nor (_29135_, _30994_, \oc8051_golden_model_1.SP [1]);
  and (_29136_, _30994_, \oc8051_golden_model_1.SP [1]);
  or (_29137_, _29136_, _29135_);
  or (_29138_, _29137_, _29134_);
  nor (_29139_, _31000_, \oc8051_golden_model_1.SP [2]);
  or (_29140_, _29139_, _29138_);
  or (_29141_, _29140_, _29130_);
  or (_29142_, _29141_, _29129_);
  and (_29143_, _31012_, \oc8051_golden_model_1.SP [4]);
  nor (_29145_, _31012_, \oc8051_golden_model_1.SP [4]);
  or (_29146_, _29145_, _29143_);
  or (_29147_, _29146_, _29142_);
  or (_29148_, _29147_, _29126_);
  or (_29149_, _29148_, _29123_);
  or (_29150_, _29149_, _29119_);
  and (_29151_, _28631_, inst_finished_r);
  and (_29152_, _29151_, property_invalid_sp_1_r);
  and (property_invalid_sp, _29152_, _29150_);
  nand (_29153_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_29155_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_29156_, _29155_, _29153_);
  and (_29157_, _26229_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_29158_, \oc8051_golden_model_1.PSW [1], _31392_);
  or (_29159_, _29158_, _29157_);
  or (_29160_, _29159_, _29156_);
  and (_29161_, _26679_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_29162_, \oc8051_golden_model_1.PSW [4], _32405_);
  or (_29163_, _29162_, _29161_);
  and (_29164_, _02974_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_29166_, \oc8051_golden_model_1.PSW [3], _32046_);
  or (_29167_, _29166_, _29164_);
  or (_29168_, _29167_, _29163_);
  or (_29169_, _29168_, _29160_);
  and (_29170_, _07288_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_29171_, \oc8051_golden_model_1.PSW [7], _31375_);
  or (_29172_, _29171_, _29170_);
  and (_29173_, _26788_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_29174_, \oc8051_golden_model_1.PSW [5], _28676_);
  or (_29175_, _29174_, _29173_);
  nand (_29177_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_29178_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_29179_, _29178_, _29177_);
  or (_29180_, _29179_, _29175_);
  or (_29181_, _29180_, _29172_);
  or (_29182_, _29181_, _29169_);
  and (_29183_, _29182_, property_invalid_psw_1_r);
  and (property_invalid_psw, _29183_, _29151_);
  or (_29184_, _28055_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  nand (_29185_, _28055_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  and (_29187_, _29185_, _29184_);
  or (_29188_, _28123_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  nand (_29189_, _28123_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  and (_29190_, _29189_, _29188_);
  or (_29191_, _29190_, _29187_);
  or (_29192_, _28198_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  nand (_29193_, _28198_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  and (_29194_, _29193_, _29192_);
  or (_29195_, _28232_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  nand (_29196_, _28232_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  and (_29198_, _29196_, _29195_);
  or (_29199_, _29198_, _29194_);
  or (_29200_, _29199_, _29191_);
  nor (_29201_, _28145_, _00237_);
  and (_29202_, _28145_, _00237_);
  or (_29203_, _29202_, _29201_);
  nor (_29204_, _10339_, _35217_);
  and (_29205_, _10339_, _35217_);
  or (_29206_, _29205_, _29204_);
  or (_29207_, _29206_, _29203_);
  nor (_29209_, _28091_, _00227_);
  and (_29210_, _28091_, _00227_);
  or (_29211_, _29210_, _29209_);
  nor (_29212_, _28171_, _00242_);
  and (_29213_, _28171_, _00242_);
  or (_29214_, _29213_, _29212_);
  or (_29215_, _29214_, _29211_);
  or (_29216_, _29215_, _29207_);
  or (_29217_, _29216_, _29200_);
  and (property_invalid_xram_data_out, _29217_, _28632_);
  or (_29219_, _28343_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  nand (_29220_, _28343_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  and (_29221_, _29220_, _29219_);
  or (_29222_, _28312_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  nand (_29223_, _28312_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  and (_29224_, _29223_, _29222_);
  nor (_29225_, _28359_, _00299_);
  and (_29226_, _28359_, _00299_);
  or (_29227_, _29226_, _29225_);
  or (_29228_, _29227_, _29224_);
  or (_29230_, _29228_, _29221_);
  and (_29231_, _28328_, _00285_);
  nor (_29232_, _28297_, _00271_);
  nor (_29233_, _28374_, _00306_);
  or (_29234_, _29233_, _29232_);
  or (_29235_, _29234_, _29231_);
  or (_29236_, _28281_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  nand (_29237_, _28281_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  and (_29238_, _29237_, _29236_);
  nor (_29239_, _28435_, _00323_);
  and (_29241_, _28435_, _00323_);
  or (_29242_, _29241_, _29239_);
  nor (_29243_, _28529_, _00343_);
  and (_29244_, _28529_, _00343_);
  or (_29245_, _29244_, _29243_);
  or (_29246_, _29245_, _29242_);
  nor (_29247_, _28495_, _00338_);
  and (_29248_, _28495_, _00338_);
  or (_29249_, _29248_, _29247_);
  nor (_29250_, _28405_, _00318_);
  and (_29252_, _28381_, _00313_);
  or (_29253_, _29252_, _29250_);
  or (_29254_, _29253_, _29249_);
  or (_29255_, _29254_, _29246_);
  nor (_29256_, _10346_, _35227_);
  and (_29257_, _10346_, _35227_);
  or (_29258_, _29257_, _29256_);
  nor (_29259_, _28484_, _00333_);
  and (_29260_, _28484_, _00333_);
  or (_29261_, _29260_, _29259_);
  or (_29262_, _29261_, _29258_);
  nor (_29263_, _28454_, _00328_);
  and (_29264_, _28454_, _00328_);
  or (_29265_, _29264_, _29263_);
  nor (_29266_, _28381_, _00313_);
  and (_29267_, _28405_, _00318_);
  or (_29268_, _29267_, _29266_);
  or (_29269_, _29268_, _29265_);
  or (_29270_, _29269_, _29262_);
  or (_29271_, _29270_, _29255_);
  nor (_29274_, _28265_, _00257_);
  or (_29275_, _29274_, _29271_);
  or (_29276_, _29275_, _29238_);
  and (_29277_, _28265_, _00257_);
  and (_29278_, _28297_, _00271_);
  or (_29279_, _29278_, _29277_);
  nor (_29280_, _28328_, _00285_);
  and (_29281_, _28374_, _00306_);
  or (_29282_, _29281_, _29280_);
  or (_29283_, _29282_, _29279_);
  or (_29285_, _29283_, _29276_);
  or (_29286_, _29285_, _29235_);
  or (_29287_, _29286_, _29230_);
  and (property_invalid_xram_addr, _29287_, _28632_);
  nand (_29288_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_29289_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_29290_, _29289_, _29288_);
  and (_29291_, _19057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_29292_, \oc8051_golden_model_1.P3 [2], _31960_);
  or (_29293_, _29292_, _29291_);
  or (_29295_, _29293_, _29290_);
  and (_29296_, \oc8051_golden_model_1.P3 [0], _31934_);
  and (_29297_, _18846_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_29298_, _29297_, _29296_);
  and (_29299_, _18948_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_29300_, \oc8051_golden_model_1.P3 [1], _31949_);
  or (_29301_, _29300_, _29299_);
  or (_29302_, _29301_, _29298_);
  or (_29303_, _29302_, _29295_);
  or (_29304_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_29306_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_29307_, _29306_, _29304_);
  or (_29308_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_29309_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_29310_, _29309_, _29308_);
  or (_29311_, _29310_, _29307_);
  and (_29312_, _08687_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_29313_, \oc8051_golden_model_1.P3 [7], _31648_);
  or (_29314_, _29313_, _29312_);
  nand (_29315_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_29317_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_29318_, _29317_, _29315_);
  or (_29319_, _29318_, _29314_);
  or (_29320_, _29319_, _29311_);
  or (_29321_, _29320_, _29303_);
  and (property_invalid_p3, _29321_, _29151_);
  nand (_29322_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_29323_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_29324_, _29323_, _29322_);
  and (_29325_, _18309_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_29327_, \oc8051_golden_model_1.P2 [2], _31874_);
  or (_29328_, _29327_, _29325_);
  or (_29329_, _29328_, _29324_);
  and (_29330_, \oc8051_golden_model_1.P2 [0], _31848_);
  and (_29331_, _18097_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_29332_, _29331_, _29330_);
  and (_29333_, _18200_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_29334_, \oc8051_golden_model_1.P2 [1], _31861_);
  or (_29335_, _29334_, _29333_);
  or (_29336_, _29335_, _29332_);
  or (_29338_, _29336_, _29329_);
  or (_29339_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_29340_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_29341_, _29340_, _29339_);
  or (_29342_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_29343_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_29344_, _29343_, _29342_);
  or (_29345_, _29344_, _29341_);
  and (_29346_, _08588_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_29347_, \oc8051_golden_model_1.P2 [7], _31640_);
  or (_29349_, _29347_, _29346_);
  nand (_29350_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_29351_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_29352_, _29351_, _29350_);
  or (_29353_, _29352_, _29349_);
  or (_29354_, _29353_, _29345_);
  or (_29355_, _29354_, _29338_);
  and (property_invalid_p2, _29355_, _29151_);
  nand (_29356_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_29357_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_29359_, _29357_, _29356_);
  and (_29360_, _17560_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_29361_, \oc8051_golden_model_1.P1 [2], _31787_);
  or (_29362_, _29361_, _29360_);
  or (_29363_, _29362_, _29359_);
  and (_29364_, \oc8051_golden_model_1.P1 [0], _31761_);
  and (_29365_, _17349_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_29366_, _29365_, _29364_);
  and (_29367_, _17451_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_29368_, \oc8051_golden_model_1.P1 [1], _31774_);
  or (_29370_, _29368_, _29367_);
  or (_29371_, _29370_, _29366_);
  or (_29372_, _29371_, _29363_);
  or (_29373_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_29374_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_29375_, _29374_, _29373_);
  or (_29376_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_29377_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_29378_, _29377_, _29376_);
  or (_29379_, _29378_, _29375_);
  and (_29381_, _08489_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_29382_, \oc8051_golden_model_1.P1 [7], _31622_);
  or (_29383_, _29382_, _29381_);
  nand (_29384_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_29385_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_29386_, _29385_, _29384_);
  or (_29387_, _29386_, _29383_);
  or (_29388_, _29387_, _29379_);
  or (_29389_, _29388_, _29372_);
  and (property_invalid_p1, _29389_, _29151_);
  nand (_29391_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_29392_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_29393_, _29392_, _29391_);
  and (_29394_, _16804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_29395_, \oc8051_golden_model_1.P0 [2], _31698_);
  or (_29396_, _29395_, _29394_);
  or (_29397_, _29396_, _29393_);
  and (_29398_, \oc8051_golden_model_1.P0 [0], _31671_);
  and (_29399_, _16590_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_29400_, _29399_, _29398_);
  and (_29402_, _16694_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_29403_, \oc8051_golden_model_1.P0 [1], _31682_);
  or (_29404_, _29403_, _29402_);
  or (_29405_, _29404_, _29400_);
  or (_29406_, _29405_, _29397_);
  or (_29407_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_29408_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_29409_, _29408_, _29407_);
  or (_29410_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_29411_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_29413_, _29411_, _29410_);
  or (_29414_, _29413_, _29409_);
  and (_29415_, _08389_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_29416_, \oc8051_golden_model_1.P0 [7], _31609_);
  or (_29417_, _29416_, _29415_);
  nand (_29418_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_29419_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_29420_, _29419_, _29418_);
  or (_29421_, _29420_, _29417_);
  or (_29422_, _29421_, _29414_);
  or (_29424_, _29422_, _29406_);
  and (property_invalid_p0, _29424_, _29151_);
  or (_29425_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_29426_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_29427_, _29426_, _29425_);
  nand (_29428_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_29429_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_29430_, _29429_, _29428_);
  or (_29431_, _29430_, _29427_);
  and (_29432_, _03370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_29434_, \oc8051_golden_model_1.IRAM[0] [0], _32604_);
  or (_29435_, _29434_, _29432_);
  and (_29436_, _03965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_29437_, \oc8051_golden_model_1.IRAM[0] [1], _32608_);
  or (_29438_, _29437_, _29436_);
  or (_29439_, _29438_, _29435_);
  or (_29440_, _29439_, _29431_);
  or (_29441_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand (_29442_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_29443_, _29442_, _29441_);
  nand (_29445_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_29446_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_29447_, _29446_, _29445_);
  or (_29448_, _29447_, _29443_);
  or (_29449_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_29450_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_29451_, _29450_, _29449_);
  or (_29452_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_29453_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_29454_, _29453_, _29452_);
  or (_29456_, _29454_, _29451_);
  or (_29457_, _29456_, _29448_);
  or (_29458_, _29457_, _29440_);
  or (_29459_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_29460_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_29461_, _29460_, _29459_);
  or (_29462_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_29463_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_29464_, _29463_, _29462_);
  or (_29465_, _29464_, _29461_);
  or (_29467_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand (_29468_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_29469_, _29468_, _29467_);
  nand (_29470_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_29471_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_29472_, _29471_, _29470_);
  or (_29473_, _29472_, _29469_);
  or (_29474_, _29473_, _29465_);
  and (_29475_, _05139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_29476_, \oc8051_golden_model_1.IRAM[1] [4], _32640_);
  or (_29478_, _29476_, _29475_);
  and (_29479_, _04840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_29480_, \oc8051_golden_model_1.IRAM[1] [5], _32643_);
  or (_29481_, _29480_, _29479_);
  or (_29482_, _29481_, _29478_);
  or (_29483_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand (_29484_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_29485_, _29484_, _29483_);
  nand (_29486_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_29487_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_29489_, _29487_, _29486_);
  or (_29490_, _29489_, _29485_);
  or (_29491_, _29490_, _29482_);
  or (_29492_, _29491_, _29474_);
  or (_29493_, _29492_, _29458_);
  or (_29494_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand (_29495_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_29496_, _29495_, _29494_);
  or (_29497_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand (_29498_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_29500_, _29498_, _29497_);
  or (_29501_, _29500_, _29496_);
  nand (_29502_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_29503_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_29504_, _29503_, _29502_);
  and (_29505_, _04401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_29506_, \oc8051_golden_model_1.IRAM[2] [2], _32658_);
  or (_29507_, _29506_, _29505_);
  or (_29508_, _29507_, _29504_);
  or (_29509_, _29508_, _29501_);
  and (_29511_, _05144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_29512_, \oc8051_golden_model_1.IRAM[2] [4], _32663_);
  or (_29513_, _29512_, _29511_);
  and (_29514_, _04845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_29515_, \oc8051_golden_model_1.IRAM[2] [5], _32666_);
  or (_29516_, _29515_, _29514_);
  or (_29517_, _29516_, _29513_);
  and (_29518_, _04579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_29519_, \oc8051_golden_model_1.IRAM[2] [7], _32672_);
  or (_29520_, _29519_, _29518_);
  nand (_29521_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_29522_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_29523_, _29522_, _29521_);
  or (_29524_, _29523_, _29520_);
  or (_29525_, _29524_, _29517_);
  or (_29526_, _29525_, _29509_);
  and (_29527_, \oc8051_golden_model_1.IRAM[3] [2], _32682_);
  and (_29528_, _04399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_29529_, _29528_, _29527_);
  nand (_29530_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_29533_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_29534_, _29533_, _29530_);
  or (_29535_, _29534_, _29529_);
  and (_29536_, _03784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_29537_, \oc8051_golden_model_1.IRAM[3] [0], _32676_);
  or (_29538_, _29537_, _29536_);
  and (_29539_, _03970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_29540_, \oc8051_golden_model_1.IRAM[3] [1], _32679_);
  or (_29541_, _29540_, _29539_);
  or (_29542_, _29541_, _29538_);
  or (_29544_, _29542_, _29535_);
  nand (_29545_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_29546_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_29547_, _29546_, _29545_);
  and (_29548_, _04577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_29549_, \oc8051_golden_model_1.IRAM[3] [7], _32537_);
  or (_29550_, _29549_, _29548_);
  or (_29551_, _29550_, _29547_);
  or (_29552_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_29553_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_29554_, _29553_, _29552_);
  or (_29555_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_29556_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_29557_, _29556_, _29555_);
  or (_29558_, _29557_, _29554_);
  or (_29559_, _29558_, _29551_);
  or (_29560_, _29559_, _29544_);
  or (_29561_, _29560_, _29526_);
  or (_29562_, _29561_, _29493_);
  and (_29563_, _03800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_29565_, \oc8051_golden_model_1.IRAM[4] [0], _32699_);
  or (_29566_, _29565_, _29563_);
  and (_29567_, \oc8051_golden_model_1.IRAM[4] [1], _32702_);
  and (_29568_, _03984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_29569_, _29568_, _29567_);
  or (_29570_, _29569_, _29566_);
  or (_29571_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand (_29572_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_29573_, _29572_, _29571_);
  nand (_29574_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_29576_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_29577_, _29576_, _29574_);
  or (_29578_, _29577_, _29573_);
  or (_29579_, _29578_, _29570_);
  or (_29580_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand (_29581_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_29582_, _29581_, _29580_);
  or (_29583_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand (_29584_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_29585_, _29584_, _29583_);
  or (_29587_, _29585_, _29582_);
  or (_29588_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand (_29589_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_29590_, _29589_, _29588_);
  nand (_29591_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_29592_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_29593_, _29592_, _29591_);
  or (_29594_, _29593_, _29590_);
  or (_29595_, _29594_, _29587_);
  or (_29596_, _29595_, _29579_);
  or (_29598_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand (_29599_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_29600_, _29599_, _29598_);
  or (_29601_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand (_29602_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_29603_, _29602_, _29601_);
  or (_29604_, _29603_, _29600_);
  or (_29605_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_29606_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_29607_, _29606_, _29605_);
  or (_29609_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_29610_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_29611_, _29610_, _29609_);
  or (_29612_, _29611_, _29607_);
  or (_29613_, _29612_, _29604_);
  or (_29614_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand (_29615_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_29616_, _29615_, _29614_);
  or (_29617_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nand (_29618_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_29620_, _29618_, _29617_);
  or (_29621_, _29620_, _29616_);
  and (_29622_, \oc8051_golden_model_1.IRAM[5] [4], _32729_);
  and (_29623_, _05158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_29624_, _29623_, _29622_);
  and (_29625_, \oc8051_golden_model_1.IRAM[5] [5], _32732_);
  and (_29626_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_29627_, _29626_, _29625_);
  or (_29628_, _29627_, _29624_);
  or (_29629_, _29628_, _29621_);
  or (_29631_, _29629_, _29613_);
  or (_29632_, _29631_, _29596_);
  or (_29633_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nand (_29634_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_29635_, _29634_, _29633_);
  and (_29636_, \oc8051_golden_model_1.IRAM[6] [2], _32745_);
  and (_29637_, _04409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_29638_, _29637_, _29636_);
  or (_29639_, _29638_, _29635_);
  or (_29640_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand (_29642_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_29643_, _29642_, _29640_);
  or (_29644_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand (_29645_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_29646_, _29645_, _29644_);
  or (_29647_, _29646_, _29643_);
  or (_29648_, _29647_, _29639_);
  or (_29649_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nand (_29650_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_29651_, _29650_, _29649_);
  and (_29653_, _04588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_29654_, \oc8051_golden_model_1.IRAM[6] [7], _32758_);
  or (_29655_, _29654_, _29653_);
  or (_29656_, _29655_, _29651_);
  and (_29657_, \oc8051_golden_model_1.IRAM[6] [5], _32753_);
  and (_29658_, _04853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_29659_, _29658_, _29657_);
  and (_29660_, _05152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_29661_, \oc8051_golden_model_1.IRAM[6] [4], _32750_);
  or (_29662_, _29661_, _29660_);
  or (_29664_, _29662_, _29659_);
  or (_29665_, _29664_, _29656_);
  or (_29666_, _29665_, _29648_);
  and (_29667_, _03978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_29668_, \oc8051_golden_model_1.IRAM[7] [1], _32765_);
  or (_29669_, _29668_, _29667_);
  and (_29670_, _03794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_29671_, \oc8051_golden_model_1.IRAM[7] [0], _32762_);
  or (_29672_, _29671_, _29670_);
  or (_29673_, _29672_, _29669_);
  and (_29675_, _04407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_29676_, \oc8051_golden_model_1.IRAM[7] [2], _32768_);
  or (_29677_, _29676_, _29675_);
  nand (_29678_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_29679_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_29680_, _29679_, _29678_);
  or (_29681_, _29680_, _29677_);
  or (_29682_, _29681_, _29673_);
  or (_29683_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_29684_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_29686_, _29684_, _29683_);
  or (_29687_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_29688_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_29689_, _29688_, _29687_);
  or (_29690_, _29689_, _29686_);
  and (_29691_, _04586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_29692_, \oc8051_golden_model_1.IRAM[7] [7], _32549_);
  or (_29693_, _29692_, _29691_);
  nand (_29694_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_29695_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_29697_, _29695_, _29694_);
  or (_29698_, _29697_, _29693_);
  or (_29699_, _29698_, _29690_);
  or (_29700_, _29699_, _29682_);
  or (_29701_, _29700_, _29666_);
  or (_29702_, _29701_, _29632_);
  or (_29703_, _29702_, _29562_);
  and (_29704_, _03999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_29705_, \oc8051_golden_model_1.IRAM[8] [1], _32788_);
  or (_29706_, _29705_, _29704_);
  and (_29708_, _03817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_29709_, \oc8051_golden_model_1.IRAM[8] [0], _32785_);
  or (_29710_, _29709_, _29708_);
  or (_29711_, _29710_, _29706_);
  or (_29712_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand (_29713_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_29714_, _29713_, _29712_);
  nand (_29715_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_29716_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_29717_, _29716_, _29715_);
  or (_29719_, _29717_, _29714_);
  or (_29720_, _29719_, _29711_);
  or (_29721_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand (_29722_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_29723_, _29722_, _29721_);
  or (_29724_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand (_29725_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_29726_, _29725_, _29724_);
  or (_29727_, _29726_, _29723_);
  or (_29728_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_29730_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_29731_, _29730_, _29728_);
  nand (_29732_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_29733_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_29734_, _29733_, _29732_);
  or (_29735_, _29734_, _29731_);
  or (_29736_, _29735_, _29727_);
  or (_29737_, _29736_, _29720_);
  or (_29738_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand (_29739_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_29741_, _29739_, _29738_);
  nand (_29742_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_29743_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_29744_, _29743_, _29742_);
  or (_29745_, _29744_, _29741_);
  or (_29746_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand (_29747_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_29748_, _29747_, _29746_);
  or (_29749_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand (_29750_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_29752_, _29750_, _29749_);
  or (_29753_, _29752_, _29748_);
  or (_29754_, _29753_, _29745_);
  or (_29755_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand (_29756_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_29757_, _29756_, _29755_);
  nand (_29758_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_29759_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_29760_, _29759_, _29758_);
  or (_29761_, _29760_, _29757_);
  and (_29763_, _05172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_29764_, \oc8051_golden_model_1.IRAM[9] [4], _32816_);
  or (_29765_, _29764_, _29763_);
  and (_29766_, _04873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_29767_, \oc8051_golden_model_1.IRAM[9] [5], _32819_);
  or (_29768_, _29767_, _29766_);
  or (_29769_, _29768_, _29765_);
  or (_29770_, _29769_, _29761_);
  or (_29771_, _29770_, _29754_);
  or (_29772_, _29771_, _29737_);
  and (_29774_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_29775_, \oc8051_golden_model_1.IRAM[10] [2], _32832_);
  or (_29776_, _29775_, _29774_);
  nand (_29777_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_29778_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_29779_, _29778_, _29777_);
  or (_29780_, _29779_, _29776_);
  or (_29781_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nand (_29782_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_29783_, _29782_, _29781_);
  or (_29785_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nand (_29786_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_29787_, _29786_, _29785_);
  or (_29788_, _29787_, _29783_);
  or (_29789_, _29788_, _29780_);
  and (_29790_, _04604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_29791_, \oc8051_golden_model_1.IRAM[10] [7], _32563_);
  or (_29792_, _29791_, _29790_);
  nand (_29793_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_29794_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_29796_, _29794_, _29793_);
  or (_29797_, _29796_, _29792_);
  and (_29798_, _05167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_29799_, \oc8051_golden_model_1.IRAM[10] [4], _32838_);
  or (_29800_, _29799_, _29798_);
  and (_29801_, \oc8051_golden_model_1.IRAM[10] [5], _32841_);
  and (_29802_, _04868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_29803_, _29802_, _29801_);
  or (_29804_, _29803_, _29800_);
  or (_29805_, _29804_, _29797_);
  or (_29807_, _29805_, _29789_);
  and (_29808_, _03811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_29809_, \oc8051_golden_model_1.IRAM[11] [0], _32850_);
  or (_29810_, _29809_, _29808_);
  and (_29811_, _03994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_29812_, \oc8051_golden_model_1.IRAM[11] [1], _32853_);
  or (_29813_, _29812_, _29811_);
  or (_29814_, _29813_, _29810_);
  and (_29815_, _04423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_29816_, \oc8051_golden_model_1.IRAM[11] [2], _32856_);
  or (_29818_, _29816_, _29815_);
  nand (_29819_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_29820_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_29821_, _29820_, _29819_);
  or (_29822_, _29821_, _29818_);
  or (_29823_, _29822_, _29814_);
  or (_29824_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_29825_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_29826_, _29825_, _29824_);
  or (_29827_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_29828_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_29829_, _29828_, _29827_);
  or (_29830_, _29829_, _29826_);
  and (_29831_, \oc8051_golden_model_1.IRAM[11] [7], _32868_);
  and (_29832_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_29833_, _29832_, _29831_);
  nand (_29834_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_29835_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_29836_, _29835_, _29834_);
  or (_29837_, _29836_, _29833_);
  or (_29840_, _29837_, _29830_);
  or (_29841_, _29840_, _29823_);
  or (_29842_, _29841_, _29807_);
  or (_29843_, _29842_, _29772_);
  or (_29844_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand (_29845_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_29846_, _29845_, _29844_);
  nand (_29847_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_29848_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_29849_, _29848_, _29847_);
  or (_29851_, _29849_, _29846_);
  and (_29852_, \oc8051_golden_model_1.IRAM[12] [1], _32875_);
  and (_29853_, _04011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_29854_, _29853_, _29852_);
  and (_29855_, _03829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_29856_, \oc8051_golden_model_1.IRAM[12] [0], _32872_);
  or (_29857_, _29856_, _29855_);
  or (_29858_, _29857_, _29854_);
  or (_29859_, _29858_, _29851_);
  or (_29860_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_29862_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_29863_, _29862_, _29860_);
  nand (_29864_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_29865_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_29866_, _29865_, _29864_);
  or (_29867_, _29866_, _29863_);
  or (_29868_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand (_29869_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_29870_, _29869_, _29868_);
  or (_29871_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand (_29873_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_29874_, _29873_, _29871_);
  or (_29875_, _29874_, _29870_);
  or (_29876_, _29875_, _29867_);
  or (_29877_, _29876_, _29859_);
  or (_29878_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand (_29879_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_29880_, _29879_, _29878_);
  or (_29881_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand (_29882_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_29884_, _29882_, _29881_);
  or (_29885_, _29884_, _29880_);
  or (_29886_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand (_29887_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_29888_, _29887_, _29886_);
  nand (_29889_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_29890_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_29891_, _29890_, _29889_);
  or (_29892_, _29891_, _29888_);
  or (_29893_, _29892_, _29885_);
  and (_29895_, _05184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_29896_, \oc8051_golden_model_1.IRAM[13] [4], _32902_);
  or (_29897_, _29896_, _29895_);
  and (_29898_, _04886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_29899_, \oc8051_golden_model_1.IRAM[13] [5], _32905_);
  or (_29900_, _29899_, _29898_);
  or (_29901_, _29900_, _29897_);
  or (_29902_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand (_29903_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_29904_, _29903_, _29902_);
  nand (_29906_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_29907_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_29908_, _29907_, _29906_);
  or (_29909_, _29908_, _29904_);
  or (_29910_, _29909_, _29901_);
  or (_29911_, _29910_, _29893_);
  or (_29912_, _29911_, _29877_);
  or (_29913_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nand (_29914_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_29915_, _29914_, _29913_);
  or (_29917_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nand (_29918_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_29919_, _29918_, _29917_);
  or (_29920_, _29919_, _29915_);
  and (_29921_, \oc8051_golden_model_1.IRAM[14] [2], _32919_);
  and (_29922_, _04437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_29923_, _29922_, _29921_);
  nand (_29924_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_29925_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_29926_, _29925_, _29924_);
  or (_29928_, _29926_, _29923_);
  or (_29929_, _29928_, _29920_);
  and (_29930_, _05179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_29931_, \oc8051_golden_model_1.IRAM[14] [4], _32925_);
  or (_29932_, _29931_, _29930_);
  and (_29933_, \oc8051_golden_model_1.IRAM[14] [5], _32928_);
  and (_29934_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_29935_, _29934_, _29933_);
  or (_29936_, _29935_, _29932_);
  and (_29937_, _04616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_29939_, \oc8051_golden_model_1.IRAM[14] [7], _32574_);
  or (_29940_, _29939_, _29937_);
  nand (_29941_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_29942_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_29943_, _29942_, _29941_);
  or (_29944_, _29943_, _29940_);
  or (_29945_, _29944_, _29936_);
  or (_29946_, _29945_, _29929_);
  and (_29947_, _04006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_29948_, \oc8051_golden_model_1.IRAM[15] [1], _32939_);
  or (_29950_, _29948_, _29947_);
  and (_29951_, _03824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_29952_, \oc8051_golden_model_1.IRAM[15] [0], _32936_);
  or (_29953_, _29952_, _29951_);
  or (_29954_, _29953_, _29950_);
  and (_29955_, _04435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_29956_, \oc8051_golden_model_1.IRAM[15] [2], _32942_);
  or (_29957_, _29956_, _29955_);
  nand (_29958_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_29959_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_29961_, _29959_, _29958_);
  or (_29962_, _29961_, _29957_);
  or (_29963_, _29962_, _29954_);
  nand (_29964_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_29965_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_29966_, _29965_, _29964_);
  and (_29967_, \oc8051_golden_model_1.IRAM[15] [7], _32596_);
  and (_29968_, _04614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_29969_, _29968_, _29967_);
  or (_29970_, _29969_, _29966_);
  or (_29972_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_29973_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_29974_, _29973_, _29972_);
  or (_29975_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_29976_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_29977_, _29976_, _29975_);
  or (_29978_, _29977_, _29974_);
  or (_29979_, _29978_, _29970_);
  or (_29980_, _29979_, _29963_);
  or (_29981_, _29980_, _29946_);
  or (_29983_, _29981_, _29912_);
  or (_29984_, _29983_, _29843_);
  or (_29985_, _29984_, _29703_);
  and (property_invalid_iram, _29985_, _29151_);
  nand (_29986_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_29987_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_29988_, _29987_, _29986_);
  and (_29989_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_29990_, _16131_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_29991_, _29990_, _29989_);
  or (_29993_, _29991_, _29988_);
  nor (_29994_, _09380_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_29995_, _09380_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_29996_, _29995_, _29994_);
  and (_29997_, _16039_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_29998_, _16039_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_29999_, _29998_, _29997_);
  or (_30000_, _29999_, _29996_);
  or (_30001_, _30000_, _29993_);
  or (_30002_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_30004_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_30005_, _30004_, _30002_);
  or (_30006_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_30007_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_30008_, _30007_, _30006_);
  or (_30009_, _30008_, _30005_);
  and (_30010_, _08295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_30011_, _08295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_30012_, _30011_, _30010_);
  nand (_30013_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_30015_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_30016_, _30015_, _30013_);
  or (_30017_, _30016_, _30012_);
  or (_30018_, _30017_, _30009_);
  or (_30019_, _30018_, _30001_);
  and (property_invalid_dph, _30019_, _29151_);
  nand (_30020_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_30021_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_30022_, _30021_, _30020_);
  and (_30023_, _15494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_30025_, \oc8051_golden_model_1.DPL [2], _31356_);
  or (_30026_, _30025_, _30023_);
  or (_30027_, _30026_, _30022_);
  and (_30028_, \oc8051_golden_model_1.DPL [0], _31348_);
  and (_30029_, _15315_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_30030_, _30029_, _30028_);
  and (_30031_, _15402_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_30032_, \oc8051_golden_model_1.DPL [1], _31352_);
  or (_30033_, _30032_, _30031_);
  or (_30034_, _30033_, _30030_);
  or (_30036_, _30034_, _30027_);
  or (_30037_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_30038_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_30039_, _30038_, _30037_);
  or (_30040_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_30041_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_30042_, _30041_, _30040_);
  or (_30043_, _30042_, _30039_);
  and (_30044_, _08200_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_30045_, \oc8051_golden_model_1.DPL [7], _31127_);
  or (_30047_, _30045_, _30044_);
  nand (_30048_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_30049_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_30050_, _30049_, _30048_);
  or (_30051_, _30050_, _30047_);
  or (_30052_, _30051_, _30043_);
  or (_30053_, _30052_, _30036_);
  and (property_invalid_dpl, _30053_, _29151_);
  nand (_30054_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_30055_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_30057_, _30055_, _30054_);
  and (_30058_, _06951_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_30059_, \oc8051_golden_model_1.B [2], _30056_);
  or (_30060_, _30059_, _30058_);
  or (_30061_, _30060_, _30057_);
  and (_30062_, \oc8051_golden_model_1.B [0], _28772_);
  and (_30063_, _06798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_30064_, _30063_, _30062_);
  and (_30065_, _06793_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_30066_, \oc8051_golden_model_1.B [1], _29412_);
  or (_30068_, _30066_, _30065_);
  or (_30069_, _30068_, _30064_);
  or (_30070_, _30069_, _30061_);
  or (_30071_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_30072_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_30073_, _30072_, _30071_);
  or (_30074_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_30075_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_30076_, _30075_, _30074_);
  or (_30077_, _30076_, _30073_);
  and (_30079_, _06211_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_30080_, \oc8051_golden_model_1.B [7], _27722_);
  or (_30081_, _30080_, _30079_);
  nand (_30082_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_30083_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_30084_, _30083_, _30082_);
  or (_30085_, _30084_, _30081_);
  or (_30086_, _30085_, _30077_);
  or (_30087_, _30086_, _30070_);
  and (property_invalid_b_reg, _30087_, _29151_);
  nand (_30089_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_30090_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_30091_, _30090_, _30089_);
  and (_30092_, _06964_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_30093_, _06964_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_30094_, _30093_, _30092_);
  or (_30095_, _30094_, _30091_);
  nor (_30096_, _02543_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_30097_, _02543_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_30098_, _30097_, _30096_);
  and (_30100_, _02696_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_30101_, _02696_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_30102_, _30101_, _30100_);
  or (_30103_, _30102_, _30098_);
  or (_30104_, _30103_, _30095_);
  or (_30105_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_30106_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_30107_, _30106_, _30105_);
  or (_30108_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_30109_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_30111_, _30109_, _30108_);
  or (_30112_, _30111_, _30107_);
  and (_30113_, _06807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_30114_, _06807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_30115_, _30114_, _30113_);
  nand (_30116_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_30117_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_30118_, _30117_, _30116_);
  or (_30119_, _30118_, _30115_);
  or (_30120_, _30119_, _30112_);
  or (_30122_, _30120_, _30104_);
  and (property_invalid_acc, _30122_, _29151_);
  and (_30123_, _20271_, _35249_);
  nor (_30124_, _20271_, _35249_);
  or (_30125_, _30124_, _30123_);
  nor (_30126_, _20627_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_30127_, _20627_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_30128_, _30127_, _30126_);
  or (_30129_, _30128_, _30125_);
  and (_30130_, _22087_, _35268_);
  nor (_30132_, _22087_, _35268_);
  nor (_30133_, _20986_, _35256_);
  and (_30134_, _21732_, _35264_);
  and (_30135_, _20986_, _35256_);
  or (_30136_, _30135_, _30134_);
  or (_30137_, _30136_, _30133_);
  and (_30138_, _22454_, _35272_);
  and (_30139_, _21349_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_30140_, _21349_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_30141_, _24699_, _31065_);
  nand (_30143_, _24699_, _31065_);
  and (_30144_, _30143_, _30141_);
  and (_30145_, _24070_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_30146_, _24070_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_30147_, _23439_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_30148_, _23439_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_30149_, _30148_, _30147_);
  nand (_30150_, _22783_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_30151_, _22783_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_30152_, _30151_, _30150_);
  nand (_30153_, _23758_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_30154_, _23758_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_30155_, _30154_, _30153_);
  nor (_30156_, _19873_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_30157_, _19873_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_30158_, _30157_, _30156_);
  and (_30159_, _24388_, _31034_);
  nor (_30160_, _24388_, _31034_);
  or (_30161_, _30160_, _30159_);
  or (_30162_, _30161_, _30158_);
  or (_30165_, _30162_, _30155_);
  nor (_30166_, _09769_, _31070_);
  and (_30167_, _09769_, _31070_);
  or (_30168_, _30167_, _30166_);
  or (_30169_, _30168_, _30165_);
  or (_30170_, _30169_, _30152_);
  or (_30171_, _30170_, _30149_);
  or (_30172_, _30171_, _30146_);
  or (_30173_, _30172_, _30145_);
  or (_30174_, _30173_, _30144_);
  nor (_30176_, _23113_, _31048_);
  and (_30177_, _23113_, _31048_);
  or (_30178_, _30177_, _30176_);
  or (_30179_, _30178_, _30174_);
  or (_30180_, _30179_, _30140_);
  or (_30181_, _30180_, _30139_);
  or (_30182_, _30181_, _30138_);
  nor (_30183_, _22454_, _35272_);
  nor (_30184_, _21732_, _35264_);
  or (_30185_, _30184_, _30183_);
  or (_30187_, _30185_, _30182_);
  or (_30188_, _30187_, _30137_);
  or (_30189_, _30188_, _30132_);
  or (_30190_, _30189_, _30130_);
  or (_30191_, _30190_, _30129_);
  and (property_invalid_pc, _30191_, _28632_);
  buf (_35798_, _35796_);
  buf (_35812_, _35796_);
  buf (_35814_, _35796_);
  buf (_35816_, _35796_);
  buf (_35818_, _35796_);
  buf (_35820_, _35796_);
  buf (_35822_, _35796_);
  buf (_35824_, _35796_);
  buf (_35826_, _35796_);
  buf (_35800_, _35796_);
  buf (_35802_, _35796_);
  buf (_35804_, _35796_);
  buf (_35806_, _35796_);
  buf (_35808_, _35796_);
  buf (_35810_, _35796_);
  buf (_36006_[7], _35984_[7]);
  buf (_36007_[7], _35985_[7]);
  buf (_36018_[7], _35984_[7]);
  buf (_36019_[7], _35985_[7]);
  buf (_36006_[0], _35984_[0]);
  buf (_36006_[1], _35984_[1]);
  buf (_36006_[2], _35984_[2]);
  buf (_36006_[3], _35984_[3]);
  buf (_36006_[4], _35984_[4]);
  buf (_36006_[5], _35984_[5]);
  buf (_36006_[6], _35984_[6]);
  buf (_36007_[0], _35985_[0]);
  buf (_36007_[1], _35985_[1]);
  buf (_36007_[2], _35985_[2]);
  buf (_36007_[3], _35985_[3]);
  buf (_36007_[4], _35985_[4]);
  buf (_36007_[5], _35985_[5]);
  buf (_36007_[6], _35985_[6]);
  buf (_36018_[0], _35984_[0]);
  buf (_36018_[1], _35984_[1]);
  buf (_36018_[2], _35984_[2]);
  buf (_36018_[3], _35984_[3]);
  buf (_36018_[4], _35984_[4]);
  buf (_36018_[5], _35984_[5]);
  buf (_36018_[6], _35984_[6]);
  buf (_36019_[0], _35985_[0]);
  buf (_36019_[1], _35985_[1]);
  buf (_36019_[2], _35985_[2]);
  buf (_36019_[3], _35985_[3]);
  buf (_36019_[4], _35985_[4]);
  buf (_36019_[5], _35985_[5]);
  buf (_36019_[6], _35985_[6]);
  buf (_36138_, _35999_);
  buf (_36038_, _35999_);
  dff (xram_data_in_reg[0], _00008_[0]);
  dff (xram_data_in_reg[1], _00008_[1]);
  dff (xram_data_in_reg[2], _00008_[2]);
  dff (xram_data_in_reg[3], _00008_[3]);
  dff (xram_data_in_reg[4], _00008_[4]);
  dff (xram_data_in_reg[5], _00008_[5]);
  dff (xram_data_in_reg[6], _00008_[6]);
  dff (xram_data_in_reg[7], _00008_[7]);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (property_invalid_psw_1_r, _00006_);
  dff (property_invalid_sp_1_r, _00007_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _35795_[0]);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _35795_[1]);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _35795_[2]);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _35795_[3]);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _35795_[4]);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _35795_[5]);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _35795_[6]);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _35795_[7]);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _35796_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _35797_[0]);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _35797_[1]);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _35797_[2]);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _35797_[3]);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _35797_[4]);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _35797_[5]);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _35797_[6]);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _35797_[7]);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _35798_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _35799_[0]);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _35799_[1]);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _35799_[2]);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _35799_[3]);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _35799_[4]);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _35799_[5]);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _35799_[6]);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _35799_[7]);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _35800_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _35801_[0]);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _35801_[1]);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _35801_[2]);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _35801_[3]);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _35801_[4]);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _35801_[5]);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _35801_[6]);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _35801_[7]);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _35802_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _35803_[0]);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _35803_[1]);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _35803_[2]);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _35803_[3]);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _35803_[4]);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _35803_[5]);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _35803_[6]);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _35803_[7]);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _35804_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _35805_[0]);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _35805_[1]);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _35805_[2]);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _35805_[3]);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _35805_[4]);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _35805_[5]);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _35805_[6]);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _35805_[7]);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _35806_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _35807_[0]);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _35807_[1]);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _35807_[2]);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _35807_[3]);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _35807_[4]);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _35807_[5]);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _35807_[6]);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _35807_[7]);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _35808_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _35809_[0]);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _35809_[1]);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _35809_[2]);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _35809_[3]);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _35809_[4]);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _35809_[5]);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _35809_[6]);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _35809_[7]);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _35810_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _35811_[0]);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _35811_[1]);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _35811_[2]);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _35811_[3]);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _35811_[4]);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _35811_[5]);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _35811_[6]);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _35811_[7]);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _35812_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _35813_[0]);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _35813_[1]);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _35813_[2]);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _35813_[3]);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _35813_[4]);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _35813_[5]);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _35813_[6]);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _35813_[7]);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _35814_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _35815_[0]);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _35815_[1]);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _35815_[2]);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _35815_[3]);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _35815_[4]);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _35815_[5]);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _35815_[6]);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _35815_[7]);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _35816_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _35817_[0]);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _35817_[1]);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _35817_[2]);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _35817_[3]);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _35817_[4]);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _35817_[5]);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _35817_[6]);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _35817_[7]);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _35818_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _35819_[0]);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _35819_[1]);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _35819_[2]);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _35819_[3]);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _35819_[4]);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _35819_[5]);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _35819_[6]);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _35819_[7]);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _35820_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _35821_[0]);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _35821_[1]);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _35821_[2]);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _35821_[3]);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _35821_[4]);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _35821_[5]);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _35821_[6]);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _35821_[7]);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _35822_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _35823_[0]);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _35823_[1]);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _35823_[2]);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _35823_[3]);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _35823_[4]);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _35823_[5]);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _35823_[6]);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _35823_[7]);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _35824_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _35825_[0]);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _35825_[1]);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _35825_[2]);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _35825_[3]);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _35825_[4]);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _35825_[5]);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _35825_[6]);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _35825_[7]);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _35826_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _35903_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _35904_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _35905_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _35906_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _35907_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _35908_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _35909_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _35910_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _35895_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _35896_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _35897_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _35898_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _35899_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _35900_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _35901_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _35902_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _35887_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _35888_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _35889_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _35890_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _35891_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _35892_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _35893_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _35894_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _35879_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _35880_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _35881_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _35882_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _35883_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _35884_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _35885_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _35886_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _35871_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _35872_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _35873_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _35874_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _35875_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _35876_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _35877_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _35878_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _35863_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _35864_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _35865_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _35866_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _35867_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _35868_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _35869_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _35870_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _35975_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _35976_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _35977_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _35978_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _35979_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _35980_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _35981_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _35982_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _35967_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _35968_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _35969_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _35970_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _35971_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _35972_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _35973_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _35974_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _35959_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _35960_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _35961_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _35962_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _35963_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _35964_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _35965_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _35966_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _35951_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _35952_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _35953_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _35954_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _35955_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _35956_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _35957_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _35958_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _35943_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _35944_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _35945_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _35946_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _35947_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _35948_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _35949_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _35950_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _35935_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _35936_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _35937_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _35938_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _35939_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _35940_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _35941_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _35942_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _35927_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _35928_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _35929_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _35930_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _35931_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _35932_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _35933_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _35934_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _35919_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _35920_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _35921_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _35922_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _35923_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _35924_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _35925_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _35926_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _35911_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _35912_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _35913_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _35914_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _35915_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _35916_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _35917_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _35918_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _35855_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _35856_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _35857_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _35858_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _35859_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _35860_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _35861_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _35862_);
  dff (\oc8051_golden_model_1.B [0], _35828_[0]);
  dff (\oc8051_golden_model_1.B [1], _35828_[1]);
  dff (\oc8051_golden_model_1.B [2], _35828_[2]);
  dff (\oc8051_golden_model_1.B [3], _35828_[3]);
  dff (\oc8051_golden_model_1.B [4], _35828_[4]);
  dff (\oc8051_golden_model_1.B [5], _35828_[5]);
  dff (\oc8051_golden_model_1.B [6], _35828_[6]);
  dff (\oc8051_golden_model_1.B [7], _35828_[7]);
  dff (\oc8051_golden_model_1.ACC [0], _35827_[0]);
  dff (\oc8051_golden_model_1.ACC [1], _35827_[1]);
  dff (\oc8051_golden_model_1.ACC [2], _35827_[2]);
  dff (\oc8051_golden_model_1.ACC [3], _35827_[3]);
  dff (\oc8051_golden_model_1.ACC [4], _35827_[4]);
  dff (\oc8051_golden_model_1.ACC [5], _35827_[5]);
  dff (\oc8051_golden_model_1.ACC [6], _35827_[6]);
  dff (\oc8051_golden_model_1.ACC [7], _35827_[7]);
  dff (\oc8051_golden_model_1.DPL [0], _35830_[0]);
  dff (\oc8051_golden_model_1.DPL [1], _35830_[1]);
  dff (\oc8051_golden_model_1.DPL [2], _35830_[2]);
  dff (\oc8051_golden_model_1.DPL [3], _35830_[3]);
  dff (\oc8051_golden_model_1.DPL [4], _35830_[4]);
  dff (\oc8051_golden_model_1.DPL [5], _35830_[5]);
  dff (\oc8051_golden_model_1.DPL [6], _35830_[6]);
  dff (\oc8051_golden_model_1.DPL [7], _35830_[7]);
  dff (\oc8051_golden_model_1.DPH [0], _35829_[0]);
  dff (\oc8051_golden_model_1.DPH [1], _35829_[1]);
  dff (\oc8051_golden_model_1.DPH [2], _35829_[2]);
  dff (\oc8051_golden_model_1.DPH [3], _35829_[3]);
  dff (\oc8051_golden_model_1.DPH [4], _35829_[4]);
  dff (\oc8051_golden_model_1.DPH [5], _35829_[5]);
  dff (\oc8051_golden_model_1.DPH [6], _35829_[6]);
  dff (\oc8051_golden_model_1.DPH [7], _35829_[7]);
  dff (\oc8051_golden_model_1.IE [0], _35831_[0]);
  dff (\oc8051_golden_model_1.IE [1], _35831_[1]);
  dff (\oc8051_golden_model_1.IE [2], _35831_[2]);
  dff (\oc8051_golden_model_1.IE [3], _35831_[3]);
  dff (\oc8051_golden_model_1.IE [4], _35831_[4]);
  dff (\oc8051_golden_model_1.IE [5], _35831_[5]);
  dff (\oc8051_golden_model_1.IE [6], _35831_[6]);
  dff (\oc8051_golden_model_1.IE [7], _35831_[7]);
  dff (\oc8051_golden_model_1.IP [0], _35832_[0]);
  dff (\oc8051_golden_model_1.IP [1], _35832_[1]);
  dff (\oc8051_golden_model_1.IP [2], _35832_[2]);
  dff (\oc8051_golden_model_1.IP [3], _35832_[3]);
  dff (\oc8051_golden_model_1.IP [4], _35832_[4]);
  dff (\oc8051_golden_model_1.IP [5], _35832_[5]);
  dff (\oc8051_golden_model_1.IP [6], _35832_[6]);
  dff (\oc8051_golden_model_1.IP [7], _35832_[7]);
  dff (\oc8051_golden_model_1.P0 [0], _35834_[0]);
  dff (\oc8051_golden_model_1.P0 [1], _35834_[1]);
  dff (\oc8051_golden_model_1.P0 [2], _35834_[2]);
  dff (\oc8051_golden_model_1.P0 [3], _35834_[3]);
  dff (\oc8051_golden_model_1.P0 [4], _35834_[4]);
  dff (\oc8051_golden_model_1.P0 [5], _35834_[5]);
  dff (\oc8051_golden_model_1.P0 [6], _35834_[6]);
  dff (\oc8051_golden_model_1.P0 [7], _35834_[7]);
  dff (\oc8051_golden_model_1.P1 [0], _35836_[0]);
  dff (\oc8051_golden_model_1.P1 [1], _35836_[1]);
  dff (\oc8051_golden_model_1.P1 [2], _35836_[2]);
  dff (\oc8051_golden_model_1.P1 [3], _35836_[3]);
  dff (\oc8051_golden_model_1.P1 [4], _35836_[4]);
  dff (\oc8051_golden_model_1.P1 [5], _35836_[5]);
  dff (\oc8051_golden_model_1.P1 [6], _35836_[6]);
  dff (\oc8051_golden_model_1.P1 [7], _35836_[7]);
  dff (\oc8051_golden_model_1.P2 [0], _35838_[0]);
  dff (\oc8051_golden_model_1.P2 [1], _35838_[1]);
  dff (\oc8051_golden_model_1.P2 [2], _35838_[2]);
  dff (\oc8051_golden_model_1.P2 [3], _35838_[3]);
  dff (\oc8051_golden_model_1.P2 [4], _35838_[4]);
  dff (\oc8051_golden_model_1.P2 [5], _35838_[5]);
  dff (\oc8051_golden_model_1.P2 [6], _35838_[6]);
  dff (\oc8051_golden_model_1.P2 [7], _35838_[7]);
  dff (\oc8051_golden_model_1.P3 [0], _35840_[0]);
  dff (\oc8051_golden_model_1.P3 [1], _35840_[1]);
  dff (\oc8051_golden_model_1.P3 [2], _35840_[2]);
  dff (\oc8051_golden_model_1.P3 [3], _35840_[3]);
  dff (\oc8051_golden_model_1.P3 [4], _35840_[4]);
  dff (\oc8051_golden_model_1.P3 [5], _35840_[5]);
  dff (\oc8051_golden_model_1.P3 [6], _35840_[6]);
  dff (\oc8051_golden_model_1.P3 [7], _35840_[7]);
  dff (\oc8051_golden_model_1.PC [0], _35842_[0]);
  dff (\oc8051_golden_model_1.PC [1], _35842_[1]);
  dff (\oc8051_golden_model_1.PC [2], _35842_[2]);
  dff (\oc8051_golden_model_1.PC [3], _35842_[3]);
  dff (\oc8051_golden_model_1.PC [4], _35842_[4]);
  dff (\oc8051_golden_model_1.PC [5], _35842_[5]);
  dff (\oc8051_golden_model_1.PC [6], _35842_[6]);
  dff (\oc8051_golden_model_1.PC [7], _35842_[7]);
  dff (\oc8051_golden_model_1.PC [8], _35842_[8]);
  dff (\oc8051_golden_model_1.PC [9], _35842_[9]);
  dff (\oc8051_golden_model_1.PC [10], _35842_[10]);
  dff (\oc8051_golden_model_1.PC [11], _35842_[11]);
  dff (\oc8051_golden_model_1.PC [12], _35842_[12]);
  dff (\oc8051_golden_model_1.PC [13], _35842_[13]);
  dff (\oc8051_golden_model_1.PC [14], _35842_[14]);
  dff (\oc8051_golden_model_1.PC [15], _35842_[15]);
  dff (\oc8051_golden_model_1.PSW [0], _35843_[0]);
  dff (\oc8051_golden_model_1.PSW [1], _35843_[1]);
  dff (\oc8051_golden_model_1.PSW [2], _35843_[2]);
  dff (\oc8051_golden_model_1.PSW [3], _35843_[3]);
  dff (\oc8051_golden_model_1.PSW [4], _35843_[4]);
  dff (\oc8051_golden_model_1.PSW [5], _35843_[5]);
  dff (\oc8051_golden_model_1.PSW [6], _35843_[6]);
  dff (\oc8051_golden_model_1.PSW [7], _35843_[7]);
  dff (\oc8051_golden_model_1.PCON [0], _35841_[0]);
  dff (\oc8051_golden_model_1.PCON [1], _35841_[1]);
  dff (\oc8051_golden_model_1.PCON [2], _35841_[2]);
  dff (\oc8051_golden_model_1.PCON [3], _35841_[3]);
  dff (\oc8051_golden_model_1.PCON [4], _35841_[4]);
  dff (\oc8051_golden_model_1.PCON [5], _35841_[5]);
  dff (\oc8051_golden_model_1.PCON [6], _35841_[6]);
  dff (\oc8051_golden_model_1.PCON [7], _35841_[7]);
  dff (\oc8051_golden_model_1.SBUF [0], _35844_[0]);
  dff (\oc8051_golden_model_1.SBUF [1], _35844_[1]);
  dff (\oc8051_golden_model_1.SBUF [2], _35844_[2]);
  dff (\oc8051_golden_model_1.SBUF [3], _35844_[3]);
  dff (\oc8051_golden_model_1.SBUF [4], _35844_[4]);
  dff (\oc8051_golden_model_1.SBUF [5], _35844_[5]);
  dff (\oc8051_golden_model_1.SBUF [6], _35844_[6]);
  dff (\oc8051_golden_model_1.SBUF [7], _35844_[7]);
  dff (\oc8051_golden_model_1.SCON [0], _35845_[0]);
  dff (\oc8051_golden_model_1.SCON [1], _35845_[1]);
  dff (\oc8051_golden_model_1.SCON [2], _35845_[2]);
  dff (\oc8051_golden_model_1.SCON [3], _35845_[3]);
  dff (\oc8051_golden_model_1.SCON [4], _35845_[4]);
  dff (\oc8051_golden_model_1.SCON [5], _35845_[5]);
  dff (\oc8051_golden_model_1.SCON [6], _35845_[6]);
  dff (\oc8051_golden_model_1.SCON [7], _35845_[7]);
  dff (\oc8051_golden_model_1.SP [0], _35846_[0]);
  dff (\oc8051_golden_model_1.SP [1], _35846_[1]);
  dff (\oc8051_golden_model_1.SP [2], _35846_[2]);
  dff (\oc8051_golden_model_1.SP [3], _35846_[3]);
  dff (\oc8051_golden_model_1.SP [4], _35846_[4]);
  dff (\oc8051_golden_model_1.SP [5], _35846_[5]);
  dff (\oc8051_golden_model_1.SP [6], _35846_[6]);
  dff (\oc8051_golden_model_1.SP [7], _35846_[7]);
  dff (\oc8051_golden_model_1.TCON [0], _35847_[0]);
  dff (\oc8051_golden_model_1.TCON [1], _35847_[1]);
  dff (\oc8051_golden_model_1.TCON [2], _35847_[2]);
  dff (\oc8051_golden_model_1.TCON [3], _35847_[3]);
  dff (\oc8051_golden_model_1.TCON [4], _35847_[4]);
  dff (\oc8051_golden_model_1.TCON [5], _35847_[5]);
  dff (\oc8051_golden_model_1.TCON [6], _35847_[6]);
  dff (\oc8051_golden_model_1.TCON [7], _35847_[7]);
  dff (\oc8051_golden_model_1.TH0 [0], _35848_[0]);
  dff (\oc8051_golden_model_1.TH0 [1], _35848_[1]);
  dff (\oc8051_golden_model_1.TH0 [2], _35848_[2]);
  dff (\oc8051_golden_model_1.TH0 [3], _35848_[3]);
  dff (\oc8051_golden_model_1.TH0 [4], _35848_[4]);
  dff (\oc8051_golden_model_1.TH0 [5], _35848_[5]);
  dff (\oc8051_golden_model_1.TH0 [6], _35848_[6]);
  dff (\oc8051_golden_model_1.TH0 [7], _35848_[7]);
  dff (\oc8051_golden_model_1.TH1 [0], _35849_[0]);
  dff (\oc8051_golden_model_1.TH1 [1], _35849_[1]);
  dff (\oc8051_golden_model_1.TH1 [2], _35849_[2]);
  dff (\oc8051_golden_model_1.TH1 [3], _35849_[3]);
  dff (\oc8051_golden_model_1.TH1 [4], _35849_[4]);
  dff (\oc8051_golden_model_1.TH1 [5], _35849_[5]);
  dff (\oc8051_golden_model_1.TH1 [6], _35849_[6]);
  dff (\oc8051_golden_model_1.TH1 [7], _35849_[7]);
  dff (\oc8051_golden_model_1.TL0 [0], _35850_[0]);
  dff (\oc8051_golden_model_1.TL0 [1], _35850_[1]);
  dff (\oc8051_golden_model_1.TL0 [2], _35850_[2]);
  dff (\oc8051_golden_model_1.TL0 [3], _35850_[3]);
  dff (\oc8051_golden_model_1.TL0 [4], _35850_[4]);
  dff (\oc8051_golden_model_1.TL0 [5], _35850_[5]);
  dff (\oc8051_golden_model_1.TL0 [6], _35850_[6]);
  dff (\oc8051_golden_model_1.TL0 [7], _35850_[7]);
  dff (\oc8051_golden_model_1.TL1 [0], _35851_[0]);
  dff (\oc8051_golden_model_1.TL1 [1], _35851_[1]);
  dff (\oc8051_golden_model_1.TL1 [2], _35851_[2]);
  dff (\oc8051_golden_model_1.TL1 [3], _35851_[3]);
  dff (\oc8051_golden_model_1.TL1 [4], _35851_[4]);
  dff (\oc8051_golden_model_1.TL1 [5], _35851_[5]);
  dff (\oc8051_golden_model_1.TL1 [6], _35851_[6]);
  dff (\oc8051_golden_model_1.TL1 [7], _35851_[7]);
  dff (\oc8051_golden_model_1.TMOD [0], _35852_[0]);
  dff (\oc8051_golden_model_1.TMOD [1], _35852_[1]);
  dff (\oc8051_golden_model_1.TMOD [2], _35852_[2]);
  dff (\oc8051_golden_model_1.TMOD [3], _35852_[3]);
  dff (\oc8051_golden_model_1.TMOD [4], _35852_[4]);
  dff (\oc8051_golden_model_1.TMOD [5], _35852_[5]);
  dff (\oc8051_golden_model_1.TMOD [6], _35852_[6]);
  dff (\oc8051_golden_model_1.TMOD [7], _35852_[7]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [0], _35854_[0]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [1], _35854_[1]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [2], _35854_[2]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [3], _35854_[3]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [4], _35854_[4]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [5], _35854_[5]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [6], _35854_[6]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [7], _35854_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [0], _35853_[0]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [1], _35853_[1]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [2], _35853_[2]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [3], _35853_[3]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [4], _35853_[4]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [5], _35853_[5]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [6], _35853_[6]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [7], _35853_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [8], _35853_[8]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [9], _35853_[9]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [10], _35853_[10]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [11], _35853_[11]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [12], _35853_[12]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [13], _35853_[13]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [14], _35853_[14]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [15], _35853_[15]);
  dff (\oc8051_golden_model_1.P0INREG [0], _35833_[0]);
  dff (\oc8051_golden_model_1.P0INREG [1], _35833_[1]);
  dff (\oc8051_golden_model_1.P0INREG [2], _35833_[2]);
  dff (\oc8051_golden_model_1.P0INREG [3], _35833_[3]);
  dff (\oc8051_golden_model_1.P0INREG [4], _35833_[4]);
  dff (\oc8051_golden_model_1.P0INREG [5], _35833_[5]);
  dff (\oc8051_golden_model_1.P0INREG [6], _35833_[6]);
  dff (\oc8051_golden_model_1.P0INREG [7], _35833_[7]);
  dff (\oc8051_golden_model_1.P1INREG [0], _35835_[0]);
  dff (\oc8051_golden_model_1.P1INREG [1], _35835_[1]);
  dff (\oc8051_golden_model_1.P1INREG [2], _35835_[2]);
  dff (\oc8051_golden_model_1.P1INREG [3], _35835_[3]);
  dff (\oc8051_golden_model_1.P1INREG [4], _35835_[4]);
  dff (\oc8051_golden_model_1.P1INREG [5], _35835_[5]);
  dff (\oc8051_golden_model_1.P1INREG [6], _35835_[6]);
  dff (\oc8051_golden_model_1.P1INREG [7], _35835_[7]);
  dff (\oc8051_golden_model_1.P2INREG [0], _35837_[0]);
  dff (\oc8051_golden_model_1.P2INREG [1], _35837_[1]);
  dff (\oc8051_golden_model_1.P2INREG [2], _35837_[2]);
  dff (\oc8051_golden_model_1.P2INREG [3], _35837_[3]);
  dff (\oc8051_golden_model_1.P2INREG [4], _35837_[4]);
  dff (\oc8051_golden_model_1.P2INREG [5], _35837_[5]);
  dff (\oc8051_golden_model_1.P2INREG [6], _35837_[6]);
  dff (\oc8051_golden_model_1.P2INREG [7], _35837_[7]);
  dff (\oc8051_golden_model_1.P3INREG [0], _35839_[0]);
  dff (\oc8051_golden_model_1.P3INREG [1], _35839_[1]);
  dff (\oc8051_golden_model_1.P3INREG [2], _35839_[2]);
  dff (\oc8051_golden_model_1.P3INREG [3], _35839_[3]);
  dff (\oc8051_golden_model_1.P3INREG [4], _35839_[4]);
  dff (\oc8051_golden_model_1.P3INREG [5], _35839_[5]);
  dff (\oc8051_golden_model_1.P3INREG [6], _35839_[6]);
  dff (\oc8051_golden_model_1.P3INREG [7], _35839_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02918_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02929_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02950_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02972_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02993_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00945_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03004_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00915_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03015_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03026_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03037_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03048_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03059_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03070_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03081_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00965_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02556_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _24509_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02757_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02961_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03172_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03373_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03574_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03775_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03976_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04177_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04278_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04379_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04480_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04581_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04682_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04783_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04884_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _26705_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _35983_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _35983_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _35983_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _35983_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _35983_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _35983_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _35983_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _35983_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _35984_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _35984_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _35984_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _35984_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _35984_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _35984_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _35984_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _35984_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _35985_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _35985_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _35985_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _35985_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _35985_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _35985_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _35985_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _35985_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _35990_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _35991_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _35991_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _35992_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _35992_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _35993_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _35993_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _35993_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _35994_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _35994_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _35994_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _35995_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _35995_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _35996_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _35996_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _35996_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _35996_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _35997_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _35997_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _35998_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _35986_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _35986_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _35986_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _35987_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _35987_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _35987_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _35988_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _35988_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _35989_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _35989_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _35989_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _35989_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _35989_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _35989_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _35989_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _35989_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _35999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _36000_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _36000_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _36000_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _36000_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _36000_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _36000_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _36000_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _36000_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _36000_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _36000_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _36000_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _36000_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _36000_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _36000_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _36000_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _36000_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _36001_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _36001_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _36001_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _36001_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _36001_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _36001_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _36001_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _36001_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _36001_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _36001_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _36001_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _36001_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _36001_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _36001_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _36001_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _36001_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _36025_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _36025_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _36025_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _36025_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _36025_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _36025_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _36025_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _36025_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _36025_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _36025_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _36025_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _36025_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _36025_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _36025_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _36025_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _36025_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _36025_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _36025_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _36025_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _36025_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _36025_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _36025_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _36025_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _36025_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _36025_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _36025_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _36025_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _36025_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _36025_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _36025_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _36025_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _36025_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _36002_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , _36003_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _36004_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _36004_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _36004_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _36004_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _36004_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _36005_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _36005_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _36005_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _36005_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _36005_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _36005_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _36005_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _36005_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _36006_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _36006_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _36006_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _36006_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _36006_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _36006_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _36006_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _36006_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _36007_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _36007_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _36007_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _36007_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _36007_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _36007_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _36007_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _36007_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _36008_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _36009_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _36010_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _36010_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _36010_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _36010_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _36010_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _36010_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _36010_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _36010_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _36011_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _36011_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _36011_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _36011_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _36011_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _36011_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _36011_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _36011_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _36011_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _36011_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _36011_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _36011_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _36011_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _36011_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _36011_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _36011_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _36012_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _36012_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _36012_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _36012_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _36012_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _36012_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _36012_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _36012_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _36012_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _36012_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _36012_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _36012_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _36012_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _36012_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _36012_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _36012_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _36013_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _36015_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _36014_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _36016_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _36016_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _36016_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _36016_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _36016_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _36016_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _36016_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _36016_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _36017_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _36017_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _36017_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _36018_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _36018_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _36018_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _36018_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _36018_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _36018_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _36018_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _36018_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _36019_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _36019_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _36019_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _36019_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _36019_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _36019_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _36019_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _36019_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _36020_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _36021_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _36021_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _36021_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _36021_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _36021_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _36021_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _36021_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _36021_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _36022_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _36023_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _36024_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _36024_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _36024_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _36024_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _36026_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _36026_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _36026_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _36026_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _36026_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _36026_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _36026_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _36026_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _36026_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _36026_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _36026_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _36026_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _36026_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _36026_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _36026_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _36026_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _36026_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _36026_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _36026_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _36026_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _36026_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _36026_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _36026_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _36026_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _36026_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _36026_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _36026_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _36026_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _36026_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _36026_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _36026_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _36026_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _36027_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _36027_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _36027_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _36027_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _36027_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _36027_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _36027_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _36027_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _36028_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _36029_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _36030_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _36030_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _36030_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _36030_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _36030_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _36030_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _36030_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _36030_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _36030_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _36030_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _36030_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _36030_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _36030_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _36030_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _36030_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _36030_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _36031_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _36032_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _36033_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _36034_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _36034_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _36034_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _36034_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _36034_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _36034_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _36034_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _36034_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _36034_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _36034_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _36034_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _36034_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _36034_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _36034_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _36034_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _36034_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _36035_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _36036_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _36037_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _36037_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _36037_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _36037_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _36037_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _36037_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _36037_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _36037_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _36038_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _36039_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _36039_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _36039_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _33667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _33672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _33677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _33682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _33687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _33693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _33698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _33701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _36118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _36119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _36120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _36121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _36122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _36123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _36124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _36125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _33707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _33711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _33714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _33718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _33721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _33725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _33728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _33731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _36110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _36111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _36112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _36113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _36114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _36115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _36116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _36117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _36102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _36103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _36104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _36105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _36106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _36107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _36108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _36109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _36094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _36095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _36096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _36097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _36098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _36099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _36100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _36101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _33797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _36087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _36088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _36089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _36090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _36091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _36092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _36093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _33767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _33770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _33774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _33777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _33781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _33784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _33788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _33791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _33738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _33741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _33745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _33748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _33752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _33756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _33759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _33762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _36126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _36127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _36128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _36129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _36130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _36131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _36132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _36133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _36072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _36073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _36074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _36075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _36076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _36077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _36078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _36079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _36064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _36065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _36066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _36067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _36068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _36069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _36070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _36071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _36056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _36057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _36058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _36059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _36060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _36061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _36062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _36063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _36048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _36049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _36050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _36051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _36052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _36053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _36054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _36055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _36040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _36041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _36042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _36043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _36044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _36045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _36046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _36047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _36080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _36081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _36082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _36083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _36084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _36085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _36086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _33424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _36134_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _36134_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _36134_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _36134_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _36134_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _36134_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _36134_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _33414_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _36135_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _36136_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _36137_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _36137_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _36137_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _36137_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _36137_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _36137_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _36137_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _36137_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _36138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24099_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22201_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08838_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06574_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13391_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13402_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13413_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13446_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13468_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13490_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13501_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13511_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13522_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13533_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12477_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _33289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _33290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _33292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _33294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _33296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _33298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _33300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _30648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _33302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _33303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _33305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _33307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _33309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _33311_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _33313_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _30651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _33314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _33316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _33318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _33320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _33322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _33324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _33325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _30654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _33327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _33329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _33331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _33333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _33335_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _33336_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _33338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _30657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21361_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21373_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21397_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16434_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09422_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10566_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10577_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10588_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09443_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.dack_i , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [0], xram_data_in_reg[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [1], xram_data_in_reg[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [2], xram_data_in_reg[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [3], xram_data_in_reg[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [4], xram_data_in_reg[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [5], xram_data_in_reg[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [6], xram_data_in_reg[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [7], xram_data_in_reg[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.SBUF_next [0], \oc8051_golden_model_1.SBUF [0]);
  buf(\oc8051_golden_model_1.SBUF_next [1], \oc8051_golden_model_1.SBUF [1]);
  buf(\oc8051_golden_model_1.SBUF_next [2], \oc8051_golden_model_1.SBUF [2]);
  buf(\oc8051_golden_model_1.SBUF_next [3], \oc8051_golden_model_1.SBUF [3]);
  buf(\oc8051_golden_model_1.SBUF_next [4], \oc8051_golden_model_1.SBUF [4]);
  buf(\oc8051_golden_model_1.SBUF_next [5], \oc8051_golden_model_1.SBUF [5]);
  buf(\oc8051_golden_model_1.SBUF_next [6], \oc8051_golden_model_1.SBUF [6]);
  buf(\oc8051_golden_model_1.SBUF_next [7], \oc8051_golden_model_1.SBUF [7]);
  buf(\oc8051_golden_model_1.SCON_next [0], \oc8051_golden_model_1.SCON [0]);
  buf(\oc8051_golden_model_1.SCON_next [1], \oc8051_golden_model_1.SCON [1]);
  buf(\oc8051_golden_model_1.SCON_next [2], \oc8051_golden_model_1.SCON [2]);
  buf(\oc8051_golden_model_1.SCON_next [3], \oc8051_golden_model_1.SCON [3]);
  buf(\oc8051_golden_model_1.SCON_next [4], \oc8051_golden_model_1.SCON [4]);
  buf(\oc8051_golden_model_1.SCON_next [5], \oc8051_golden_model_1.SCON [5]);
  buf(\oc8051_golden_model_1.SCON_next [6], \oc8051_golden_model_1.SCON [6]);
  buf(\oc8051_golden_model_1.SCON_next [7], \oc8051_golden_model_1.SCON [7]);
  buf(\oc8051_golden_model_1.PCON_next [0], \oc8051_golden_model_1.PCON [0]);
  buf(\oc8051_golden_model_1.PCON_next [1], \oc8051_golden_model_1.PCON [1]);
  buf(\oc8051_golden_model_1.PCON_next [2], \oc8051_golden_model_1.PCON [2]);
  buf(\oc8051_golden_model_1.PCON_next [3], \oc8051_golden_model_1.PCON [3]);
  buf(\oc8051_golden_model_1.PCON_next [4], \oc8051_golden_model_1.PCON [4]);
  buf(\oc8051_golden_model_1.PCON_next [5], \oc8051_golden_model_1.PCON [5]);
  buf(\oc8051_golden_model_1.PCON_next [6], \oc8051_golden_model_1.PCON [6]);
  buf(\oc8051_golden_model_1.PCON_next [7], \oc8051_golden_model_1.PCON [7]);
  buf(\oc8051_golden_model_1.TCON_next [0], \oc8051_golden_model_1.TCON [0]);
  buf(\oc8051_golden_model_1.TCON_next [1], \oc8051_golden_model_1.TCON [1]);
  buf(\oc8051_golden_model_1.TCON_next [2], \oc8051_golden_model_1.TCON [2]);
  buf(\oc8051_golden_model_1.TCON_next [3], \oc8051_golden_model_1.TCON [3]);
  buf(\oc8051_golden_model_1.TCON_next [4], \oc8051_golden_model_1.TCON [4]);
  buf(\oc8051_golden_model_1.TCON_next [5], \oc8051_golden_model_1.TCON [5]);
  buf(\oc8051_golden_model_1.TCON_next [6], \oc8051_golden_model_1.TCON [6]);
  buf(\oc8051_golden_model_1.TCON_next [7], \oc8051_golden_model_1.TCON [7]);
  buf(\oc8051_golden_model_1.TL0_next [0], \oc8051_golden_model_1.TL0 [0]);
  buf(\oc8051_golden_model_1.TL0_next [1], \oc8051_golden_model_1.TL0 [1]);
  buf(\oc8051_golden_model_1.TL0_next [2], \oc8051_golden_model_1.TL0 [2]);
  buf(\oc8051_golden_model_1.TL0_next [3], \oc8051_golden_model_1.TL0 [3]);
  buf(\oc8051_golden_model_1.TL0_next [4], \oc8051_golden_model_1.TL0 [4]);
  buf(\oc8051_golden_model_1.TL0_next [5], \oc8051_golden_model_1.TL0 [5]);
  buf(\oc8051_golden_model_1.TL0_next [6], \oc8051_golden_model_1.TL0 [6]);
  buf(\oc8051_golden_model_1.TL0_next [7], \oc8051_golden_model_1.TL0 [7]);
  buf(\oc8051_golden_model_1.TL1_next [0], \oc8051_golden_model_1.TL1 [0]);
  buf(\oc8051_golden_model_1.TL1_next [1], \oc8051_golden_model_1.TL1 [1]);
  buf(\oc8051_golden_model_1.TL1_next [2], \oc8051_golden_model_1.TL1 [2]);
  buf(\oc8051_golden_model_1.TL1_next [3], \oc8051_golden_model_1.TL1 [3]);
  buf(\oc8051_golden_model_1.TL1_next [4], \oc8051_golden_model_1.TL1 [4]);
  buf(\oc8051_golden_model_1.TL1_next [5], \oc8051_golden_model_1.TL1 [5]);
  buf(\oc8051_golden_model_1.TL1_next [6], \oc8051_golden_model_1.TL1 [6]);
  buf(\oc8051_golden_model_1.TL1_next [7], \oc8051_golden_model_1.TL1 [7]);
  buf(\oc8051_golden_model_1.TH0_next [0], \oc8051_golden_model_1.TH0 [0]);
  buf(\oc8051_golden_model_1.TH0_next [1], \oc8051_golden_model_1.TH0 [1]);
  buf(\oc8051_golden_model_1.TH0_next [2], \oc8051_golden_model_1.TH0 [2]);
  buf(\oc8051_golden_model_1.TH0_next [3], \oc8051_golden_model_1.TH0 [3]);
  buf(\oc8051_golden_model_1.TH0_next [4], \oc8051_golden_model_1.TH0 [4]);
  buf(\oc8051_golden_model_1.TH0_next [5], \oc8051_golden_model_1.TH0 [5]);
  buf(\oc8051_golden_model_1.TH0_next [6], \oc8051_golden_model_1.TH0 [6]);
  buf(\oc8051_golden_model_1.TH0_next [7], \oc8051_golden_model_1.TH0 [7]);
  buf(\oc8051_golden_model_1.TH1_next [0], \oc8051_golden_model_1.TH1 [0]);
  buf(\oc8051_golden_model_1.TH1_next [1], \oc8051_golden_model_1.TH1 [1]);
  buf(\oc8051_golden_model_1.TH1_next [2], \oc8051_golden_model_1.TH1 [2]);
  buf(\oc8051_golden_model_1.TH1_next [3], \oc8051_golden_model_1.TH1 [3]);
  buf(\oc8051_golden_model_1.TH1_next [4], \oc8051_golden_model_1.TH1 [4]);
  buf(\oc8051_golden_model_1.TH1_next [5], \oc8051_golden_model_1.TH1 [5]);
  buf(\oc8051_golden_model_1.TH1_next [6], \oc8051_golden_model_1.TH1 [6]);
  buf(\oc8051_golden_model_1.TH1_next [7], \oc8051_golden_model_1.TH1 [7]);
  buf(\oc8051_golden_model_1.TMOD_next [0], \oc8051_golden_model_1.TMOD [0]);
  buf(\oc8051_golden_model_1.TMOD_next [1], \oc8051_golden_model_1.TMOD [1]);
  buf(\oc8051_golden_model_1.TMOD_next [2], \oc8051_golden_model_1.TMOD [2]);
  buf(\oc8051_golden_model_1.TMOD_next [3], \oc8051_golden_model_1.TMOD [3]);
  buf(\oc8051_golden_model_1.TMOD_next [4], \oc8051_golden_model_1.TMOD [4]);
  buf(\oc8051_golden_model_1.TMOD_next [5], \oc8051_golden_model_1.TMOD [5]);
  buf(\oc8051_golden_model_1.TMOD_next [6], \oc8051_golden_model_1.TMOD [6]);
  buf(\oc8051_golden_model_1.TMOD_next [7], \oc8051_golden_model_1.TMOD [7]);
  buf(\oc8051_golden_model_1.IE_next [0], \oc8051_golden_model_1.IE [0]);
  buf(\oc8051_golden_model_1.IE_next [1], \oc8051_golden_model_1.IE [1]);
  buf(\oc8051_golden_model_1.IE_next [2], \oc8051_golden_model_1.IE [2]);
  buf(\oc8051_golden_model_1.IE_next [3], \oc8051_golden_model_1.IE [3]);
  buf(\oc8051_golden_model_1.IE_next [4], \oc8051_golden_model_1.IE [4]);
  buf(\oc8051_golden_model_1.IE_next [5], \oc8051_golden_model_1.IE [5]);
  buf(\oc8051_golden_model_1.IE_next [6], \oc8051_golden_model_1.IE [6]);
  buf(\oc8051_golden_model_1.IE_next [7], \oc8051_golden_model_1.IE [7]);
  buf(\oc8051_golden_model_1.IP_next [0], \oc8051_golden_model_1.IP [0]);
  buf(\oc8051_golden_model_1.IP_next [1], \oc8051_golden_model_1.IP [1]);
  buf(\oc8051_golden_model_1.IP_next [2], \oc8051_golden_model_1.IP [2]);
  buf(\oc8051_golden_model_1.IP_next [3], \oc8051_golden_model_1.IP [3]);
  buf(\oc8051_golden_model_1.IP_next [4], \oc8051_golden_model_1.IP [4]);
  buf(\oc8051_golden_model_1.IP_next [5], \oc8051_golden_model_1.IP [5]);
  buf(\oc8051_golden_model_1.IP_next [6], \oc8051_golden_model_1.IP [6]);
  buf(\oc8051_golden_model_1.IP_next [7], \oc8051_golden_model_1.IP [7]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [0], xram_data_in_reg[0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [1], xram_data_in_reg[1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [2], xram_data_in_reg[2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [3], xram_data_in_reg[3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [4], xram_data_in_reg[4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [5], xram_data_in_reg[5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [6], xram_data_in_reg[6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [7], xram_data_in_reg[7]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e0 [0], xram_data_in_reg[0]);
  buf(\oc8051_golden_model_1.ACC_e0 [1], xram_data_in_reg[1]);
  buf(\oc8051_golden_model_1.ACC_e0 [2], xram_data_in_reg[2]);
  buf(\oc8051_golden_model_1.ACC_e0 [3], xram_data_in_reg[3]);
  buf(\oc8051_golden_model_1.ACC_e0 [4], xram_data_in_reg[4]);
  buf(\oc8051_golden_model_1.ACC_e0 [5], xram_data_in_reg[5]);
  buf(\oc8051_golden_model_1.ACC_e0 [6], xram_data_in_reg[6]);
  buf(\oc8051_golden_model_1.ACC_e0 [7], xram_data_in_reg[7]);
  buf(\oc8051_golden_model_1.ACC_e2 [0], xram_data_in_reg[0]);
  buf(\oc8051_golden_model_1.ACC_e2 [1], xram_data_in_reg[1]);
  buf(\oc8051_golden_model_1.ACC_e2 [2], xram_data_in_reg[2]);
  buf(\oc8051_golden_model_1.ACC_e2 [3], xram_data_in_reg[3]);
  buf(\oc8051_golden_model_1.ACC_e2 [4], xram_data_in_reg[4]);
  buf(\oc8051_golden_model_1.ACC_e2 [5], xram_data_in_reg[5]);
  buf(\oc8051_golden_model_1.ACC_e2 [6], xram_data_in_reg[6]);
  buf(\oc8051_golden_model_1.ACC_e2 [7], xram_data_in_reg[7]);
  buf(\oc8051_golden_model_1.ACC_e3 [0], xram_data_in_reg[0]);
  buf(\oc8051_golden_model_1.ACC_e3 [1], xram_data_in_reg[1]);
  buf(\oc8051_golden_model_1.ACC_e3 [2], xram_data_in_reg[2]);
  buf(\oc8051_golden_model_1.ACC_e3 [3], xram_data_in_reg[3]);
  buf(\oc8051_golden_model_1.ACC_e3 [4], xram_data_in_reg[4]);
  buf(\oc8051_golden_model_1.ACC_e3 [5], xram_data_in_reg[5]);
  buf(\oc8051_golden_model_1.ACC_e3 [6], xram_data_in_reg[6]);
  buf(\oc8051_golden_model_1.ACC_e3 [7], xram_data_in_reg[7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1041 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1058 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1262 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1279 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1328 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1369 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1425 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1551 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1620 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1653 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1653 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1702 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1702 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1702 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1702 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1747 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1764 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1781 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1781 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1812 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1812 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1812 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1812 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1812 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1812 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1812 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1857 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1874 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1891 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1891 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n1984 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2001 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2018 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2018 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2116 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2302 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2332 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2362 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2362 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2428 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2537 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2664 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2686 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2686 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e0 [0], \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.PSW_e0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e2 [0], \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.PSW_e2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e2 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e3 [0], \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.PSW_e3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2722 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2723 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f2 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f2 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2740 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1002 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1002 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1002 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1002 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1002 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1002 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1002 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1004 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1005 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1006 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1007 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1008 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1018 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1018 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1018 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1018 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1018 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1018 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1018 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1018 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1025 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1025 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1025 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1025 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1025 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1025 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1025 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1025 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1027 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1028 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1029 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1030 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1040 , \oc8051_golden_model_1.n1041 [0]);
  buf(\oc8051_golden_model_1.n1041 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1041 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1041 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1041 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1041 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1041 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1041 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1057 , \oc8051_golden_model_1.n1058 [0]);
  buf(\oc8051_golden_model_1.n1058 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1058 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1058 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1058 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1058 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1058 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1058 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1139 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1139 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1139 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1139 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1141 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1143 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1144 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1144 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1145 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1146 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1147 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1148 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1148 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1148 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1149 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1149 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1149 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1195 , \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1239 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1239 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1239 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1239 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1239 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1239 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1239 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1239 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1239 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1240 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1240 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1240 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1240 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1240 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1240 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1240 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1241 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1242 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1242 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1242 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1243 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1244 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1244 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1245 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1245 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1245 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1245 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1245 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1245 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1245 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1245 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1246 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1247 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1248 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1249 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1251 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1252 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1253 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1254 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 , \oc8051_golden_model_1.n1262 [0]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1278 , \oc8051_golden_model_1.n1279 [0]);
  buf(\oc8051_golden_model_1.n1279 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1279 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1279 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1279 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1279 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1279 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1279 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1310 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1310 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1310 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1310 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1310 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n1310 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n1310 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n1310 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1310 [8], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1310 [9], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1310 [10], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1310 [11], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1310 [12], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n1310 [13], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n1310 [14], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n1310 [15], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1312 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1312 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1312 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1312 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1312 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1312 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1312 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1312 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1313 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1314 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1315 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1316 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1318 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1319 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1320 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1327 , \oc8051_golden_model_1.n1328 [0]);
  buf(\oc8051_golden_model_1.n1328 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1328 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1328 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1328 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1328 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1328 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1328 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1330 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1330 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1330 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1330 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1330 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1330 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1330 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1330 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1330 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1334 [8], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1335 , \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1336 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1336 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1336 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1336 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1337 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1337 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1337 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1337 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1337 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.n1352 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1352 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1352 [2], \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.n1352 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1352 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1352 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1352 [6], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1352 [7], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1353 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1353 [1], \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.n1353 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1353 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1353 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1353 [5], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1353 [6], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1369 [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1369 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1369 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1392 [8], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1393 , \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1398 [4], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1399 , \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1407 , \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.n1408 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1408 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1408 [2], \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.n1408 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1408 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1408 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1408 [6], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1408 [7], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1409 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1409 [1], \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.n1409 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1409 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1409 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1409 [5], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1409 [6], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1424 , \oc8051_golden_model_1.n1425 [0]);
  buf(\oc8051_golden_model_1.n1425 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1425 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1425 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1425 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1427 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1427 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1427 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1427 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1427 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n1427 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n1427 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n1427 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1427 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1429 [8], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1430 , \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1431 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1431 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1431 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1431 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1432 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1432 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1432 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1432 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1432 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1434 [4], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1435 , \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1436 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1436 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1436 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1436 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1436 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n1436 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n1436 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n1436 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1436 [8], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1443 , \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.n1444 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1444 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1444 [2], \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.n1444 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1444 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1444 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1444 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1444 [7], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1445 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1445 [1], \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.n1445 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1445 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1445 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1445 [5], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1445 [6], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1460 , \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.n1461 [0], \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.n1461 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1461 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1461 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1461 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1461 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1463 [8], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1464 , \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1471 , \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.n1472 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1472 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1472 [2], \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.n1472 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1472 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1472 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1472 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1472 [7], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1473 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1473 [1], \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.n1473 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1473 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1473 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1473 [5], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1473 [6], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1474 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1474 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1474 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1474 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1476 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1478 [8], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1479 , \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1480 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1480 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1480 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1480 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1480 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1482 [4], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1483 , \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1484 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1484 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1484 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1484 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1484 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n1484 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n1484 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n1484 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1484 [8], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1491 , \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1492 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1492 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1492 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1492 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1492 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1492 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1492 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1492 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1508 , \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1511 [4], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1513 [6], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1513 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1514 [1], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1514 [5], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1514 [6], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1515 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.n1515 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1515 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1515 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1518 , \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1525 , \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1526 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1527 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1527 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1527 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1527 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1527 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1527 [5], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1527 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1531 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1531 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1531 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1531 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1531 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1531 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1531 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1531 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1531 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1532 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1532 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1532 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1532 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1532 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1532 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1532 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1532 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1532 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1533 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1533 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1533 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1533 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1533 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1533 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1533 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1533 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1534 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1534 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1534 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1534 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1534 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1534 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1534 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1534 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1535 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1535 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1535 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1535 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1535 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1535 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1535 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1536 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1537 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1538 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1539 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1540 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1542 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1543 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1550 , \oc8051_golden_model_1.n1551 [0]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1551 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1552 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1552 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1555 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1557 [8], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1559 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1559 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1559 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1559 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1562 , \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1569 , \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1586 , \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1591 [8], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1592 , \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1594 [4], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1595 , \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1602 , \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.n1603 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1603 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1603 [2], \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.n1603 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1603 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1603 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1603 [6], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1603 [7], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1604 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1604 [1], \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.n1604 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1604 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1604 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1604 [5], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1604 [6], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1619 , \oc8051_golden_model_1.n1620 [0]);
  buf(\oc8051_golden_model_1.n1620 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1620 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1620 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1620 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1624 [8], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1625 , \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1627 [4], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1628 , \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1635 , \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.n1636 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1636 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1636 [2], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.n1636 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1636 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1636 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1636 [6], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1636 [7], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1637 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1637 [1], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.n1637 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1637 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1637 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1637 [5], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1637 [6], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1652 , \oc8051_golden_model_1.n1653 [0]);
  buf(\oc8051_golden_model_1.n1653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1657 [8], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1658 , \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1660 [4], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1668 , \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.n1669 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1669 [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.n1669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1669 [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1669 [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1670 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1670 [1], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.n1670 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1670 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1670 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1670 [5], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1670 [6], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.n1686 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1686 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1686 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1686 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1700 [1], \oc8051_golden_model_1.n1702 [1]);
  buf(\oc8051_golden_model_1.n1700 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1700 [3], \oc8051_golden_model_1.n1702 [3]);
  buf(\oc8051_golden_model_1.n1700 [4], \oc8051_golden_model_1.n1702 [4]);
  buf(\oc8051_golden_model_1.n1700 [5], \oc8051_golden_model_1.n1702 [5]);
  buf(\oc8051_golden_model_1.n1700 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1700 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1701 [0], \oc8051_golden_model_1.n1702 [1]);
  buf(\oc8051_golden_model_1.n1701 [1], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1701 [2], \oc8051_golden_model_1.n1702 [3]);
  buf(\oc8051_golden_model_1.n1701 [3], \oc8051_golden_model_1.n1702 [4]);
  buf(\oc8051_golden_model_1.n1701 [4], \oc8051_golden_model_1.n1702 [5]);
  buf(\oc8051_golden_model_1.n1701 [5], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1701 [6], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1702 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1746 , \oc8051_golden_model_1.n1747 [0]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1747 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1747 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1747 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1763 , \oc8051_golden_model_1.n1764 [0]);
  buf(\oc8051_golden_model_1.n1764 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1764 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1764 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1764 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1764 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1764 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1764 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1780 , \oc8051_golden_model_1.n1781 [0]);
  buf(\oc8051_golden_model_1.n1781 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1781 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1781 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1781 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1781 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1781 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1781 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1797 , \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.n1798 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1798 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1798 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1798 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1798 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1798 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1798 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1810 [1], \oc8051_golden_model_1.n1812 [1]);
  buf(\oc8051_golden_model_1.n1810 [2], \oc8051_golden_model_1.n1812 [2]);
  buf(\oc8051_golden_model_1.n1810 [3], \oc8051_golden_model_1.n1812 [3]);
  buf(\oc8051_golden_model_1.n1810 [4], \oc8051_golden_model_1.n1812 [4]);
  buf(\oc8051_golden_model_1.n1810 [5], \oc8051_golden_model_1.n1812 [5]);
  buf(\oc8051_golden_model_1.n1810 [6], \oc8051_golden_model_1.n1812 [6]);
  buf(\oc8051_golden_model_1.n1810 [7], \oc8051_golden_model_1.n1812 [7]);
  buf(\oc8051_golden_model_1.n1811 [0], \oc8051_golden_model_1.n1812 [1]);
  buf(\oc8051_golden_model_1.n1811 [1], \oc8051_golden_model_1.n1812 [2]);
  buf(\oc8051_golden_model_1.n1811 [2], \oc8051_golden_model_1.n1812 [3]);
  buf(\oc8051_golden_model_1.n1811 [3], \oc8051_golden_model_1.n1812 [4]);
  buf(\oc8051_golden_model_1.n1811 [4], \oc8051_golden_model_1.n1812 [5]);
  buf(\oc8051_golden_model_1.n1811 [5], \oc8051_golden_model_1.n1812 [6]);
  buf(\oc8051_golden_model_1.n1811 [6], \oc8051_golden_model_1.n1812 [7]);
  buf(\oc8051_golden_model_1.n1812 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1856 , \oc8051_golden_model_1.n1857 [0]);
  buf(\oc8051_golden_model_1.n1857 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1857 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1857 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1857 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1857 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1857 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1857 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1873 , \oc8051_golden_model_1.n1874 [0]);
  buf(\oc8051_golden_model_1.n1874 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1874 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1874 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1874 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1874 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1874 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1874 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1890 , \oc8051_golden_model_1.n1891 [0]);
  buf(\oc8051_golden_model_1.n1891 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1891 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1891 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1891 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1891 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1891 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1891 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1907 , \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.n1908 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1908 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1908 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1908 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1908 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1908 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1908 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1983 , \oc8051_golden_model_1.n1984 [0]);
  buf(\oc8051_golden_model_1.n1984 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1984 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1984 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1984 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1984 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1984 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1984 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2000 , \oc8051_golden_model_1.n2001 [0]);
  buf(\oc8051_golden_model_1.n2001 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2001 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2001 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2001 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2001 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2001 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2001 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2017 , \oc8051_golden_model_1.n2018 [0]);
  buf(\oc8051_golden_model_1.n2018 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2018 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2018 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2018 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2018 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2018 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2018 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2034 , \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.n2035 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2035 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2035 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2035 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2035 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2039 , \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.n2040 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2040 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2040 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2040 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2040 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2040 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2040 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2041 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2041 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2041 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2041 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2041 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2041 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2041 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2041 [7], \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.n2042 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2042 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2042 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2042 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2042 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2042 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2042 [6], \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.n2043 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2043 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2043 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2043 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2043 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2043 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2043 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2058 , \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.n2059 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2059 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2059 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2059 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2059 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2059 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2059 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2087 , \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.n2088 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2088 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2088 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2088 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2088 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2088 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2088 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2088 [7], \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.n2089 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2089 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2089 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2089 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2089 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2089 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2089 [6], \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.n2090 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2090 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2090 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2090 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2090 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2090 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2090 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2097 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2097 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2097 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2097 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2098 , \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.n2099 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2099 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2099 [2], \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.n2099 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2099 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2099 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2099 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2099 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2100 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2100 [1], \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.n2100 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2100 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2100 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2100 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2100 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2115 , \oc8051_golden_model_1.n2116 [0]);
  buf(\oc8051_golden_model_1.n2116 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2116 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2116 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2116 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2116 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2116 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2273 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2276 , \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.n2278 , \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.n2284 , \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.n2285 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2285 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2285 [2], \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.n2285 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2285 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2285 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2285 [6], \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.n2285 [7], \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.n2286 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2286 [1], \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.n2286 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2286 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2286 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2286 [5], \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.n2286 [6], \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.n2301 , \oc8051_golden_model_1.n2302 [0]);
  buf(\oc8051_golden_model_1.n2302 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2302 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2302 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2302 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2306 , \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.n2308 , \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.n2314 , \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.n2315 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2315 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2315 [2], \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.n2315 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2315 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2315 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2315 [6], \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.n2315 [7], \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.n2316 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2316 [1], \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.n2316 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2316 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2316 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2316 [5], \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.n2316 [6], \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.n2331 , \oc8051_golden_model_1.n2332 [0]);
  buf(\oc8051_golden_model_1.n2332 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2332 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2332 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2332 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2336 , \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.n2338 , \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.n2344 , \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.n2345 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2345 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2345 [2], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.n2345 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2345 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2345 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2345 [6], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.n2345 [7], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.n2346 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2346 [1], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.n2346 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2346 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2346 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2346 [5], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.n2346 [6], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.n2361 , \oc8051_golden_model_1.n2362 [0]);
  buf(\oc8051_golden_model_1.n2362 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2362 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2362 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2362 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2366 , \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.n2368 , \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.n2374 , \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.n2375 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2375 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2375 [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.n2375 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2375 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2375 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2375 [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.n2375 [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.n2376 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2376 [1], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.n2376 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2376 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2376 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2376 [5], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.n2376 [6], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.n2391 , \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.n2392 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2392 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2392 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2392 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2394 , \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.n2395 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2395 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2395 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2395 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2395 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2395 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2395 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2395 [7], \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.n2396 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2396 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2396 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2396 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2396 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2396 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2396 [6], \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.n2397 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2397 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2397 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2397 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2397 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2397 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2397 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2398 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2398 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2398 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2398 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2398 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2398 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2398 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2398 [7], \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.n2399 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2399 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2399 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2399 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2399 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2399 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2399 [6], \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.n2400 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2400 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2400 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2400 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2400 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2400 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2400 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2404 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2404 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2404 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2404 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2404 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2404 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2404 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2404 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2404 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2410 , \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.n2411 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2411 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2411 [2], \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.n2411 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2411 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2411 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2411 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2411 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2412 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2412 [1], \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.n2412 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2412 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2412 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2412 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2412 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2427 , \oc8051_golden_model_1.n2428 [0]);
  buf(\oc8051_golden_model_1.n2428 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2428 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2428 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2428 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2428 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2428 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2430 , \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.n2431 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2431 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2431 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2431 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2431 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2431 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2431 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2431 [7], \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.n2432 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2432 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2432 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2432 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2432 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2432 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2432 [6], \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.n2433 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2433 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2433 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2433 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2433 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2433 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2433 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2461 , \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.n2462 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2462 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2462 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2462 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2462 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2462 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2462 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2462 [7], \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.n2463 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2463 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2463 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2463 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2463 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2463 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2463 [6], \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.n2464 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2464 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2464 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2464 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2464 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2464 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2464 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.n2470 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2470 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2470 [7], \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.n2471 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2471 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2471 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2471 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2471 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2471 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2471 [6], \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.n2472 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2472 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2472 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2472 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2472 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2472 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2472 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2477 , \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2478 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2478 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2478 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2478 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2478 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2478 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2478 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2478 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2479 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2479 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2479 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2479 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2479 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2479 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2479 [6], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2480 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2480 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2480 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2480 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2480 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2480 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2480 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2485 , \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.n2486 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2486 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2486 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2486 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2486 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2486 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2486 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2486 [7], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.n2487 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2487 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2487 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2487 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2487 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2487 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2487 [6], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.n2488 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2488 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2488 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2488 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2488 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2488 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2488 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2493 , \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.n2494 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2494 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2494 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2494 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2494 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2494 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2494 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2494 [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.n2495 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2495 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2495 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2495 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2495 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2495 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2495 [6], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.n2496 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2496 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2496 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2496 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2496 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2496 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2496 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2517 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2517 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2517 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2517 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2517 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2517 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2517 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2517 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2518 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2518 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2518 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2518 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2518 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2518 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2518 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2519 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2519 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2519 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2519 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2519 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2519 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2519 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2519 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2520 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2520 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2520 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2520 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2521 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2521 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2521 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2521 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2521 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2521 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2521 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2521 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2522 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2523 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2524 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2525 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2526 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2527 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2528 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.n2537 [0]);
  buf(\oc8051_golden_model_1.n2537 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2537 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2537 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2537 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2537 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2537 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2537 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2546 [1], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.n2546 [2], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.n2546 [3], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.n2546 [4], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.n2546 [5], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.n2546 [6], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.n2546 [7], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.n2547 [0], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.n2547 [2], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.n2547 [6], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.n2562 , \oc8051_golden_model_1.n2723 [0]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.n2723 [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.n2564 , \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n2565 , \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n2566 , \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n2567 , \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n2568 , \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n2569 , \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n2570 , \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n2571 , \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2580 , \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n2581 , \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n2582 , \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n2583 , \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n2584 , \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n2585 , \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n2586 , \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n2587 , \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n2594 , \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.n2595 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2595 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2595 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2595 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2595 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2595 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2595 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2625 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2625 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2625 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2625 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2625 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2625 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2625 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2625 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2626 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2626 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2626 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2626 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2626 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2626 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2626 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2627 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2627 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2627 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2627 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2627 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2627 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2627 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2627 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2646 , \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.n2647 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2647 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2647 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2647 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2647 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2647 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2647 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2647 [7], \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.n2648 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2648 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2648 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2648 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2648 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2648 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2648 [6], \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.n2663 , \oc8051_golden_model_1.n2664 [0]);
  buf(\oc8051_golden_model_1.n2664 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2664 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2664 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2664 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2664 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2664 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2668 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n2670 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2670 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2670 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2670 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2671 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2672 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2673 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2674 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2685 , \oc8051_golden_model_1.n2686 [0]);
  buf(\oc8051_golden_model_1.n2686 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2686 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2686 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2686 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2686 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2686 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2686 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2690 , xram_data_in_reg[7]);
  buf(\oc8051_golden_model_1.n2691 , xram_data_in_reg[6]);
  buf(\oc8051_golden_model_1.n2692 , xram_data_in_reg[5]);
  buf(\oc8051_golden_model_1.n2693 , xram_data_in_reg[4]);
  buf(\oc8051_golden_model_1.n2694 , xram_data_in_reg[3]);
  buf(\oc8051_golden_model_1.n2695 , xram_data_in_reg[2]);
  buf(\oc8051_golden_model_1.n2696 , xram_data_in_reg[1]);
  buf(\oc8051_golden_model_1.n2697 , xram_data_in_reg[0]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.n2705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2705 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2705 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2705 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2706 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2721 , \oc8051_golden_model_1.n2722 [0]);
  buf(\oc8051_golden_model_1.n2722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2722 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2722 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2722 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2723 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2723 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2723 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2723 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2723 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2723 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2723 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2739 , \oc8051_golden_model_1.n2740 [0]);
  buf(\oc8051_golden_model_1.n2740 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2740 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2740 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2740 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2740 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2740 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2740 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wbd_ack_i , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.wbd_dat_i [0], xram_data_in_reg[0]);
  buf(\oc8051_top_1.wbd_dat_i [1], xram_data_in_reg[1]);
  buf(\oc8051_top_1.wbd_dat_i [2], xram_data_in_reg[2]);
  buf(\oc8051_top_1.wbd_dat_i [3], xram_data_in_reg[3]);
  buf(\oc8051_top_1.wbd_dat_i [4], xram_data_in_reg[4]);
  buf(\oc8051_top_1.wbd_dat_i [5], xram_data_in_reg[5]);
  buf(\oc8051_top_1.wbd_dat_i [6], xram_data_in_reg[6]);
  buf(\oc8051_top_1.wbd_dat_i [7], xram_data_in_reg[7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(xram_data_in_model[0], xram_data_in_reg[0]);
  buf(xram_data_in_model[1], xram_data_in_reg[1]);
  buf(xram_data_in_model[2], xram_data_in_reg[2]);
  buf(xram_data_in_model[3], xram_data_in_reg[3]);
  buf(xram_data_in_model[4], xram_data_in_reg[4]);
  buf(xram_data_in_model[5], xram_data_in_reg[5]);
  buf(xram_data_in_model[6], xram_data_in_reg[6]);
  buf(xram_data_in_model[7], xram_data_in_reg[7]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(xram_addr_gm[0], \oc8051_golden_model_1.XRAM_ADDR [0]);
  buf(xram_addr_gm[1], \oc8051_golden_model_1.XRAM_ADDR [1]);
  buf(xram_addr_gm[2], \oc8051_golden_model_1.XRAM_ADDR [2]);
  buf(xram_addr_gm[3], \oc8051_golden_model_1.XRAM_ADDR [3]);
  buf(xram_addr_gm[4], \oc8051_golden_model_1.XRAM_ADDR [4]);
  buf(xram_addr_gm[5], \oc8051_golden_model_1.XRAM_ADDR [5]);
  buf(xram_addr_gm[6], \oc8051_golden_model_1.XRAM_ADDR [6]);
  buf(xram_addr_gm[7], \oc8051_golden_model_1.XRAM_ADDR [7]);
  buf(xram_addr_gm[8], \oc8051_golden_model_1.XRAM_ADDR [8]);
  buf(xram_addr_gm[9], \oc8051_golden_model_1.XRAM_ADDR [9]);
  buf(xram_addr_gm[10], \oc8051_golden_model_1.XRAM_ADDR [10]);
  buf(xram_addr_gm[11], \oc8051_golden_model_1.XRAM_ADDR [11]);
  buf(xram_addr_gm[12], \oc8051_golden_model_1.XRAM_ADDR [12]);
  buf(xram_addr_gm[13], \oc8051_golden_model_1.XRAM_ADDR [13]);
  buf(xram_addr_gm[14], \oc8051_golden_model_1.XRAM_ADDR [14]);
  buf(xram_addr_gm[15], \oc8051_golden_model_1.XRAM_ADDR [15]);
  buf(xram_data_out_gm[0], \oc8051_golden_model_1.XRAM_DATA_OUT [0]);
  buf(xram_data_out_gm[1], \oc8051_golden_model_1.XRAM_DATA_OUT [1]);
  buf(xram_data_out_gm[2], \oc8051_golden_model_1.XRAM_DATA_OUT [2]);
  buf(xram_data_out_gm[3], \oc8051_golden_model_1.XRAM_DATA_OUT [3]);
  buf(xram_data_out_gm[4], \oc8051_golden_model_1.XRAM_DATA_OUT [4]);
  buf(xram_data_out_gm[5], \oc8051_golden_model_1.XRAM_DATA_OUT [5]);
  buf(xram_data_out_gm[6], \oc8051_golden_model_1.XRAM_DATA_OUT [6]);
  buf(xram_data_out_gm[7], \oc8051_golden_model_1.XRAM_DATA_OUT [7]);
  buf(TMOD_gm_next[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm_next[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm_next[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm_next[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm_next[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm_next[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm_next[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm_next[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm_next[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm_next[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm_next[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm_next[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm_next[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm_next[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm_next[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm_next[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm_next[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm_next[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm_next[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm_next[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm_next[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm_next[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm_next[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm_next[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm_next[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm_next[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm_next[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm_next[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm_next[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm_next[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm_next[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm_next[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm_next[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm_next[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm_next[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm_next[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm_next[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm_next[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm_next[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm_next[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm_next[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm_next[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm_next[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm_next[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm_next[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm_next[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm_next[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm_next[7], \oc8051_golden_model_1.TCON [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm_next[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm_next[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm_next[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm_next[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm_next[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm_next[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm_next[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm_next[7], \oc8051_golden_model_1.SCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm_next[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm_next[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm_next[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm_next[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm_next[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm_next[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm_next[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm_next[7], \oc8051_golden_model_1.SBUF [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm_next[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm_next[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm_next[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm_next[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm_next[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm_next[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm_next[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm_next[7], \oc8051_golden_model_1.PCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm_next[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm_next[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm_next[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm_next[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm_next[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm_next[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm_next[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm_next[7], \oc8051_golden_model_1.IP [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm_next[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm_next[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm_next[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm_next[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm_next[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm_next[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm_next[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm_next[7], \oc8051_golden_model_1.IE [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(PC_gm[0], \oc8051_golden_model_1.PC [0]);
  buf(PC_gm[1], \oc8051_golden_model_1.PC [1]);
  buf(PC_gm[2], \oc8051_golden_model_1.PC [2]);
  buf(PC_gm[3], \oc8051_golden_model_1.PC [3]);
  buf(PC_gm[4], \oc8051_golden_model_1.PC [4]);
  buf(PC_gm[5], \oc8051_golden_model_1.PC [5]);
  buf(PC_gm[6], \oc8051_golden_model_1.PC [6]);
  buf(PC_gm[7], \oc8051_golden_model_1.PC [7]);
  buf(PC_gm[8], \oc8051_golden_model_1.PC [8]);
  buf(PC_gm[9], \oc8051_golden_model_1.PC [9]);
  buf(PC_gm[10], \oc8051_golden_model_1.PC [10]);
  buf(PC_gm[11], \oc8051_golden_model_1.PC [11]);
  buf(PC_gm[12], \oc8051_golden_model_1.PC [12]);
  buf(PC_gm[13], \oc8051_golden_model_1.PC [13]);
  buf(PC_gm[14], \oc8051_golden_model_1.PC [14]);
  buf(PC_gm[15], \oc8051_golden_model_1.PC [15]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc_impl[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc_impl[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc_impl[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc_impl[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc_impl[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc_impl[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc_impl[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc_impl[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc_impl[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc_impl[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc_impl[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc_impl[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc_impl[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc_impl[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc_impl[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc_impl[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(wbd_ack_i, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_i[0], xram_data_in_reg[0]);
  buf(wbd_dat_i[1], xram_data_in_reg[1]);
  buf(wbd_dat_i[2], xram_data_in_reg[2]);
  buf(wbd_dat_i[3], xram_data_in_reg[3]);
  buf(wbd_dat_i[4], xram_data_in_reg[4]);
  buf(wbd_dat_i[5], xram_data_in_reg[5]);
  buf(wbd_dat_i[6], xram_data_in_reg[6]);
  buf(wbd_dat_i[7], xram_data_in_reg[7]);
  buf(property_invalid_dec_rom_pc, 1'b0);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
