
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire _44061_;
  wire _44062_;
  wire _44063_;
  wire _44064_;
  wire _44065_;
  wire _44066_;
  wire _44067_;
  wire _44068_;
  wire _44069_;
  wire _44070_;
  wire _44071_;
  wire _44072_;
  wire _44073_;
  wire _44074_;
  wire _44075_;
  wire _44076_;
  wire _44077_;
  wire _44078_;
  wire _44079_;
  wire _44080_;
  wire _44081_;
  wire _44082_;
  wire _44083_;
  wire _44084_;
  wire _44085_;
  wire _44086_;
  wire _44087_;
  wire _44088_;
  wire _44089_;
  wire _44090_;
  wire _44091_;
  wire _44092_;
  wire _44093_;
  wire _44094_;
  wire _44095_;
  wire _44096_;
  wire _44097_;
  wire _44098_;
  wire _44099_;
  wire _44100_;
  wire _44101_;
  wire _44102_;
  wire _44103_;
  wire _44104_;
  wire _44105_;
  wire _44106_;
  wire _44107_;
  wire _44108_;
  wire _44109_;
  wire _44110_;
  wire _44111_;
  wire _44112_;
  wire _44113_;
  wire _44114_;
  wire _44115_;
  wire _44116_;
  wire _44117_;
  wire _44118_;
  wire _44119_;
  wire _44120_;
  wire _44121_;
  wire _44122_;
  wire _44123_;
  wire _44124_;
  wire _44125_;
  wire _44126_;
  wire _44127_;
  wire _44128_;
  wire _44129_;
  wire _44130_;
  wire _44131_;
  wire _44132_;
  wire _44133_;
  wire _44134_;
  wire _44135_;
  wire _44136_;
  wire _44137_;
  wire _44138_;
  wire _44139_;
  wire _44140_;
  wire _44141_;
  wire _44142_;
  wire _44143_;
  wire _44144_;
  wire _44145_;
  wire _44146_;
  wire _44147_;
  wire _44148_;
  wire _44149_;
  wire _44150_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1071 ;
  wire [3:0] \oc8051_golden_model_1.n1073 ;
  wire [3:0] \oc8051_golden_model_1.n1075 ;
  wire [3:0] \oc8051_golden_model_1.n1076 ;
  wire [3:0] \oc8051_golden_model_1.n1077 ;
  wire [3:0] \oc8051_golden_model_1.n1078 ;
  wire [3:0] \oc8051_golden_model_1.n1079 ;
  wire [3:0] \oc8051_golden_model_1.n1080 ;
  wire [3:0] \oc8051_golden_model_1.n1081 ;
  wire \oc8051_golden_model_1.n1118 ;
  wire \oc8051_golden_model_1.n1146 ;
  wire [8:0] \oc8051_golden_model_1.n1147 ;
  wire [8:0] \oc8051_golden_model_1.n1148 ;
  wire [7:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1150 ;
  wire \oc8051_golden_model_1.n1151 ;
  wire [2:0] \oc8051_golden_model_1.n1152 ;
  wire \oc8051_golden_model_1.n1153 ;
  wire [1:0] \oc8051_golden_model_1.n1154 ;
  wire [7:0] \oc8051_golden_model_1.n1155 ;
  wire [15:0] \oc8051_golden_model_1.n1181 ;
  wire [7:0] \oc8051_golden_model_1.n1183 ;
  wire [8:0] \oc8051_golden_model_1.n1185 ;
  wire [8:0] \oc8051_golden_model_1.n1189 ;
  wire \oc8051_golden_model_1.n1190 ;
  wire [3:0] \oc8051_golden_model_1.n1191 ;
  wire [4:0] \oc8051_golden_model_1.n1192 ;
  wire [4:0] \oc8051_golden_model_1.n1196 ;
  wire \oc8051_golden_model_1.n1197 ;
  wire [8:0] \oc8051_golden_model_1.n1198 ;
  wire \oc8051_golden_model_1.n1206 ;
  wire [7:0] \oc8051_golden_model_1.n1207 ;
  wire [8:0] \oc8051_golden_model_1.n1211 ;
  wire \oc8051_golden_model_1.n1212 ;
  wire [4:0] \oc8051_golden_model_1.n1217 ;
  wire \oc8051_golden_model_1.n1218 ;
  wire \oc8051_golden_model_1.n1226 ;
  wire [7:0] \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1229 ;
  wire [8:0] \oc8051_golden_model_1.n1231 ;
  wire \oc8051_golden_model_1.n1232 ;
  wire [3:0] \oc8051_golden_model_1.n1233 ;
  wire [4:0] \oc8051_golden_model_1.n1234 ;
  wire [4:0] \oc8051_golden_model_1.n1236 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [7:0] \oc8051_golden_model_1.n1246 ;
  wire [8:0] \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1257 ;
  wire [7:0] \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [4:0] \oc8051_golden_model_1.n1278 ;
  wire \oc8051_golden_model_1.n1279 ;
  wire [7:0] \oc8051_golden_model_1.n1280 ;
  wire [8:0] \oc8051_golden_model_1.n1282 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1290 ;
  wire [7:0] \oc8051_golden_model_1.n1291 ;
  wire [7:0] \oc8051_golden_model_1.n1292 ;
  wire [8:0] \oc8051_golden_model_1.n1295 ;
  wire [8:0] \oc8051_golden_model_1.n1296 ;
  wire [7:0] \oc8051_golden_model_1.n1297 ;
  wire \oc8051_golden_model_1.n1298 ;
  wire [7:0] \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [8:0] \oc8051_golden_model_1.n1303 ;
  wire [8:0] \oc8051_golden_model_1.n1305 ;
  wire \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1307 ;
  wire [4:0] \oc8051_golden_model_1.n1309 ;
  wire \oc8051_golden_model_1.n1310 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire [7:0] \oc8051_golden_model_1.n1318 ;
  wire [8:0] \oc8051_golden_model_1.n1322 ;
  wire \oc8051_golden_model_1.n1323 ;
  wire [4:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire [7:0] \oc8051_golden_model_1.n1334 ;
  wire [8:0] \oc8051_golden_model_1.n1338 ;
  wire \oc8051_golden_model_1.n1339 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire [7:0] \oc8051_golden_model_1.n1350 ;
  wire [8:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [4:0] \oc8051_golden_model_1.n1357 ;
  wire \oc8051_golden_model_1.n1358 ;
  wire \oc8051_golden_model_1.n1365 ;
  wire [7:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1520 ;
  wire [6:0] \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [3:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire [7:0] \oc8051_golden_model_1.n1555 ;
  wire [7:0] \oc8051_golden_model_1.n1680 ;
  wire \oc8051_golden_model_1.n1683 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire \oc8051_golden_model_1.n1691 ;
  wire [7:0] \oc8051_golden_model_1.n1692 ;
  wire \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1698 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire \oc8051_golden_model_1.n1709 ;
  wire \oc8051_golden_model_1.n1711 ;
  wire \oc8051_golden_model_1.n1717 ;
  wire [7:0] \oc8051_golden_model_1.n1718 ;
  wire \oc8051_golden_model_1.n1722 ;
  wire \oc8051_golden_model_1.n1724 ;
  wire \oc8051_golden_model_1.n1730 ;
  wire [7:0] \oc8051_golden_model_1.n1731 ;
  wire \oc8051_golden_model_1.n1733 ;
  wire [7:0] \oc8051_golden_model_1.n1734 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire [15:0] \oc8051_golden_model_1.n1739 ;
  wire \oc8051_golden_model_1.n1745 ;
  wire [7:0] \oc8051_golden_model_1.n1746 ;
  wire \oc8051_golden_model_1.n1749 ;
  wire [7:0] \oc8051_golden_model_1.n1750 ;
  wire \oc8051_golden_model_1.n1765 ;
  wire [7:0] \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1771 ;
  wire [7:0] \oc8051_golden_model_1.n1772 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire [7:0] \oc8051_golden_model_1.n1778 ;
  wire \oc8051_golden_model_1.n1783 ;
  wire [7:0] \oc8051_golden_model_1.n1784 ;
  wire \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [7:0] \oc8051_golden_model_1.n1791 ;
  wire [3:0] \oc8051_golden_model_1.n1792 ;
  wire [7:0] \oc8051_golden_model_1.n1793 ;
  wire [7:0] \oc8051_golden_model_1.n1828 ;
  wire \oc8051_golden_model_1.n1847 ;
  wire [7:0] \oc8051_golden_model_1.n1848 ;
  wire [7:0] \oc8051_golden_model_1.n1852 ;
  wire [3:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1854 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_43223_, rst);
  not (_18778_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_18789_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18800_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18789_);
  and (_18811_, _18800_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_18822_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18789_);
  and (_18833_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18789_);
  nor (_18844_, _18833_, _18822_);
  and (_18855_, _18844_, _18811_);
  nor (_18866_, _18855_, _18778_);
  and (_18877_, _18778_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18888_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_18899_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18888_);
  nor (_18910_, _18899_, _18877_);
  not (_18921_, _18910_);
  and (_18932_, _18921_, _18855_);
  or (_18943_, _18932_, _18866_);
  and (_22107_, _18943_, _43223_);
  nor (_18964_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18975_, _18964_);
  and (_18986_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_18997_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_19008_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_19019_, _19008_);
  not (_19030_, _18899_);
  nor (_19040_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_19051_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_19062_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _19051_);
  nor (_19073_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_19084_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_19095_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _19084_);
  nor (_19106_, _19095_, _19073_);
  nor (_19117_, _19106_, _19062_);
  not (_19128_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_19139_, _19062_, _19128_);
  nor (_19150_, _19139_, _19117_);
  and (_19161_, _19150_, _19040_);
  not (_19172_, _19161_);
  and (_19183_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19194_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_19205_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19216_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _19205_);
  and (_19227_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_19238_, _19227_, _19194_);
  and (_19249_, _19238_, _19172_);
  nor (_19260_, _19249_, _19030_);
  not (_19271_, _18877_);
  nor (_19282_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_19293_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _19084_);
  nor (_19304_, _19293_, _19282_);
  nor (_19315_, _19304_, _19062_);
  not (_19326_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_19337_, _19062_, _19326_);
  nor (_19348_, _19337_, _19315_);
  and (_19359_, _19348_, _19040_);
  not (_19370_, _19359_);
  and (_19380_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_19391_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_19402_, _19391_, _19380_);
  and (_19413_, _19402_, _19370_);
  nor (_19424_, _19413_, _19271_);
  nor (_19435_, _19424_, _19260_);
  nor (_19446_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_19456_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _19084_);
  nor (_19467_, _19456_, _19446_);
  nor (_19478_, _19467_, _19062_);
  not (_19489_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_19500_, _19062_, _19489_);
  nor (_19511_, _19500_, _19478_);
  and (_19522_, _19511_, _19040_);
  not (_19533_, _19522_);
  and (_19543_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_19554_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_19565_, _19554_, _19543_);
  and (_19576_, _19565_, _19533_);
  nor (_19587_, _19576_, _18921_);
  nor (_19598_, _19587_, _18964_);
  and (_19609_, _19598_, _19435_);
  nor (_19620_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_19630_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _19084_);
  nor (_19641_, _19630_, _19620_);
  nor (_19652_, _19641_, _19062_);
  not (_19663_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_19674_, _19062_, _19663_);
  nor (_19685_, _19674_, _19652_);
  and (_19696_, _19685_, _19040_);
  not (_19707_, _19696_);
  and (_19717_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_19728_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_19750_, _19728_, _19717_);
  and (_19762_, _19750_, _19707_);
  and (_19774_, _19762_, _18964_);
  nor (_19786_, _19774_, _19609_);
  not (_19797_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19809_, _19797_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19821_, _19809_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19822_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_19833_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19844_, _19833_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19855_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_19866_, _19855_, _19822_);
  nor (_19877_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19887_, _19877_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19898_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_19909_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19920_, _19809_, _19909_);
  and (_19931_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_19942_, _19931_, _19898_);
  and (_19953_, _19942_, _19866_);
  and (_19964_, _19877_, _19797_);
  and (_19974_, _19964_, _19685_);
  and (_19985_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19996_, _19985_, _19909_);
  and (_20007_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_20018_, _19985_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_20029_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_20040_, _20029_, _20007_);
  not (_20050_, _20040_);
  nor (_20061_, _20050_, _19974_);
  and (_20072_, _20061_, _19953_);
  not (_20083_, _20072_);
  and (_20094_, _20083_, _19786_);
  not (_20105_, _20094_);
  nor (_20116_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_20127_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _19084_);
  nor (_20137_, _20127_, _20116_);
  nor (_20148_, _20137_, _19062_);
  not (_20159_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_20170_, _19062_, _20159_);
  nor (_20181_, _20170_, _20148_);
  and (_20192_, _20181_, _19040_);
  not (_20203_, _20192_);
  and (_20214_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_20224_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_20235_, _20224_, _20214_);
  and (_20246_, _20235_, _20203_);
  nor (_20257_, _20246_, _19030_);
  nor (_20268_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_20279_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _19084_);
  nor (_20290_, _20279_, _20268_);
  nor (_20301_, _20290_, _19062_);
  not (_20311_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_20322_, _19062_, _20311_);
  nor (_20333_, _20322_, _20301_);
  and (_20344_, _20333_, _19040_);
  not (_20355_, _20344_);
  and (_20366_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_20377_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_20388_, _20377_, _20366_);
  and (_20398_, _20388_, _20355_);
  nor (_20409_, _20398_, _19271_);
  nor (_20420_, _20409_, _20257_);
  nor (_20431_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_20442_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _19084_);
  nor (_20453_, _20442_, _20431_);
  nor (_20464_, _20453_, _19062_);
  not (_20474_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_20485_, _19062_, _20474_);
  nor (_20496_, _20485_, _20464_);
  and (_20507_, _20496_, _19040_);
  not (_20518_, _20507_);
  and (_20529_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_20540_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_20551_, _20540_, _20529_);
  and (_20561_, _20551_, _20518_);
  nor (_20572_, _20561_, _18921_);
  nor (_20583_, _20572_, _18964_);
  and (_20594_, _20583_, _20420_);
  nor (_20605_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_20616_, _19084_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_20627_, _20616_, _20605_);
  nor (_20638_, _20627_, _19062_);
  not (_20658_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_20669_, _19062_, _20658_);
  nor (_20670_, _20669_, _20638_);
  and (_20681_, _20670_, _19040_);
  not (_20702_, _20681_);
  and (_20713_, _19183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20714_, _19216_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_20735_, _20714_, _20713_);
  and (_20745_, _20735_, _20702_);
  and (_20746_, _20745_, _18964_);
  nor (_20757_, _20746_, _20594_);
  and (_20768_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_20779_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_20800_, _20779_, _20768_);
  and (_20801_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20812_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_20823_, _20812_, _20801_);
  and (_20834_, _20823_, _20800_);
  and (_20844_, _20670_, _19964_);
  and (_20855_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_20866_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_20877_, _20866_, _20855_);
  not (_20888_, _20877_);
  nor (_20899_, _20888_, _20844_);
  and (_20910_, _20899_, _20834_);
  not (_20930_, _20910_);
  and (_20931_, _20930_, _20757_);
  and (_20942_, _20931_, _20105_);
  not (_20953_, _20942_);
  and (_20964_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_20975_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_20986_, _20975_, _20964_);
  and (_20997_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_21008_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_21019_, _21008_, _20997_);
  and (_21029_, _21019_, _20986_);
  and (_21040_, _20333_, _19964_);
  and (_21051_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_21062_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_21073_, _21062_, _21051_);
  not (_21084_, _21073_);
  nor (_21105_, _21084_, _21040_);
  and (_21106_, _21105_, _21029_);
  not (_21116_, _21106_);
  and (_21127_, _21116_, _20757_);
  and (_21138_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_21149_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_21160_, _21149_, _21138_);
  and (_21171_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_21182_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_21193_, _21182_, _21171_);
  and (_21204_, _21193_, _21160_);
  and (_21214_, _19964_, _19348_);
  and (_21225_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_21236_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_21247_, _21236_, _21225_);
  not (_21258_, _21247_);
  nor (_21269_, _21258_, _21214_);
  and (_21280_, _21269_, _21204_);
  not (_21300_, _21280_);
  and (_21301_, _21300_, _19786_);
  and (_21312_, _21301_, _21127_);
  and (_21323_, _21312_, _20083_);
  nor (_21334_, _21312_, _20094_);
  nor (_21345_, _21334_, _21323_);
  and (_21356_, _21345_, _21127_);
  and (_21367_, _20931_, _20094_);
  and (_21378_, _20757_, _20083_);
  and (_21389_, _20930_, _19786_);
  nor (_21399_, _21389_, _21378_);
  nor (_21410_, _21399_, _21367_);
  and (_21421_, _21410_, _21356_);
  nor (_21432_, _21410_, _21356_);
  nor (_21443_, _21432_, _21421_);
  and (_21454_, _21443_, _21323_);
  nor (_21465_, _21454_, _21421_);
  nor (_21476_, _21465_, _20953_);
  and (_21486_, _21465_, _20953_);
  nor (_21497_, _21486_, _21476_);
  not (_21508_, _21497_);
  and (_21519_, _21300_, _20757_);
  and (_21530_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_21541_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_21552_, _21541_, _21530_);
  and (_21563_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_21574_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_21584_, _21574_, _21563_);
  and (_21595_, _21584_, _21552_);
  and (_21606_, _20181_, _19964_);
  and (_21617_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_21628_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_21649_, _21628_, _21617_);
  not (_21650_, _21649_);
  nor (_21661_, _21650_, _21606_);
  and (_21672_, _21661_, _21595_);
  not (_21682_, _21672_);
  and (_21693_, _21682_, _19786_);
  and (_21704_, _21693_, _21519_);
  and (_21715_, _21116_, _19786_);
  nor (_21726_, _21715_, _21519_);
  nor (_21737_, _21726_, _21312_);
  and (_21758_, _21737_, _21704_);
  nor (_21759_, _21127_, _20094_);
  nor (_21769_, _21759_, _21356_);
  and (_21780_, _21769_, _21758_);
  nor (_21791_, _21443_, _21323_);
  nor (_21802_, _21791_, _21454_);
  and (_21813_, _21802_, _21780_);
  nor (_21824_, _21802_, _21780_);
  nor (_21835_, _21824_, _21813_);
  not (_21846_, _21835_);
  and (_21857_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_21867_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_21878_, _21867_, _21857_);
  and (_21889_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_21900_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_21911_, _21900_, _21889_);
  and (_21922_, _21911_, _21878_);
  and (_21933_, _20496_, _19964_);
  and (_21943_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_21954_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_21965_, _21954_, _21943_);
  not (_21976_, _21965_);
  nor (_21987_, _21976_, _21933_);
  and (_21998_, _21987_, _21922_);
  not (_22009_, _21998_);
  and (_22020_, _22009_, _20757_);
  and (_22030_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_22041_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_22052_, _22041_, _22030_);
  and (_22063_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_22074_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_22085_, _22074_, _22063_);
  and (_22096_, _22085_, _22052_);
  and (_22108_, _19964_, _19150_);
  and (_22118_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_22129_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_22140_, _22129_, _22118_);
  not (_22151_, _22140_);
  nor (_22162_, _22151_, _22108_);
  and (_22173_, _22162_, _22096_);
  not (_22184_, _22173_);
  and (_22204_, _22184_, _19786_);
  and (_22205_, _22204_, _22020_);
  and (_22216_, _22009_, _19786_);
  not (_22227_, _22216_);
  and (_22238_, _22184_, _20757_);
  and (_22249_, _22238_, _22227_);
  and (_22260_, _22249_, _21693_);
  nor (_22271_, _22260_, _22205_);
  and (_22282_, _21682_, _20757_);
  nor (_22292_, _22282_, _21301_);
  nor (_22303_, _22292_, _21704_);
  not (_22314_, _22303_);
  nor (_22325_, _22314_, _22271_);
  nor (_22336_, _21737_, _21704_);
  nor (_22347_, _22336_, _21758_);
  and (_22358_, _22347_, _22325_);
  nor (_22369_, _21769_, _21758_);
  nor (_22379_, _22369_, _21780_);
  and (_22390_, _22379_, _22358_);
  and (_22401_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_22412_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_22423_, _22412_, _22401_);
  and (_22434_, _19887_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_22445_, _19920_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_22455_, _22445_, _22434_);
  and (_22466_, _22455_, _22423_);
  and (_22477_, _19964_, _19511_);
  and (_22498_, _20018_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_22499_, _19996_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_22510_, _22499_, _22498_);
  not (_22521_, _22510_);
  nor (_22532_, _22521_, _22477_);
  and (_22542_, _22532_, _22466_);
  not (_22553_, _22542_);
  and (_22564_, _22553_, _20757_);
  and (_22575_, _22564_, _22216_);
  nor (_22586_, _22204_, _22020_);
  nor (_22607_, _22586_, _22205_);
  and (_22608_, _22607_, _22575_);
  nor (_22618_, _22249_, _21693_);
  nor (_22629_, _22618_, _22260_);
  and (_22640_, _22629_, _22608_);
  and (_22651_, _22314_, _22271_);
  nor (_22662_, _22651_, _22325_);
  and (_22673_, _22662_, _22640_);
  nor (_22684_, _22347_, _22325_);
  nor (_22695_, _22684_, _22358_);
  and (_22705_, _22695_, _22673_);
  nor (_22716_, _22379_, _22358_);
  nor (_22727_, _22716_, _22390_);
  and (_22738_, _22727_, _22705_);
  nor (_22749_, _22738_, _22390_);
  nor (_22760_, _22749_, _21846_);
  nor (_22771_, _22760_, _21813_);
  nor (_22782_, _22771_, _21508_);
  or (_22792_, _22782_, _21367_);
  nor (_22803_, _22792_, _21476_);
  nor (_22824_, _22803_, _19019_);
  and (_22825_, _22803_, _19019_);
  nor (_22836_, _22825_, _22824_);
  not (_22847_, _22836_);
  and (_22858_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_22869_, _22771_, _21508_);
  nor (_22879_, _22869_, _22782_);
  and (_22890_, _22879_, _22858_);
  and (_22901_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_22912_, _22749_, _21846_);
  nor (_22923_, _22912_, _22760_);
  and (_22934_, _22923_, _22901_);
  nor (_22945_, _22923_, _22901_);
  nor (_22956_, _22945_, _22934_);
  not (_22966_, _22956_);
  and (_22977_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_22988_, _22727_, _22705_);
  nor (_22999_, _22988_, _22738_);
  and (_23010_, _22999_, _22977_);
  nor (_23021_, _22999_, _22977_);
  nor (_23032_, _23021_, _23010_);
  not (_23042_, _23032_);
  and (_23053_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_23064_, _22695_, _22673_);
  nor (_23085_, _23064_, _22705_);
  and (_23086_, _23085_, _23053_);
  nor (_23097_, _23085_, _23053_);
  nor (_23108_, _23097_, _23086_);
  not (_23119_, _23108_);
  and (_23130_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_23141_, _22662_, _22640_);
  nor (_23151_, _23141_, _22673_);
  and (_23162_, _23151_, _23130_);
  and (_23173_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_23184_, _22629_, _22608_);
  nor (_23195_, _23184_, _22640_);
  and (_23206_, _23195_, _23173_);
  and (_23217_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_23228_, _22607_, _22575_);
  nor (_23239_, _23228_, _22608_);
  and (_23250_, _23239_, _23217_);
  nor (_23260_, _23195_, _23173_);
  nor (_23271_, _23260_, _23206_);
  and (_23282_, _23271_, _23250_);
  nor (_23293_, _23282_, _23206_);
  not (_23304_, _23293_);
  nor (_23315_, _23151_, _23130_);
  nor (_23326_, _23315_, _23162_);
  and (_23337_, _23326_, _23304_);
  nor (_23348_, _23337_, _23162_);
  nor (_23369_, _23348_, _23119_);
  nor (_23370_, _23369_, _23086_);
  nor (_23380_, _23370_, _23042_);
  nor (_23391_, _23380_, _23010_);
  nor (_23402_, _23391_, _22966_);
  nor (_23413_, _23402_, _22934_);
  nor (_23424_, _22879_, _22858_);
  nor (_23435_, _23424_, _22890_);
  not (_23446_, _23435_);
  nor (_23457_, _23446_, _23413_);
  nor (_23468_, _23457_, _22890_);
  nor (_23479_, _23468_, _22847_);
  nor (_23489_, _23479_, _22824_);
  not (_23500_, _23489_);
  and (_23511_, _23500_, _18997_);
  and (_23522_, _23511_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_23533_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_23544_, _23533_, _23522_);
  and (_23555_, _23544_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_23566_, _23555_, _18986_);
  not (_23577_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_23588_, _18964_, _23577_);
  or (_23598_, _23588_, _23566_);
  nand (_23609_, _23566_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and (_23620_, _23609_, _23598_);
  and (_24267_, _23620_, _43223_);
  nor (_23641_, _18855_, _18888_);
  and (_23652_, _18855_, _18888_);
  or (_23663_, _23652_, _23641_);
  and (_02346_, _23663_, _43223_);
  and (_23684_, _22553_, _19786_);
  and (_02538_, _23684_, _43223_);
  nor (_23704_, _22564_, _22216_);
  nor (_23715_, _23704_, _22575_);
  and (_02716_, _23715_, _43223_);
  nor (_23736_, _23239_, _23217_);
  nor (_23747_, _23736_, _23250_);
  and (_02889_, _23747_, _43223_);
  nor (_23768_, _23271_, _23250_);
  nor (_23779_, _23768_, _23282_);
  and (_03129_, _23779_, _43223_);
  nor (_23800_, _23326_, _23304_);
  nor (_23810_, _23800_, _23337_);
  and (_03335_, _23810_, _43223_);
  and (_23831_, _23348_, _23119_);
  nor (_23842_, _23831_, _23369_);
  and (_03513_, _23842_, _43223_);
  and (_23863_, _23370_, _23042_);
  nor (_23874_, _23863_, _23380_);
  and (_03714_, _23874_, _43223_);
  and (_23894_, _23391_, _22966_);
  nor (_23905_, _23894_, _23402_);
  and (_03913_, _23905_, _43223_);
  and (_23926_, _23446_, _23413_);
  nor (_23937_, _23926_, _23457_);
  and (_04014_, _23937_, _43223_);
  and (_23958_, _23468_, _22847_);
  nor (_23978_, _23958_, _23479_);
  and (_04110_, _23978_, _43223_);
  nor (_23989_, _23500_, _18997_);
  nor (_24000_, _23989_, _23511_);
  and (_04209_, _24000_, _43223_);
  and (_24021_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_24032_, _24021_, _23511_);
  nor (_24043_, _24032_, _23522_);
  and (_04309_, _24043_, _43223_);
  nor (_24063_, _23533_, _23522_);
  nor (_24074_, _24063_, _23544_);
  and (_04408_, _24074_, _43223_);
  and (_24095_, _18975_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_24106_, _24095_, _23544_);
  nor (_24117_, _24106_, _23555_);
  and (_04502_, _24117_, _43223_);
  nor (_24137_, _23555_, _18986_);
  nor (_24148_, _24137_, _23566_);
  and (_04600_, _24148_, _43223_);
  and (_24169_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18789_);
  nor (_24180_, _24169_, _18800_);
  not (_24191_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_24202_, _18822_, _24191_);
  and (_24213_, _24202_, _24180_);
  and (_24223_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24234_, _24223_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24245_, _24223_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24256_, _24245_, _24234_);
  and (_00924_, _24256_, _43223_);
  and (_00953_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _43223_);
  not (_24288_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_24299_, _20561_, _24288_);
  and (_24309_, _20246_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24320_, _24309_, _24299_);
  nor (_24331_, _24320_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24342_, _20398_, _24288_);
  and (_24353_, _20745_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24364_, _24353_, _24342_);
  and (_24375_, _24364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24385_, _24375_, _24331_);
  nor (_24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24407_, _24396_, _20910_);
  nor (_24418_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_24429_, _24418_, _24407_);
  not (_24440_, _24429_);
  and (_24451_, _19576_, _24288_);
  and (_24461_, _19249_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24472_, _24461_, _24451_);
  nor (_24483_, _24472_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24504_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24505_, _19413_, _24288_);
  and (_24516_, _19762_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24527_, _24516_, _24505_);
  nor (_24538_, _24527_, _24504_);
  nor (_24548_, _24538_, _24483_);
  nor (_24559_, _24548_, _24440_);
  and (_24570_, _24548_, _24440_);
  nor (_24581_, _24570_, _24559_);
  and (_24592_, _24396_, _20072_);
  nor (_24603_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_24614_, _24603_, _24592_);
  not (_24625_, _24614_);
  nor (_24635_, _20561_, _24288_);
  nor (_24646_, _24635_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24657_, _20246_, _24288_);
  and (_24668_, _20398_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24679_, _24668_, _24657_);
  nor (_24690_, _24679_, _24504_);
  nor (_24701_, _24690_, _24646_);
  nor (_24712_, _24701_, _24625_);
  and (_24722_, _24701_, _24625_);
  nor (_24733_, _24722_, _24712_);
  not (_24744_, _24733_);
  and (_24755_, _24396_, _21106_);
  nor (_24766_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor (_24777_, _24766_, _24755_);
  not (_24788_, _24777_);
  nor (_24799_, _19576_, _24288_);
  nor (_24809_, _24799_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24820_, _19249_, _24288_);
  and (_24831_, _19413_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24842_, _24831_, _24820_);
  nor (_24853_, _24842_, _24504_);
  nor (_24864_, _24853_, _24809_);
  nor (_24875_, _24864_, _24788_);
  and (_24886_, _24864_, _24788_);
  and (_24896_, _24320_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24907_, _24896_);
  nor (_24918_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_24929_, _24396_, _21280_);
  nor (_24940_, _24929_, _24918_);
  and (_24951_, _24940_, _24907_);
  and (_24962_, _24472_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24972_, _24962_);
  nor (_24983_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  and (_24994_, _24396_, _21672_);
  nor (_25005_, _24994_, _24983_);
  and (_25016_, _25005_, _24972_);
  nor (_25027_, _25005_, _24972_);
  nor (_25048_, _25027_, _25016_);
  not (_25049_, _25048_);
  and (_25060_, _24635_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25071_, _25060_);
  and (_25082_, _24396_, _22173_);
  nor (_25093_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_25104_, _25093_, _25082_);
  and (_25115_, _25104_, _25071_);
  and (_25126_, _24799_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25137_, _25126_);
  and (_25148_, _24396_, _21998_);
  nor (_25159_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  nor (_25170_, _25159_, _25148_);
  nor (_25181_, _25170_, _25137_);
  not (_25192_, _25181_);
  nor (_25203_, _25104_, _25071_);
  nor (_25214_, _25203_, _25115_);
  and (_25225_, _25214_, _25192_);
  nor (_25235_, _25225_, _25115_);
  nor (_25246_, _25235_, _25049_);
  nor (_25257_, _25246_, _25016_);
  nor (_25268_, _24940_, _24907_);
  nor (_25279_, _25268_, _24951_);
  not (_25290_, _25279_);
  nor (_25311_, _25290_, _25257_);
  nor (_25312_, _25311_, _24951_);
  nor (_25323_, _25312_, _24886_);
  nor (_25334_, _25323_, _24875_);
  nor (_25345_, _25334_, _24744_);
  nor (_25356_, _25345_, _24712_);
  not (_25367_, _25356_);
  and (_25378_, _25367_, _24581_);
  or (_25389_, _25378_, _24559_);
  and (_25400_, _20745_, _19762_);
  or (_25411_, _25400_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_25422_, _24527_);
  and (_25433_, _24364_, _25422_);
  nor (_25444_, _24842_, _24679_);
  and (_25455_, _25444_, _25433_);
  or (_25466_, _25455_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_25477_, _25466_, _25411_);
  and (_25488_, _25477_, _25389_);
  and (_25499_, _25488_, _24385_);
  nor (_25510_, _25367_, _24581_);
  or (_25521_, _25510_, _25378_);
  and (_25532_, _25521_, _25499_);
  nor (_25543_, _25499_, _24429_);
  nor (_25554_, _25543_, _25532_);
  not (_25565_, _25554_);
  and (_25576_, _25554_, _24385_);
  not (_25587_, _24548_);
  nor (_25598_, _25499_, _24625_);
  and (_25619_, _25334_, _24744_);
  nor (_25620_, _25619_, _25345_);
  and (_25631_, _25620_, _25499_);
  or (_25641_, _25631_, _25598_);
  and (_25652_, _25641_, _25587_);
  nor (_25663_, _25641_, _25587_);
  nor (_25674_, _25663_, _25652_);
  not (_25685_, _25674_);
  not (_25696_, _24701_);
  nor (_25707_, _25499_, _24788_);
  nor (_25718_, _24886_, _24875_);
  nor (_25729_, _25718_, _25312_);
  and (_25740_, _25718_, _25312_);
  or (_25751_, _25740_, _25729_);
  and (_25762_, _25751_, _25499_);
  or (_25773_, _25762_, _25707_);
  and (_25784_, _25773_, _25696_);
  nor (_25795_, _25773_, _25696_);
  not (_25806_, _24864_);
  and (_25817_, _25290_, _25257_);
  or (_25828_, _25817_, _25311_);
  and (_25839_, _25828_, _25499_);
  nor (_25850_, _25499_, _24940_);
  nor (_25861_, _25850_, _25839_);
  and (_25872_, _25861_, _25806_);
  and (_25883_, _25235_, _25049_);
  nor (_25894_, _25883_, _25246_);
  not (_25905_, _25894_);
  and (_25916_, _25905_, _25499_);
  nor (_25927_, _25499_, _25005_);
  nor (_25948_, _25927_, _25916_);
  and (_25949_, _25948_, _24907_);
  nor (_25960_, _25948_, _24907_);
  nor (_25971_, _25960_, _25949_);
  not (_25982_, _25971_);
  nor (_25993_, _25214_, _25192_);
  nor (_26004_, _25993_, _25225_);
  not (_26014_, _26004_);
  and (_26025_, _26014_, _25499_);
  nor (_26036_, _25499_, _25104_);
  nor (_26047_, _26036_, _26025_);
  and (_26058_, _26047_, _24972_);
  not (_26069_, _25170_);
  and (_26080_, _25499_, _25126_);
  or (_26091_, _26080_, _26069_);
  nand (_26102_, _25499_, _25126_);
  or (_26113_, _26102_, _25170_);
  and (_26124_, _26113_, _26091_);
  nor (_26135_, _26124_, _25060_);
  and (_26146_, _26124_, _25060_);
  nor (_26157_, _26146_, _26135_);
  and (_26168_, _24396_, _22542_);
  nor (_26179_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_26190_, _26179_, _26168_);
  nor (_26201_, _26190_, _25137_);
  not (_26212_, _26201_);
  and (_26223_, _26212_, _26157_);
  nor (_26234_, _26223_, _26135_);
  nor (_26245_, _26047_, _24972_);
  nor (_26256_, _26245_, _26058_);
  not (_26267_, _26256_);
  nor (_26278_, _26267_, _26234_);
  nor (_26289_, _26278_, _26058_);
  nor (_26300_, _26289_, _25982_);
  nor (_26311_, _26300_, _25949_);
  nor (_26322_, _25861_, _25806_);
  nor (_26333_, _26322_, _25872_);
  not (_26344_, _26333_);
  nor (_26354_, _26344_, _26311_);
  nor (_26365_, _26354_, _25872_);
  nor (_26376_, _26365_, _25795_);
  nor (_26387_, _26376_, _25784_);
  nor (_26398_, _26387_, _25685_);
  or (_26409_, _26398_, _25652_);
  or (_26430_, _26409_, _25576_);
  and (_26431_, _26430_, _25477_);
  nor (_26442_, _26431_, _25565_);
  and (_26453_, _25576_, _25477_);
  and (_26464_, _26453_, _26409_);
  or (_26475_, _26464_, _26442_);
  and (_00973_, _26475_, _43223_);
  or (_26496_, _25554_, _24385_);
  and (_26507_, _26496_, _26431_);
  and (_02843_, _26507_, _43223_);
  and (_02854_, _25499_, _43223_);
  and (_02876_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _43223_);
  and (_02902_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _43223_);
  and (_02927_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _43223_);
  or (_26568_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_26579_, _24223_, rst);
  and (_02938_, _26579_, _26568_);
  and (_26600_, _26507_, _25126_);
  or (_26611_, _26600_, _26190_);
  nand (_26622_, _26600_, _26190_);
  and (_26633_, _26622_, _26611_);
  and (_02951_, _26633_, _43223_);
  nor (_26654_, _26507_, _26124_);
  nor (_26665_, _26212_, _26157_);
  nor (_26676_, _26665_, _26223_);
  and (_26687_, _26676_, _26507_);
  or (_26697_, _26687_, _26654_);
  and (_02963_, _26697_, _43223_);
  and (_26718_, _26267_, _26234_);
  or (_26729_, _26718_, _26278_);
  nand (_26740_, _26729_, _26507_);
  or (_26751_, _26507_, _26047_);
  and (_26762_, _26751_, _26740_);
  and (_02975_, _26762_, _43223_);
  and (_26783_, _26289_, _25982_);
  or (_26794_, _26783_, _26300_);
  nand (_26805_, _26794_, _26507_);
  or (_26816_, _26507_, _25948_);
  and (_26827_, _26816_, _26805_);
  and (_02988_, _26827_, _43223_);
  and (_26848_, _26344_, _26311_);
  or (_26859_, _26848_, _26354_);
  nand (_26870_, _26859_, _26507_);
  or (_26881_, _26507_, _25861_);
  and (_26892_, _26881_, _26870_);
  and (_03000_, _26892_, _43223_);
  or (_26913_, _25795_, _25784_);
  and (_26924_, _26913_, _26365_);
  nor (_26935_, _26913_, _26365_);
  or (_26946_, _26935_, _26924_);
  nand (_26957_, _26946_, _26507_);
  or (_26968_, _26507_, _25773_);
  and (_26979_, _26968_, _26957_);
  and (_03011_, _26979_, _43223_);
  and (_27000_, _26387_, _25685_);
  or (_27011_, _27000_, _26398_);
  nand (_27022_, _27011_, _26507_);
  or (_27033_, _26507_, _25641_);
  and (_27043_, _27033_, _27022_);
  and (_03024_, _27043_, _43223_);
  not (_27064_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27075_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18789_);
  and (_27086_, _27075_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_27097_, _27086_, _27064_);
  and (_27108_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27119_, _27108_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_27130_, _27108_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_27141_, _27130_, _27119_);
  and (_27152_, _27141_, _27097_);
  not (_27163_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_27174_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18789_);
  and (_27185_, _27174_, _27064_);
  and (_27196_, _27185_, _27163_);
  and (_27207_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_27228_, _27207_, _27152_);
  not (_27229_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_27240_, _27075_, _27229_);
  and (_27251_, _27240_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27262_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_27273_, _27240_, _27064_);
  and (_27284_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_27295_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27306_, _27295_, _18789_);
  nor (_27317_, _27306_, _27075_);
  and (_27328_, _27317_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_27339_, _27328_, _27284_);
  nor (_27350_, _27339_, _27262_);
  and (_27361_, _27350_, _27228_);
  nor (_27372_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_27383_, _27372_, _27108_);
  and (_27393_, _27383_, _27097_);
  and (_27404_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_27415_, _27404_, _27393_);
  and (_27426_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_27437_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_27448_, _27317_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_27459_, _27448_, _27437_);
  nor (_27470_, _27459_, _27426_);
  and (_27481_, _27470_, _27415_);
  and (_27492_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_27503_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_27514_, _27503_, _27492_);
  and (_27525_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_27536_, _27525_);
  not (_27547_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27558_, _27097_, _27547_);
  and (_27569_, _27317_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_27580_, _27569_, _27558_);
  and (_27591_, _27580_, _27536_);
  and (_27602_, _27591_, _27514_);
  and (_27613_, _27602_, _27481_);
  and (_27624_, _27613_, _27361_);
  and (_27635_, _27119_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_27646_, _27635_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_27657_, _27646_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_27668_, _27657_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_27679_, _27668_);
  not (_27690_, _27097_);
  nor (_27701_, _27657_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_27712_, _27701_, _27690_);
  and (_27723_, _27712_, _27679_);
  not (_27734_, _27723_);
  and (_27744_, _27086_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27755_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_27766_, _27755_, _27744_);
  and (_27777_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_27788_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_27799_, _27788_, _27777_);
  and (_27810_, _27799_, _27766_);
  and (_27821_, _27810_, _27734_);
  nor (_27832_, _27646_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_27843_, _27832_);
  nor (_27864_, _27657_, _27690_);
  and (_27865_, _27864_, _27843_);
  not (_27876_, _27865_);
  and (_27887_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_27898_, _27887_, _27744_);
  and (_27909_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_27920_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_27931_, _27920_, _27909_);
  and (_27942_, _27931_, _27898_);
  and (_27953_, _27942_, _27876_);
  nor (_27964_, _27953_, _27821_);
  not (_27975_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_27986_, _27668_, _27975_);
  and (_27997_, _27668_, _27975_);
  nor (_28008_, _27997_, _27986_);
  nor (_28019_, _28008_, _27690_);
  not (_28030_, _28019_);
  and (_28041_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_28052_, _28041_);
  not (_28062_, _27744_);
  and (_28073_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_28084_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_28095_, _28084_, _28073_);
  and (_28106_, _28095_, _28062_);
  and (_28117_, _28106_, _28052_);
  and (_28128_, _28117_, _28030_);
  not (_28139_, _28128_);
  and (_28150_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_28171_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_28172_, _28171_, _28150_);
  not (_28183_, _27635_);
  nor (_28194_, _27119_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_28205_, _28194_, _27690_);
  and (_28216_, _28205_, _28183_);
  and (_28227_, _27317_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_28238_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_28249_, _28238_, _28227_);
  not (_28260_, _28249_);
  nor (_28271_, _28260_, _28216_);
  and (_28282_, _28271_, _28172_);
  not (_28293_, _28282_);
  and (_28304_, _27251_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_28315_, _28304_, _27744_);
  nor (_28326_, _27635_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_28337_, _28326_, _27690_);
  nor (_28348_, _28337_, _27646_);
  and (_28359_, _27273_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_28370_, _28359_, _28348_);
  and (_28381_, _28370_, _28315_);
  and (_28391_, _27317_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_28402_, _27196_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_28413_, _28402_, _28391_);
  and (_28424_, _28413_, _28381_);
  nor (_28435_, _28424_, _28293_);
  and (_28446_, _28435_, _28139_);
  and (_28457_, _28446_, _27964_);
  nand (_28468_, _28457_, _27624_);
  and (_28479_, _26475_, _24213_);
  not (_28490_, _28479_);
  and (_28501_, _23620_, _18855_);
  not (_28522_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_28523_, _18800_, _28522_);
  and (_28534_, _28523_, _18844_);
  not (_28545_, _28534_);
  nor (_28556_, _20910_, _20745_);
  and (_28567_, _20910_, _20745_);
  nor (_28578_, _28567_, _28556_);
  not (_28589_, _19762_);
  nor (_28600_, _20072_, _28589_);
  nor (_28611_, _20072_, _19762_);
  and (_28622_, _20072_, _19762_);
  nor (_28633_, _28622_, _28611_);
  not (_28644_, _20398_);
  nor (_28655_, _21106_, _28644_);
  nor (_28666_, _21106_, _20398_);
  and (_28677_, _21106_, _20398_);
  nor (_28688_, _28677_, _28666_);
  not (_28698_, _19413_);
  and (_28709_, _21280_, _28698_);
  nor (_28720_, _28709_, _28688_);
  nor (_28731_, _28720_, _28655_);
  nor (_28742_, _28731_, _28633_);
  nor (_28753_, _28742_, _28600_);
  and (_28764_, _28731_, _28633_);
  nor (_28775_, _28764_, _28742_);
  not (_28786_, _28775_);
  and (_28797_, _28709_, _28688_);
  nor (_28808_, _28797_, _28720_);
  not (_28819_, _28808_);
  nor (_28830_, _21280_, _19413_);
  and (_28841_, _21280_, _19413_);
  nor (_28852_, _28841_, _28830_);
  not (_28863_, _28852_);
  and (_28874_, _21672_, _20246_);
  nor (_28895_, _21672_, _20246_);
  nor (_28896_, _28895_, _28874_);
  nor (_28907_, _22173_, _19249_);
  and (_28918_, _22173_, _19249_);
  nor (_28929_, _28918_, _28907_);
  nor (_28940_, _21998_, _20561_);
  and (_28951_, _21998_, _20561_);
  nor (_28962_, _28951_, _28940_);
  not (_28973_, _19576_);
  and (_28984_, _22542_, _28973_);
  nor (_28995_, _28984_, _28962_);
  not (_29006_, _20561_);
  nor (_29017_, _21998_, _29006_);
  nor (_29027_, _29017_, _28995_);
  nor (_29038_, _29027_, _28929_);
  not (_29049_, _19249_);
  nor (_29060_, _22173_, _29049_);
  nor (_29071_, _29060_, _29038_);
  nor (_29082_, _29071_, _28896_);
  and (_29093_, _29071_, _28896_);
  nor (_29104_, _29093_, _29082_);
  not (_29115_, _29104_);
  nor (_29126_, _22542_, _19576_);
  and (_29137_, _22542_, _19576_);
  nor (_29148_, _29137_, _29126_);
  not (_29159_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_29170_, _19062_, _29159_);
  not (_29181_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_29192_, _29181_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29203_, _29192_, _19106_);
  nor (_29214_, _29203_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_29225_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29236_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _29225_);
  and (_29247_, _29236_, _20453_);
  not (_29258_, _29247_);
  and (_29269_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29280_, _29269_, _20137_);
  nor (_29291_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29302_, _29291_, _19467_);
  nor (_29313_, _29302_, _29280_);
  and (_29324_, _29313_, _29258_);
  and (_29334_, _29324_, _29214_);
  not (_29345_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_29356_, _29192_, _19641_);
  nor (_29367_, _29356_, _29345_);
  and (_29378_, _29291_, _19304_);
  not (_29389_, _29378_);
  and (_29400_, _29269_, _20627_);
  and (_29421_, _29236_, _20290_);
  nor (_29422_, _29421_, _29400_);
  and (_29433_, _29422_, _29389_);
  and (_29444_, _29433_, _29367_);
  nor (_29455_, _29444_, _29334_);
  nor (_29466_, _29455_, _19062_);
  nor (_29477_, _29466_, _29170_);
  and (_29488_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_29499_, _29488_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_29510_, _29499_);
  and (_29521_, _29510_, _29477_);
  and (_29532_, _29510_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_29543_, _29532_, _29521_);
  nor (_29554_, _29543_, _29148_);
  and (_29565_, _29027_, _28929_);
  nor (_29576_, _29565_, _29038_);
  and (_29587_, _28984_, _28962_);
  nor (_29598_, _29587_, _28995_);
  nor (_29609_, _29598_, _29576_);
  and (_29620_, _29609_, _29554_);
  and (_29631_, _29620_, _29115_);
  not (_29641_, _20246_);
  or (_29652_, _21672_, _29641_);
  and (_29663_, _21672_, _29641_);
  or (_29674_, _29071_, _29663_);
  and (_29695_, _29674_, _29652_);
  or (_29696_, _29695_, _29631_);
  and (_29707_, _29696_, _28863_);
  and (_29718_, _29707_, _28819_);
  and (_29729_, _29718_, _28786_);
  nor (_29740_, _29729_, _28753_);
  nor (_29751_, _29740_, _28578_);
  and (_29762_, _29740_, _28578_);
  nor (_29773_, _29762_, _29751_);
  nor (_29784_, _29773_, _28545_);
  not (_29795_, _29784_);
  not (_29806_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_29817_, _24169_, _29806_);
  and (_29828_, _29817_, _18844_);
  not (_29839_, _28578_);
  not (_29850_, _28633_);
  and (_29861_, _28830_, _28688_);
  nor (_29872_, _29861_, _28666_);
  nor (_29883_, _29872_, _29850_);
  not (_29894_, _28929_);
  and (_29905_, _29126_, _28962_);
  nor (_29916_, _29905_, _28940_);
  nor (_29927_, _29916_, _29894_);
  nor (_29938_, _29927_, _28907_);
  nor (_29948_, _29938_, _28896_);
  and (_29959_, _29938_, _28896_);
  nor (_29970_, _29959_, _29948_);
  not (_29981_, _29148_);
  nor (_29992_, _29543_, _29981_);
  and (_30003_, _29992_, _28962_);
  and (_30014_, _29916_, _29894_);
  nor (_30025_, _30014_, _29927_);
  and (_30036_, _30025_, _30003_);
  not (_30047_, _30036_);
  nor (_30057_, _30047_, _29970_);
  nor (_30068_, _29938_, _28874_);
  or (_30079_, _30068_, _28895_);
  or (_30090_, _30079_, _30057_);
  and (_30101_, _30090_, _28852_);
  nor (_30112_, _28830_, _28688_);
  nor (_30123_, _30112_, _29861_);
  and (_30134_, _30123_, _30101_);
  and (_30145_, _29872_, _29850_);
  nor (_30156_, _30145_, _29883_);
  and (_30166_, _30156_, _30134_);
  or (_30177_, _30166_, _29883_);
  nor (_30188_, _30177_, _28611_);
  nor (_30199_, _30188_, _29839_);
  and (_30210_, _30188_, _29839_);
  nor (_30221_, _30210_, _30199_);
  and (_30232_, _30221_, _29828_);
  and (_30243_, _18833_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30254_, _30243_, _28523_);
  nor (_30265_, _22542_, _21998_);
  and (_30275_, _30265_, _22184_);
  and (_30286_, _30275_, _21682_);
  and (_30297_, _30286_, _21300_);
  and (_30318_, _30297_, _21116_);
  and (_30319_, _30318_, _20083_);
  and (_30330_, _30319_, _29543_);
  not (_30341_, _29543_);
  and (_30352_, _21106_, _20072_);
  and (_30363_, _22542_, _21998_);
  and (_30374_, _30363_, _22173_);
  and (_30384_, _30374_, _21672_);
  and (_30395_, _30384_, _21280_);
  and (_30406_, _30395_, _30352_);
  and (_30417_, _30406_, _30341_);
  nor (_30428_, _30417_, _30330_);
  and (_30439_, _30428_, _20910_);
  nor (_30450_, _30428_, _20910_);
  nor (_30461_, _30450_, _30439_);
  and (_30472_, _30461_, _30254_);
  not (_30483_, _20745_);
  nor (_30493_, _29543_, _30483_);
  not (_30504_, _30493_);
  and (_30515_, _29543_, _20910_);
  and (_30526_, _30243_, _18811_);
  not (_30537_, _30526_);
  nor (_30548_, _30537_, _30515_);
  and (_30559_, _30548_, _30504_);
  nor (_30570_, _30559_, _30472_);
  and (_30581_, _29817_, _24202_);
  not (_30592_, _30581_);
  and (_30603_, _22173_, _21998_);
  nor (_30613_, _30603_, _21672_);
  and (_30624_, _30613_, _30581_);
  and (_30635_, _30624_, _21300_);
  nor (_30646_, _30635_, _21116_);
  and (_30657_, _30646_, _20072_);
  nor (_30668_, _30352_, _20910_);
  nor (_30679_, _30668_, _30624_);
  and (_30690_, _30679_, _29543_);
  nor (_30701_, _30690_, _30657_);
  and (_30712_, _30701_, _20910_);
  nor (_30722_, _30701_, _20910_);
  nor (_30733_, _30722_, _30712_);
  nor (_30744_, _30733_, _30592_);
  and (_30755_, _30243_, _29817_);
  not (_30766_, _30755_);
  nor (_30777_, _30766_, _29543_);
  not (_30788_, _30777_);
  not (_30799_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30810_, _18833_, _30799_);
  and (_30820_, _30810_, _29817_);
  not (_30831_, _30820_);
  nor (_30842_, _30831_, _28567_);
  and (_30853_, _30810_, _24180_);
  and (_30864_, _30853_, _28578_);
  nor (_30875_, _30864_, _30842_);
  and (_30886_, _24202_, _18811_);
  and (_30897_, _30886_, _28556_);
  and (_30908_, _28523_, _24202_);
  and (_30919_, _30908_, _20910_);
  nor (_30930_, _30919_, _30897_);
  and (_30940_, _24180_, _18844_);
  not (_30951_, _30940_);
  nor (_30962_, _30951_, _20910_);
  and (_30973_, _30243_, _24180_);
  not (_30984_, _30973_);
  nor (_30995_, _30984_, _22542_);
  and (_31006_, _30810_, _18800_);
  not (_31028_, _31006_);
  nor (_31029_, _31028_, _20072_);
  or (_31050_, _31029_, _30995_);
  nor (_31051_, _31050_, _30962_);
  and (_31073_, _31051_, _30930_);
  and (_31074_, _31073_, _30875_);
  and (_31096_, _31074_, _30788_);
  not (_31097_, _31096_);
  nor (_31108_, _31097_, _30744_);
  and (_31119_, _31108_, _30570_);
  not (_31130_, _31119_);
  nor (_31151_, _31130_, _30232_);
  and (_31152_, _31151_, _29795_);
  not (_31172_, _31152_);
  nor (_31173_, _31172_, _28501_);
  and (_31194_, _31173_, _28490_);
  not (_31195_, _31194_);
  or (_31216_, _31195_, _28468_);
  not (_31217_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31238_, \oc8051_top_1.oc8051_decoder1.wr , _18789_);
  not (_31239_, _31238_);
  nor (_31260_, _31239_, _27185_);
  and (_31261_, _31260_, _31217_);
  not (_31281_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_31282_, _28468_, _31281_);
  and (_31303_, _31282_, _31261_);
  and (_31304_, _31303_, _31216_);
  nor (_31325_, _31260_, _31281_);
  not (_31326_, _29828_);
  nor (_31347_, _30199_, _28556_);
  nor (_31348_, _31347_, _31326_);
  not (_31369_, _31348_);
  and (_31370_, _20910_, _30483_);
  nor (_31390_, _31370_, _29751_);
  nor (_31391_, _31390_, _28545_);
  and (_31412_, _29543_, _20072_);
  and (_31413_, _31412_, _30646_);
  nor (_31434_, _31413_, _30515_);
  nor (_31435_, _29543_, _20910_);
  not (_31456_, _31435_);
  nor (_31457_, _31456_, _30657_);
  nor (_31478_, _31457_, _30592_);
  and (_31479_, _31478_, _31434_);
  or (_31499_, _31479_, _30624_);
  not (_31500_, _31499_);
  nor (_31521_, _29532_, _29477_);
  not (_31522_, _30853_);
  nor (_31543_, _31522_, _29521_);
  nor (_31544_, _31543_, _30820_);
  nor (_31565_, _31544_, _31521_);
  not (_31566_, _31565_);
  nor (_31587_, _30951_, _29543_);
  not (_31588_, _31587_);
  and (_31608_, _29499_, _29477_);
  and (_31609_, _30810_, _28523_);
  and (_31630_, _30886_, _29477_);
  nor (_31631_, _31630_, _31609_);
  nor (_31652_, _31631_, _31608_);
  not (_31653_, _31652_);
  nor (_31674_, _30984_, _29477_);
  or (_31675_, _31674_, _29543_);
  or (_31696_, _30908_, _30341_);
  and (_31697_, _31696_, _31675_);
  nor (_31717_, _30766_, _22542_);
  and (_31718_, _30810_, _18811_);
  not (_31739_, _31718_);
  nor (_31740_, _31739_, _20910_);
  nor (_31751_, _31740_, _31717_);
  not (_31762_, _31751_);
  nor (_31773_, _31762_, _31697_);
  and (_31784_, _31773_, _31653_);
  and (_31795_, _31784_, _31588_);
  and (_31806_, _31795_, _31566_);
  and (_31817_, _31806_, _31500_);
  not (_31827_, _31817_);
  nor (_31838_, _31827_, _31391_);
  and (_31849_, _31838_, _31369_);
  not (_31860_, _27361_);
  nor (_31871_, _27602_, _27481_);
  and (_31882_, _31871_, _31860_);
  and (_31893_, _31882_, _28457_);
  nand (_31904_, _31893_, _31849_);
  or (_31915_, _31893_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_31926_, _31260_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31936_, _31926_, _31915_);
  and (_31947_, _31936_, _31904_);
  or (_31958_, _31947_, _31325_);
  or (_31969_, _31958_, _31304_);
  and (_06613_, _31969_, _43223_);
  and (_31990_, _26633_, _24213_);
  not (_32001_, _31990_);
  and (_32012_, _23937_, _18855_);
  and (_32023_, _29543_, _29981_);
  nor (_32034_, _32023_, _29992_);
  and (_32044_, _29828_, _32034_);
  not (_32055_, _32044_);
  and (_32066_, _32034_, _28534_);
  not (_32077_, _32066_);
  nor (_32088_, _31739_, _29543_);
  not (_32099_, _32088_);
  nor (_32110_, _31522_, _29126_);
  nor (_32121_, _32110_, _30820_);
  or (_32132_, _32121_, _29137_);
  and (_32143_, _30886_, _29126_);
  and (_32154_, _30908_, _22542_);
  nor (_32164_, _32154_, _32143_);
  nor (_32175_, _30537_, _19576_);
  and (_32186_, _30254_, _22542_);
  nor (_32197_, _32186_, _32175_);
  nor (_32208_, _30940_, _30581_);
  nor (_32219_, _32208_, _22542_);
  not (_32230_, _32219_);
  and (_32241_, _30243_, _29806_);
  not (_32252_, _32241_);
  nor (_32263_, _32252_, _21998_);
  and (_32273_, _31609_, _20930_);
  nor (_32284_, _32273_, _32263_);
  and (_32295_, _32284_, _32230_);
  and (_32306_, _32295_, _32197_);
  and (_32317_, _32306_, _32164_);
  and (_32328_, _32317_, _32132_);
  and (_32339_, _32328_, _32099_);
  and (_32350_, _32339_, _32077_);
  and (_32361_, _32350_, _32055_);
  not (_32371_, _32361_);
  nor (_32382_, _32371_, _32012_);
  and (_32393_, _32382_, _32001_);
  not (_32404_, _32393_);
  or (_32415_, _32404_, _28468_);
  not (_32426_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_32437_, _28468_, _32426_);
  and (_32448_, _32437_, _31261_);
  and (_32459_, _32448_, _32415_);
  nor (_32470_, _31260_, _32426_);
  not (_32481_, _31849_);
  or (_32491_, _32481_, _28468_);
  and (_32502_, _32437_, _31926_);
  and (_32513_, _32502_, _32491_);
  or (_32524_, _32513_, _32470_);
  or (_32535_, _32524_, _32459_);
  and (_08854_, _32535_, _43223_);
  and (_32556_, _26697_, _24213_);
  not (_32567_, _32556_);
  and (_32578_, _23978_, _18855_);
  nor (_32589_, _29126_, _28962_);
  or (_32599_, _32589_, _29905_);
  and (_32610_, _32599_, _29992_);
  nor (_32621_, _32599_, _29992_);
  or (_32632_, _32621_, _32610_);
  and (_32643_, _32632_, _29828_);
  not (_32654_, _29598_);
  and (_32665_, _32654_, _29554_);
  nor (_32676_, _32654_, _29554_);
  nor (_32687_, _32676_, _32665_);
  nor (_32698_, _32687_, _28545_);
  nor (_32708_, _32698_, _32643_);
  nor (_32719_, _30537_, _20561_);
  nor (_32730_, _30363_, _30265_);
  not (_32741_, _32730_);
  nor (_32752_, _32741_, _29543_);
  and (_32763_, _32741_, _29543_);
  nor (_32774_, _32763_, _32752_);
  and (_32785_, _32774_, _30254_);
  nor (_32796_, _32785_, _32719_);
  nor (_32807_, _30613_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_32817_, _32807_, _22009_);
  nor (_32828_, _32807_, _22009_);
  nor (_32839_, _32828_, _32817_);
  nor (_32850_, _32839_, _30592_);
  not (_32861_, _32850_);
  and (_32872_, _30853_, _28962_);
  nor (_32883_, _30831_, _28951_);
  not (_32894_, _32883_);
  and (_32905_, _30886_, _28940_);
  and (_32916_, _30908_, _21998_);
  nor (_32926_, _32916_, _32905_);
  nand (_32937_, _32926_, _32894_);
  nor (_32948_, _32937_, _32872_);
  nor (_32959_, _31028_, _22542_);
  not (_32970_, _32959_);
  nor (_32981_, _30951_, _21998_);
  nor (_32992_, _32252_, _22173_);
  nor (_33003_, _32992_, _32981_);
  and (_33014_, _33003_, _32970_);
  and (_33025_, _33014_, _32948_);
  and (_33036_, _33025_, _32861_);
  and (_33046_, _33036_, _32796_);
  and (_33057_, _33046_, _32708_);
  not (_33068_, _33057_);
  nor (_33079_, _33068_, _32578_);
  and (_33090_, _33079_, _32567_);
  not (_33101_, _33090_);
  or (_33112_, _33101_, _28468_);
  not (_33123_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_33134_, _28468_, _33123_);
  and (_33144_, _33134_, _31261_);
  and (_33155_, _33144_, _33112_);
  nor (_33166_, _31260_, _33123_);
  not (_33177_, _27602_);
  and (_33188_, _33177_, _27481_);
  and (_33199_, _33188_, _27361_);
  and (_33210_, _33199_, _28457_);
  nand (_33221_, _33210_, _31849_);
  or (_33232_, _33210_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_33243_, _33232_, _31926_);
  and (_33254_, _33243_, _33221_);
  or (_33264_, _33254_, _33166_);
  or (_33275_, _33264_, _33155_);
  and (_08865_, _33275_, _43223_);
  and (_33296_, _26762_, _24213_);
  not (_33307_, _33296_);
  and (_33318_, _24000_, _18855_);
  nor (_33329_, _30537_, _19249_);
  and (_33340_, _30363_, _30341_);
  and (_33351_, _30265_, _29543_);
  nor (_33362_, _33351_, _33340_);
  nor (_33372_, _33362_, _22173_);
  not (_33383_, _30254_);
  and (_33394_, _33362_, _22173_);
  or (_33405_, _33394_, _33383_);
  nor (_33416_, _33405_, _33372_);
  nor (_33427_, _33416_, _33329_);
  not (_33438_, _32665_);
  and (_33449_, _33438_, _29576_);
  nor (_33460_, _33449_, _29620_);
  nor (_33471_, _33460_, _28545_);
  not (_33481_, _33471_);
  nor (_33492_, _30025_, _30003_);
  nor (_33503_, _33492_, _31326_);
  and (_33514_, _33503_, _30047_);
  nor (_33525_, _32828_, _22173_);
  and (_33536_, _30603_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33547_, _33536_, _33525_);
  nor (_33558_, _33547_, _30592_);
  nor (_33569_, _30831_, _28918_);
  and (_33580_, _30853_, _28929_);
  nor (_33590_, _33580_, _33569_);
  and (_33601_, _30886_, _28907_);
  and (_33612_, _30908_, _22173_);
  nor (_33623_, _33612_, _33601_);
  nor (_33634_, _32252_, _21672_);
  not (_33645_, _33634_);
  nor (_33656_, _30951_, _22173_);
  nor (_33667_, _31028_, _21998_);
  nor (_33678_, _33667_, _33656_);
  and (_33689_, _33678_, _33645_);
  and (_33699_, _33689_, _33623_);
  and (_33710_, _33699_, _33590_);
  not (_33721_, _33710_);
  nor (_33732_, _33721_, _33558_);
  not (_33743_, _33732_);
  nor (_33754_, _33743_, _33514_);
  and (_33765_, _33754_, _33481_);
  and (_33776_, _33765_, _33427_);
  not (_33787_, _33776_);
  nor (_33798_, _33787_, _33318_);
  and (_33809_, _33798_, _33307_);
  not (_33819_, _33809_);
  or (_33830_, _33819_, _28468_);
  not (_33841_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_33852_, _28468_, _33841_);
  and (_33863_, _33852_, _31261_);
  and (_33874_, _33863_, _33830_);
  nor (_33885_, _31260_, _33841_);
  nand (_33896_, _28457_, _27361_);
  or (_33907_, _31871_, _33896_);
  and (_33917_, _33907_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_33928_, _27481_);
  and (_33939_, _27361_, _27602_);
  and (_33950_, _33939_, _33928_);
  not (_33961_, _33950_);
  nor (_33972_, _33961_, _31849_);
  and (_33983_, _27361_, _27481_);
  and (_33994_, _33983_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_34005_, _33994_, _33972_);
  and (_34016_, _34005_, _28457_);
  or (_34026_, _34016_, _33917_);
  and (_34037_, _34026_, _31926_);
  or (_34048_, _34037_, _33885_);
  or (_34059_, _34048_, _33874_);
  and (_08876_, _34059_, _43223_);
  and (_34080_, _26827_, _24213_);
  not (_34091_, _34080_);
  and (_34102_, _24043_, _18855_);
  nor (_34113_, _29620_, _29115_);
  nor (_34124_, _34113_, _29631_);
  nor (_34135_, _34124_, _28545_);
  not (_34145_, _34135_);
  and (_34156_, _30047_, _29970_);
  or (_34169_, _34156_, _31326_);
  nor (_34188_, _34169_, _30057_);
  not (_34199_, _34188_);
  nor (_34210_, _30537_, _20246_);
  nor (_34221_, _30374_, _29543_);
  nor (_34232_, _30275_, _30341_);
  nor (_34243_, _34232_, _34221_);
  and (_34254_, _34243_, _21682_);
  not (_34264_, _34254_);
  nor (_34275_, _34243_, _21682_);
  nor (_34286_, _34275_, _33383_);
  and (_34297_, _34286_, _34264_);
  nor (_34308_, _34297_, _34210_);
  not (_34319_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_34330_, _30603_, _34319_);
  nor (_34341_, _34330_, _21682_);
  nor (_34352_, _30951_, _21672_);
  nor (_34363_, _30613_, _30592_);
  nor (_34373_, _34363_, _34352_);
  nor (_34384_, _34373_, _34341_);
  not (_34395_, _34384_);
  and (_34406_, _30853_, _28896_);
  and (_34417_, _30886_, _28895_);
  nor (_34428_, _30831_, _28874_);
  and (_34439_, _30908_, _21672_);
  or (_34450_, _34439_, _34428_);
  or (_34461_, _34450_, _34417_);
  nor (_34472_, _34461_, _34406_);
  nor (_34482_, _32252_, _21280_);
  nor (_34493_, _31028_, _22173_);
  nor (_34504_, _34493_, _34482_);
  and (_34515_, _34504_, _34472_);
  and (_34526_, _34515_, _34395_);
  and (_34537_, _34526_, _34308_);
  and (_34548_, _34537_, _34199_);
  and (_34559_, _34548_, _34145_);
  not (_34570_, _34559_);
  nor (_34581_, _34570_, _34102_);
  and (_34591_, _34581_, _34091_);
  not (_34602_, _34591_);
  or (_34613_, _34602_, _28468_);
  not (_34624_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_34635_, _28468_, _34624_);
  and (_34646_, _34635_, _31261_);
  and (_34657_, _34646_, _34613_);
  nor (_34668_, _31260_, _34624_);
  and (_34679_, _33896_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_34690_, _31871_, _27361_);
  and (_34700_, _34690_, _32481_);
  nor (_34711_, _33983_, _33939_);
  nor (_34722_, _34711_, _34624_);
  or (_34733_, _34722_, _34700_);
  and (_34744_, _34733_, _28457_);
  or (_34755_, _34744_, _34679_);
  and (_34766_, _34755_, _31926_);
  or (_34777_, _34766_, _34668_);
  or (_34788_, _34777_, _34657_);
  and (_08887_, _34788_, _43223_);
  and (_34808_, _26892_, _24213_);
  not (_34819_, _34808_);
  and (_34830_, _24074_, _18855_);
  or (_34841_, _30090_, _28852_);
  nor (_34852_, _31326_, _30101_);
  and (_34863_, _34852_, _34841_);
  nor (_34874_, _29696_, _28852_);
  and (_34885_, _29696_, _28852_);
  nor (_34896_, _34885_, _34874_);
  and (_34907_, _34896_, _28534_);
  and (_34918_, _29543_, _21300_);
  nor (_34928_, _29543_, _19413_);
  or (_34939_, _34928_, _34918_);
  and (_34950_, _34939_, _30526_);
  and (_34961_, _30286_, _29543_);
  and (_34972_, _30384_, _30341_);
  nor (_34983_, _34972_, _34961_);
  nor (_34994_, _34983_, _21280_);
  and (_35005_, _34983_, _21280_);
  or (_35016_, _35005_, _33383_);
  nor (_35027_, _35016_, _34994_);
  nor (_35037_, _35027_, _34950_);
  or (_35048_, _30624_, _21300_);
  nor (_35059_, _30635_, _30592_);
  and (_35070_, _35059_, _35048_);
  nor (_35081_, _30831_, _28841_);
  and (_35092_, _30853_, _28852_);
  nor (_35103_, _35092_, _35081_);
  and (_35114_, _30886_, _28830_);
  and (_35125_, _30908_, _21280_);
  nor (_35136_, _35125_, _35114_);
  nor (_35146_, _32252_, _21106_);
  nor (_35157_, _30951_, _21280_);
  nor (_35168_, _31028_, _21672_);
  or (_35179_, _35168_, _35157_);
  nor (_35190_, _35179_, _35146_);
  and (_35201_, _35190_, _35136_);
  nand (_35212_, _35201_, _35103_);
  nor (_35223_, _35212_, _35070_);
  nand (_35234_, _35223_, _35037_);
  or (_35245_, _35234_, _34907_);
  or (_35255_, _35245_, _34863_);
  nor (_35266_, _35255_, _34830_);
  and (_35277_, _35266_, _34819_);
  not (_35288_, _35277_);
  or (_35299_, _35288_, _28468_);
  not (_35310_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_35321_, _28468_, _35310_);
  and (_35332_, _35321_, _31261_);
  and (_35343_, _35332_, _35299_);
  nor (_35354_, _31260_, _35310_);
  not (_35364_, _28457_);
  and (_35375_, _27613_, _31860_);
  nor (_35386_, _27613_, _31860_);
  nor (_35397_, _35386_, _35375_);
  or (_35408_, _35397_, _35364_);
  and (_35419_, _35408_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_35430_, _35375_, _32481_);
  and (_35441_, _35386_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_35451_, _35441_, _35430_);
  and (_35462_, _35451_, _28457_);
  or (_35473_, _35462_, _35419_);
  and (_35484_, _35473_, _31926_);
  or (_35495_, _35484_, _35354_);
  or (_35506_, _35495_, _35343_);
  and (_08898_, _35506_, _43223_);
  and (_35527_, _26979_, _24213_);
  not (_35538_, _35527_);
  and (_35549_, _24117_, _18855_);
  nor (_35559_, _30123_, _30101_);
  not (_35570_, _35559_);
  nor (_35581_, _31326_, _30134_);
  and (_35592_, _35581_, _35570_);
  not (_35603_, _35592_);
  nor (_35614_, _29707_, _28819_);
  nor (_35625_, _35614_, _29718_);
  nor (_35636_, _35625_, _28545_);
  nor (_35647_, _29543_, _20398_);
  and (_35658_, _29543_, _21116_);
  nor (_35669_, _35658_, _35647_);
  nor (_35679_, _35669_, _30537_);
  nor (_35690_, _30297_, _30341_);
  nor (_35701_, _30395_, _29543_);
  nor (_35712_, _35701_, _35690_);
  nor (_35723_, _35712_, _21116_);
  and (_35734_, _35712_, _21116_);
  or (_35745_, _35734_, _33383_);
  nor (_35756_, _35745_, _35723_);
  nor (_35767_, _35756_, _35679_);
  not (_35778_, _30690_);
  and (_35789_, _35778_, _30646_);
  nor (_35799_, _30690_, _30635_);
  nor (_35810_, _35799_, _21106_);
  nor (_35821_, _35810_, _35789_);
  nor (_35832_, _35821_, _30592_);
  nor (_35843_, _30831_, _28677_);
  and (_35854_, _30853_, _28688_);
  nor (_35865_, _35854_, _35843_);
  and (_35876_, _30886_, _28666_);
  and (_35887_, _30908_, _21106_);
  nor (_35898_, _35887_, _35876_);
  nor (_35909_, _30951_, _21106_);
  not (_35920_, _35909_);
  nor (_35930_, _32252_, _20072_);
  nor (_35941_, _31028_, _21280_);
  nor (_35952_, _35941_, _35930_);
  and (_35963_, _35952_, _35920_);
  and (_35974_, _35963_, _35898_);
  and (_35985_, _35974_, _35865_);
  not (_35996_, _35985_);
  nor (_36007_, _35996_, _35832_);
  and (_36018_, _36007_, _35767_);
  not (_36029_, _36018_);
  nor (_36040_, _36029_, _35636_);
  and (_36050_, _36040_, _35603_);
  not (_36061_, _36050_);
  nor (_36072_, _36061_, _35549_);
  and (_36083_, _36072_, _35538_);
  not (_36094_, _36083_);
  or (_36105_, _36094_, _28468_);
  not (_36116_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_36127_, _28468_, _36116_);
  and (_36138_, _36127_, _31261_);
  and (_36149_, _36138_, _36105_);
  nor (_36160_, _31260_, _36116_);
  and (_36171_, _33188_, _31860_);
  and (_36181_, _36171_, _28457_);
  nand (_36192_, _36181_, _31849_);
  or (_36203_, _36181_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_36214_, _36203_, _31926_);
  and (_36225_, _36214_, _36192_);
  or (_36236_, _36225_, _36160_);
  or (_36247_, _36236_, _36149_);
  and (_08909_, _36247_, _43223_);
  and (_36267_, _27043_, _24213_);
  not (_36278_, _36267_);
  and (_36289_, _24148_, _18855_);
  nor (_36300_, _30156_, _30134_);
  not (_36311_, _36300_);
  nor (_36322_, _31326_, _30166_);
  and (_36333_, _36322_, _36311_);
  not (_36343_, _36333_);
  nor (_36354_, _29718_, _28786_);
  nor (_36365_, _36354_, _29729_);
  nor (_36376_, _36365_, _28545_);
  nor (_36387_, _29543_, _28589_);
  or (_36398_, _36387_, _30537_);
  nor (_36409_, _36398_, _31412_);
  nor (_36420_, _29543_, _21116_);
  nand (_36430_, _36420_, _30395_);
  nand (_36441_, _30318_, _29543_);
  and (_36452_, _36441_, _36430_);
  and (_36463_, _36452_, _20072_);
  nor (_36474_, _36452_, _20072_);
  or (_36485_, _36474_, _33383_);
  nor (_36496_, _36485_, _36463_);
  nor (_36506_, _36496_, _36409_);
  nor (_36517_, _35789_, _20072_);
  and (_36528_, _35789_, _20072_);
  nor (_36539_, _36528_, _36517_);
  nor (_36550_, _36539_, _30592_);
  and (_36561_, _30853_, _28633_);
  nor (_36572_, _30831_, _28622_);
  not (_36583_, _36572_);
  and (_36593_, _30886_, _28611_);
  and (_36604_, _30908_, _20072_);
  nor (_36615_, _36604_, _36593_);
  nand (_36626_, _36615_, _36583_);
  nor (_36637_, _36626_, _36561_);
  nor (_36648_, _30951_, _20072_);
  not (_36659_, _36648_);
  nor (_36670_, _32252_, _20910_);
  nor (_36680_, _31028_, _21106_);
  nor (_36691_, _36680_, _36670_);
  and (_36702_, _36691_, _36659_);
  and (_36713_, _36702_, _36637_);
  not (_36724_, _36713_);
  nor (_36735_, _36724_, _36550_);
  and (_36746_, _36735_, _36506_);
  not (_36757_, _36746_);
  nor (_36767_, _36757_, _36376_);
  and (_36778_, _36767_, _36343_);
  not (_36789_, _36778_);
  nor (_36800_, _36789_, _36289_);
  and (_36811_, _36800_, _36278_);
  not (_36822_, _36811_);
  or (_36833_, _36822_, _28468_);
  not (_36844_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_36855_, _28468_, _36844_);
  and (_36865_, _36855_, _31261_);
  and (_36876_, _36865_, _36833_);
  nor (_36887_, _31260_, _36844_);
  nor (_36898_, _27361_, _27481_);
  and (_36909_, _36898_, _27602_);
  and (_36920_, _36909_, _28457_);
  nand (_36931_, _36920_, _31849_);
  or (_36942_, _36920_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_36953_, _36942_, _31926_);
  and (_36964_, _36953_, _36931_);
  or (_36975_, _36964_, _36887_);
  or (_36985_, _36975_, _36876_);
  and (_08920_, _36985_, _43223_);
  and (_37006_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37017_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_37028_, _37017_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_37039_, _37028_);
  not (_37050_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_37061_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_37072_, _37061_, _37050_);
  and (_37083_, _37017_, _18789_);
  and (_37094_, _37083_, _37072_);
  not (_37105_, _37094_);
  not (_37116_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_37127_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_37138_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37149_, _37138_, _37127_);
  and (_37160_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_37171_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37182_, _37171_, _37127_);
  and (_37193_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not (_37204_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37215_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _37204_);
  and (_37226_, _37215_, _37127_);
  and (_37236_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_37247_, _37236_, _37193_);
  or (_37258_, _37247_, _37160_);
  and (_37269_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_37280_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_37291_, _37280_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37302_, _37291_, _37127_);
  and (_37313_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_37324_, _37313_, _37269_);
  nor (_37335_, _37138_, _37127_);
  and (_37345_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_37356_, _37138_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_37367_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_37378_, _37367_, _37345_);
  or (_37389_, _37378_, _37324_);
  nor (_37400_, _37389_, _37258_);
  and (_37411_, _37400_, _37116_);
  nor (_37422_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _37116_);
  nor (_37433_, _37422_, _37411_);
  nor (_37444_, _37433_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_37454_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37465_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _37454_);
  nor (_37476_, _37465_, _37444_);
  nor (_37487_, _37476_, _37105_);
  not (_37498_, _37487_);
  not (_37509_, _37072_);
  nor (_37520_, _37083_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_37531_, _37520_, _37509_);
  and (_37542_, _37531_, _37498_);
  not (_37553_, _37542_);
  and (_37564_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37574_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37585_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_37596_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_37607_, _37596_, _37585_);
  and (_37618_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37629_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_37640_, _37629_, _37618_);
  and (_37651_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_37662_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_37673_, _37662_, _37651_);
  and (_37684_, _37673_, _37640_);
  and (_37695_, _37684_, _37607_);
  nor (_37706_, _37695_, _37269_);
  and (_37717_, _37706_, _37116_);
  or (_37728_, _37717_, _37574_);
  and (_37738_, _37728_, _37454_);
  nor (_37748_, _37738_, _37564_);
  and (_37759_, _37748_, _37094_);
  not (_37770_, _37759_);
  nor (_37781_, _37083_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_37792_, _37781_, _37509_);
  and (_37803_, _37792_, _37770_);
  and (_37814_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_37825_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  or (_37836_, _37269_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37847_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_37858_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_37869_, _37858_, _37847_);
  and (_37880_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_37891_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_37902_, _37891_, _37880_);
  and (_37913_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_37924_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_37935_, _37924_, _37913_);
  and (_37946_, _37935_, _37902_);
  and (_37957_, _37946_, _37869_);
  nor (_37968_, _37957_, _37836_);
  nor (_37979_, _37968_, _37825_);
  nor (_37990_, _37979_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_38001_, _37990_, _37814_);
  and (_38012_, _38001_, _37094_);
  not (_38023_, _38012_);
  nor (_38034_, _37083_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_38045_, _38034_, _37509_);
  and (_38056_, _38045_, _38023_);
  and (_38067_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_38078_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_38089_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_38100_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_38111_, _38100_, _38089_);
  and (_38122_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_38133_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_38144_, _38133_, _38122_);
  and (_38155_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_38166_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_38177_, _38166_, _38155_);
  and (_38188_, _38177_, _38144_);
  and (_38199_, _38188_, _38111_);
  nor (_38210_, _38199_, _37836_);
  or (_38221_, _38210_, _38078_);
  and (_38232_, _38221_, _37454_);
  nor (_38243_, _38232_, _38067_);
  and (_38254_, _38243_, _37094_);
  not (_38265_, _38254_);
  nor (_38276_, _37083_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_38287_, _38276_, _37509_);
  and (_38298_, _38287_, _38265_);
  not (_38309_, _38298_);
  and (_38320_, _38309_, _38056_);
  and (_38331_, _38320_, _37803_);
  and (_38342_, _38331_, _37553_);
  and (_38353_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_38364_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_38375_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_38386_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_38396_, _38386_, _38375_);
  and (_38407_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_38418_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_38428_, _38418_, _38407_);
  and (_38439_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_38450_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_38461_, _38450_, _38439_);
  and (_38472_, _38461_, _38428_);
  and (_38483_, _38472_, _38396_);
  nor (_38494_, _38483_, _37269_);
  and (_38496_, _38494_, _37116_);
  or (_38497_, _38496_, _38364_);
  and (_38498_, _38497_, _37454_);
  nor (_38499_, _38498_, _38353_);
  and (_38500_, _38499_, _37094_);
  not (_38501_, _38500_);
  nor (_38502_, _37083_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_38503_, _38502_, _37509_);
  and (_38504_, _38503_, _38501_);
  and (_38505_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_38506_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_38507_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_38508_, _38507_, _38506_);
  or (_38509_, _38508_, _38505_);
  and (_38510_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_38511_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_38512_, _38511_, _38510_);
  and (_38513_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_38514_, _38513_, _37269_);
  nand (_38515_, _38514_, _38512_);
  nor (_38516_, _38515_, _38509_);
  and (_38517_, _38516_, _37116_);
  nor (_38518_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _37116_);
  nor (_38519_, _38518_, _38517_);
  nor (_38520_, _38519_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_38521_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _37454_);
  nor (_38522_, _38521_, _38520_);
  nor (_38523_, _38522_, _37105_);
  not (_38524_, _38523_);
  nor (_38525_, _37083_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_38526_, _38525_, _37509_);
  and (_38527_, _38526_, _38524_);
  and (_38528_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_38529_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_38530_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_38531_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_38532_, _38531_, _38530_);
  and (_38533_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_38534_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_38535_, _38534_, _38533_);
  and (_38536_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_38537_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_38538_, _38537_, _38536_);
  and (_38539_, _38538_, _38535_);
  and (_38540_, _38539_, _38532_);
  nor (_38541_, _38540_, _37836_);
  nor (_38542_, _38541_, _38529_);
  nor (_38543_, _38542_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_38544_, _38543_, _38528_);
  nor (_38545_, _38544_, _37105_);
  and (_38546_, _37105_, \oc8051_top_1.oc8051_decoder1.op [2]);
  or (_38547_, _38546_, _38545_);
  and (_38548_, _38547_, _37072_);
  and (_38549_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_38550_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_38551_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_38552_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_38553_, _38552_, _38551_);
  and (_38554_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_38555_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_38556_, _38555_, _38554_);
  and (_38557_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_38558_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_38559_, _38558_, _38557_);
  and (_38560_, _38559_, _38556_);
  and (_38561_, _38560_, _38553_);
  nor (_38562_, _38561_, _37269_);
  and (_38563_, _38562_, _37116_);
  or (_38564_, _38563_, _38550_);
  and (_38565_, _38564_, _37454_);
  nor (_38566_, _38565_, _38549_);
  and (_38567_, _38566_, _37094_);
  not (_38568_, _38567_);
  nor (_38569_, _37083_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_38570_, _38569_, _37509_);
  and (_38571_, _38570_, _38568_);
  nor (_38572_, _38571_, _38548_);
  and (_38573_, _38572_, _38527_);
  and (_38574_, _38573_, _38504_);
  and (_38575_, _38574_, _38342_);
  not (_38576_, _38056_);
  and (_38577_, _37803_, _38298_);
  and (_38578_, _38577_, _38576_);
  and (_38579_, _38578_, _37542_);
  and (_38580_, _38574_, _38579_);
  nor (_38581_, _37803_, _38298_);
  and (_38582_, _38581_, _38056_);
  and (_38583_, _38582_, _37542_);
  and (_38584_, _38574_, _38583_);
  or (_38585_, _38584_, _38580_);
  nor (_38586_, _38585_, _38575_);
  and (_38587_, _38582_, _37553_);
  not (_38588_, _38571_);
  and (_38589_, _38588_, _38548_);
  nor (_38590_, _38504_, _38527_);
  and (_38591_, _38590_, _38589_);
  and (_38592_, _38591_, _38587_);
  and (_38593_, _38591_, _38342_);
  nor (_38594_, _38593_, _38592_);
  and (_38595_, _38594_, _38586_);
  nor (_38596_, _38595_, _37039_);
  not (_38597_, _38596_);
  not (_38598_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_38599_, _18789_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38600_, _38599_, _38598_);
  and (_38601_, _38298_, _38576_);
  and (_38602_, _38590_, _38572_);
  and (_38603_, _38602_, _38601_);
  and (_38604_, _38603_, _38600_);
  and (_38605_, _38593_, _18789_);
  and (_38606_, _38592_, _18789_);
  nor (_38607_, _38606_, _38605_);
  nor (_38608_, _38607_, _37017_);
  nor (_38609_, _38608_, _38604_);
  and (_38610_, _38609_, _38597_);
  nor (_38611_, _38610_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38612_, _38611_, _37006_);
  and (_38613_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_38614_, _38604_);
  not (_38615_, _38527_);
  and (_38616_, _38504_, _38615_);
  and (_38617_, _38616_, _38589_);
  and (_38618_, _38577_, _38056_);
  and (_38619_, _38618_, _37553_);
  and (_38620_, _38619_, _38617_);
  not (_38621_, _38620_);
  and (_38622_, _38527_, _38548_);
  and (_38623_, _38622_, _38588_);
  and (_38624_, _38623_, _37553_);
  and (_38625_, _38624_, _38331_);
  and (_38626_, _38320_, _37542_);
  and (_38627_, _38626_, _38617_);
  nor (_38628_, _38627_, _38625_);
  and (_38629_, _38628_, _38621_);
  not (_38630_, _38617_);
  nor (_38631_, _38298_, _38056_);
  and (_38632_, _38631_, _37803_);
  not (_38633_, _37803_);
  and (_38634_, _38601_, _38633_);
  and (_38635_, _38634_, _37542_);
  nor (_38636_, _38635_, _38632_);
  nor (_38637_, _38636_, _38630_);
  not (_38638_, _38637_);
  not (_38639_, _38504_);
  and (_38640_, _38573_, _38639_);
  and (_38641_, _38640_, _38632_);
  not (_38642_, _38641_);
  and (_38643_, _38631_, _38633_);
  and (_38644_, _38643_, _37553_);
  and (_38645_, _38644_, _38617_);
  and (_38646_, _38342_, _38571_);
  nor (_38647_, _38646_, _38645_);
  and (_38648_, _38647_, _38642_);
  and (_38649_, _38648_, _38638_);
  and (_38650_, _38578_, _37553_);
  and (_38651_, _38650_, _38617_);
  nor (_38652_, _37803_, _38309_);
  and (_38653_, _38652_, _38056_);
  and (_38654_, _38653_, _37553_);
  and (_38655_, _38654_, _38617_);
  nor (_38656_, _38655_, _38651_);
  and (_38657_, _38653_, _37542_);
  and (_38658_, _38657_, _38640_);
  and (_38659_, _38342_, _38640_);
  nor (_38660_, _38659_, _38658_);
  and (_38661_, _38660_, _38656_);
  and (_38662_, _38661_, _38649_);
  and (_38663_, _38662_, _38629_);
  and (_38664_, _38634_, _37553_);
  and (_38665_, _38664_, _38573_);
  not (_38666_, _38665_);
  and (_38667_, _38643_, _37542_);
  and (_38668_, _38667_, _38617_);
  and (_38669_, _38331_, _37542_);
  and (_38670_, _38602_, _38669_);
  nor (_38671_, _38670_, _38668_);
  and (_38672_, _38671_, _38666_);
  and (_38673_, _38579_, _38640_);
  and (_38674_, _38657_, _38617_);
  nor (_38675_, _38674_, _38673_);
  and (_38676_, _38675_, _38672_);
  and (_38677_, _38602_, _38342_);
  and (_38678_, _38664_, _38617_);
  nor (_38679_, _38678_, _38677_);
  and (_38680_, _38640_, _38669_);
  and (_38681_, _38654_, _38640_);
  nor (_38682_, _38681_, _38680_);
  and (_38683_, _38682_, _38679_);
  and (_38684_, _38683_, _38676_);
  and (_38685_, _38587_, _38640_);
  and (_38686_, _38573_, _38635_);
  nor (_38687_, _38686_, _38685_);
  and (_38688_, _38640_, _38583_);
  and (_38689_, _38587_, _38617_);
  nor (_38690_, _38689_, _38688_);
  and (_38691_, _38690_, _38687_);
  and (_38692_, _38632_, _37542_);
  and (_38693_, _38692_, _38602_);
  not (_38694_, _38693_);
  and (_38695_, _38632_, _37553_);
  and (_38696_, _38695_, _38602_);
  and (_38697_, _38602_, _38667_);
  nor (_38698_, _38697_, _38696_);
  and (_38699_, _38698_, _38694_);
  and (_38700_, _38602_, _38653_);
  and (_38701_, _38650_, _38573_);
  nor (_38702_, _38701_, _38700_);
  and (_38703_, _38702_, _38699_);
  and (_38704_, _38703_, _38691_);
  and (_38705_, _38704_, _38684_);
  and (_38706_, _38705_, _38663_);
  nor (_38707_, _38706_, _37039_);
  and (_38708_, \oc8051_top_1.oc8051_decoder1.state [0], _18789_);
  and (_38709_, _38708_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38710_, _38709_, _38641_);
  nor (_38711_, _38710_, _38707_);
  and (_38712_, _38711_, _38614_);
  nor (_38713_, _38712_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38714_, _38713_, _38613_);
  and (_38715_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38716_, _37553_, _38571_);
  and (_38717_, _38716_, _38622_);
  and (_38718_, _38717_, _38634_);
  and (_38719_, _38632_, _38623_);
  or (_38720_, _38719_, _38718_);
  and (_38721_, _38587_, _38623_);
  or (_38722_, _38721_, _38641_);
  and (_38723_, _38717_, _38331_);
  and (_38724_, _38643_, _38623_);
  nor (_38725_, _38724_, _38723_);
  not (_38726_, _38725_);
  or (_38727_, _38634_, _38618_);
  and (_38728_, _38727_, _38624_);
  or (_38729_, _38728_, _38726_);
  or (_38730_, _38729_, _38722_);
  or (_38731_, _38730_, _38720_);
  and (_38732_, _38602_, _38657_);
  and (_38733_, _38653_, _38623_);
  and (_38734_, _38583_, _38623_);
  nor (_38735_, _38734_, _38733_);
  not (_38736_, _38735_);
  and (_38737_, _38650_, _38623_);
  or (_38738_, _38737_, _38736_);
  nor (_38739_, _38738_, _38732_);
  nand (_38740_, _38739_, _38586_);
  nor (_38741_, _38740_, _38731_);
  nor (_38742_, _38741_, _37039_);
  and (_38743_, _38600_, _38578_);
  and (_38744_, _38743_, _38602_);
  or (_38745_, _38744_, _38710_);
  nor (_38746_, _38745_, _38742_);
  nor (_38747_, _38746_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38748_, _38747_, _38715_);
  nor (_38749_, _38748_, _38714_);
  and (_38750_, _38749_, _38612_);
  and (_09470_, _38750_, _43223_);
  and (_38751_, _31261_, _28282_);
  and (_38752_, _38751_, _27361_);
  and (_38753_, _28424_, _27953_);
  not (_38754_, _27821_);
  nor (_38755_, _38754_, _28128_);
  and (_38756_, _38755_, _38753_);
  and (_38757_, _38756_, _33188_);
  and (_38758_, _38757_, _38752_);
  not (_38759_, _38758_);
  and (_38760_, _38759_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_38761_, _24213_, _18855_);
  and (_38762_, _29817_, _24191_);
  nor (_38763_, _30940_, _38762_);
  and (_38764_, _38763_, _38761_);
  nor (_38765_, _31006_, _32241_);
  and (_38766_, _38765_, _38764_);
  nor (_38767_, _38766_, _20072_);
  not (_38768_, _38767_);
  and (_38769_, _38768_, _36637_);
  and (_38770_, _38769_, _36506_);
  nor (_38771_, _38770_, _38759_);
  nor (_38772_, _38771_, _38760_);
  and (_38773_, _38759_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38774_, _38766_, _21106_);
  not (_38775_, _38774_);
  and (_38776_, _38775_, _35898_);
  and (_38777_, _38776_, _35865_);
  and (_38778_, _38777_, _35767_);
  nor (_38779_, _38778_, _38759_);
  nor (_38780_, _38779_, _38773_);
  and (_38781_, _38759_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38782_, _38766_, _21280_);
  not (_38783_, _38782_);
  and (_38784_, _38783_, _35136_);
  and (_38785_, _38784_, _35103_);
  and (_38786_, _38785_, _35037_);
  nor (_38787_, _38786_, _38759_);
  nor (_38788_, _38787_, _38781_);
  and (_38789_, _38759_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38790_, _38766_, _21672_);
  not (_38791_, _38790_);
  and (_38792_, _38791_, _34472_);
  and (_38793_, _38792_, _34308_);
  nor (_38794_, _38793_, _38759_);
  nor (_38795_, _38794_, _38789_);
  and (_38796_, _38759_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38797_, _38766_, _22173_);
  not (_38798_, _38797_);
  and (_38799_, _38798_, _33623_);
  and (_38800_, _38799_, _33590_);
  and (_38801_, _38800_, _33427_);
  nor (_38802_, _38801_, _38759_);
  nor (_38803_, _38802_, _38796_);
  and (_38804_, _38759_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38805_, _38766_, _21998_);
  not (_38806_, _38805_);
  and (_38807_, _38806_, _32948_);
  and (_38808_, _38807_, _32796_);
  nor (_38809_, _38808_, _38759_);
  nor (_38810_, _38809_, _38804_);
  nor (_38811_, _38758_, _27547_);
  nor (_38812_, _38766_, _22542_);
  not (_38813_, _38812_);
  and (_38814_, _38813_, _32197_);
  and (_38815_, _38814_, _32164_);
  and (_38816_, _38815_, _32132_);
  not (_38817_, _38816_);
  and (_38818_, _38817_, _38758_);
  nor (_38819_, _38818_, _38811_);
  and (_38820_, _38819_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38821_, _38820_, _38810_);
  and (_38822_, _38821_, _38803_);
  and (_38823_, _38822_, _38795_);
  and (_38824_, _38823_, _38788_);
  and (_38825_, _38824_, _38780_);
  and (_38826_, _38825_, _38772_);
  nor (_38827_, _38758_, _27975_);
  nand (_38828_, _38827_, _38826_);
  or (_38829_, _38827_, _38826_);
  and (_38830_, _38829_, _27690_);
  and (_38831_, _38830_, _38828_);
  or (_38832_, _38758_, _28019_);
  or (_38833_, _38832_, _38831_);
  or (_38834_, _38766_, _20910_);
  and (_38835_, _38834_, _30930_);
  and (_38836_, _38835_, _30875_);
  and (_38837_, _38836_, _30570_);
  nand (_38838_, _38837_, _38758_);
  and (_38839_, _38838_, _38833_);
  and (_09491_, _38839_, _43223_);
  not (_38840_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38841_, _38819_, _38840_);
  nor (_38842_, _38819_, _38840_);
  nor (_38843_, _38842_, _38841_);
  and (_38844_, _38843_, _27690_);
  nor (_38845_, _38844_, _27558_);
  nor (_38846_, _38845_, _38758_);
  nor (_38847_, _38846_, _38818_);
  nand (_10647_, _38847_, _43223_);
  nor (_38848_, _38820_, _38810_);
  nor (_38849_, _38848_, _38821_);
  nor (_38850_, _38849_, _27097_);
  nor (_38851_, _38850_, _27393_);
  nor (_38852_, _38851_, _38758_);
  nor (_38853_, _38852_, _38809_);
  nand (_10658_, _38853_, _43223_);
  nor (_38854_, _38821_, _38803_);
  nor (_38855_, _38854_, _38822_);
  nor (_38856_, _38855_, _27097_);
  nor (_38857_, _38856_, _27152_);
  nor (_38858_, _38857_, _38758_);
  nor (_38859_, _38858_, _38802_);
  nand (_10669_, _38859_, _43223_);
  nor (_38860_, _38822_, _38795_);
  nor (_38861_, _38860_, _38823_);
  nor (_38862_, _38861_, _27097_);
  nor (_38863_, _38862_, _28216_);
  nor (_38864_, _38863_, _38758_);
  nor (_38865_, _38864_, _38794_);
  nor (_10680_, _38865_, rst);
  nor (_38866_, _38823_, _38788_);
  nor (_38867_, _38866_, _38824_);
  nor (_38868_, _38867_, _27097_);
  nor (_38869_, _38868_, _28348_);
  nor (_38870_, _38869_, _38758_);
  nor (_38871_, _38870_, _38787_);
  nor (_10691_, _38871_, rst);
  nor (_38872_, _38824_, _38780_);
  nor (_38873_, _38872_, _38825_);
  nor (_38874_, _38873_, _27097_);
  nor (_38875_, _38874_, _27865_);
  nor (_38876_, _38875_, _38758_);
  nor (_38877_, _38876_, _38779_);
  nor (_10702_, _38877_, rst);
  nor (_38878_, _38825_, _38772_);
  nor (_38879_, _38878_, _38826_);
  nor (_38880_, _38879_, _27097_);
  nor (_38881_, _38880_, _27723_);
  nor (_38882_, _38881_, _38758_);
  nor (_38883_, _38882_, _38771_);
  nor (_10713_, _38883_, rst);
  and (_38884_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18789_);
  and (_38885_, _38884_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_38886_, _38885_);
  nor (_38887_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38888_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38889_, _38888_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38890_, _38889_, _38887_);
  nor (_38891_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38892_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38893_, _38892_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38894_, _38893_, _38891_);
  nor (_38895_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38896_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38897_, _38896_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38898_, _38897_, _38895_);
  nor (_38899_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38900_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38901_, _38900_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38902_, _38901_, _38899_);
  nor (_38903_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38904_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38905_, _38904_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38906_, _38905_, _38903_);
  not (_38907_, _38906_);
  nor (_38908_, _38907_, _31347_);
  nor (_38909_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38910_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38911_, _38910_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38912_, _38911_, _38909_);
  and (_38913_, _38912_, _38908_);
  nor (_38914_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38915_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38916_, _38915_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38917_, _38916_, _38914_);
  and (_38918_, _38917_, _38913_);
  and (_38919_, _38918_, _38902_);
  nor (_38920_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38921_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38922_, _38921_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38923_, _38922_, _38920_);
  and (_38924_, _38923_, _38919_);
  and (_38925_, _38924_, _38898_);
  and (_38926_, _38925_, _38894_);
  or (_38927_, _38926_, _38890_);
  nand (_38928_, _38926_, _38890_);
  and (_38929_, _38928_, _38927_);
  and (_38930_, _38929_, _29828_);
  not (_38931_, _38930_);
  and (_38932_, _23905_, _18855_);
  and (_38933_, _30319_, _20930_);
  and (_38934_, _38933_, _28973_);
  and (_38935_, _38934_, _29006_);
  and (_38936_, _38935_, _29049_);
  and (_38937_, _38936_, _29641_);
  nor (_38938_, _38937_, _30341_);
  and (_38939_, _29543_, _19413_);
  nor (_38940_, _38939_, _38938_);
  and (_38941_, _30406_, _20910_);
  and (_38942_, _20246_, _19249_);
  and (_38943_, _20561_, _19576_);
  and (_38944_, _38943_, _38942_);
  and (_38945_, _38944_, _38941_);
  and (_38946_, _20398_, _19413_);
  and (_38947_, _38946_, _38945_);
  nor (_38948_, _38947_, _29543_);
  and (_38949_, _29543_, _20398_);
  nor (_38950_, _38949_, _38948_);
  and (_38951_, _38950_, _38940_);
  nor (_38952_, _29543_, _19762_);
  and (_38953_, _29543_, _19762_);
  nor (_38954_, _38953_, _38952_);
  and (_38955_, _38954_, _38951_);
  and (_38956_, _38955_, _30483_);
  nor (_38957_, _38955_, _30483_);
  nor (_38958_, _38957_, _38956_);
  and (_38959_, _38958_, _30254_);
  and (_38960_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_38961_, _29543_, _30483_);
  nor (_38962_, _38961_, _31435_);
  nor (_38963_, _38962_, _30537_);
  nor (_38964_, _31739_, _21672_);
  nor (_38965_, _30951_, _20745_);
  or (_38966_, _38965_, _38964_);
  or (_38967_, _38966_, _38963_);
  nor (_38968_, _38967_, _38960_);
  not (_38969_, _38968_);
  nor (_38970_, _38969_, _38959_);
  not (_38971_, _38970_);
  nor (_38972_, _38971_, _38932_);
  and (_38973_, _38972_, _38931_);
  nor (_38974_, _38973_, _38886_);
  and (_38975_, _38756_, _34690_);
  and (_38976_, _38975_, _38751_);
  or (_38977_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_38978_, _38977_, _38886_);
  nand (_38979_, _38976_, _31194_);
  and (_38980_, _38979_, _38978_);
  or (_38981_, _38980_, _38974_);
  and (_12664_, _38981_, _43223_);
  and (_38982_, _38751_, _33950_);
  and (_38983_, _38982_, _38756_);
  nor (_38984_, _38983_, _38885_);
  not (_38985_, _38984_);
  nand (_38986_, _38985_, _31194_);
  or (_38987_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38988_, _38987_, _43223_);
  and (_12685_, _38988_, _38986_);
  and (_38989_, _26507_, _24213_);
  not (_38990_, _38989_);
  and (_38991_, _38907_, _31347_);
  nor (_38992_, _38991_, _38908_);
  and (_38993_, _38992_, _29828_);
  nor (_38994_, _31435_, _30515_);
  not (_38995_, _38994_);
  nor (_38996_, _38995_, _30428_);
  nor (_38997_, _38996_, _28973_);
  and (_38998_, _38996_, _28973_);
  or (_38999_, _38998_, _33383_);
  nor (_39000_, _38999_, _38997_);
  nor (_39001_, _30951_, _19576_);
  and (_39002_, _23684_, _18855_);
  nor (_39003_, _31739_, _21280_);
  nor (_39004_, _30537_, _22542_);
  or (_39005_, _39004_, _39003_);
  or (_39006_, _39005_, _39002_);
  nor (_39007_, _39006_, _39001_);
  not (_39008_, _39007_);
  nor (_39009_, _39008_, _39000_);
  not (_39010_, _39009_);
  nor (_39011_, _39010_, _38993_);
  and (_39012_, _39011_, _38990_);
  nor (_39013_, _39012_, _38886_);
  or (_39014_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_39015_, _39014_, _38886_);
  nand (_39016_, _38976_, _32393_);
  and (_39017_, _39016_, _39015_);
  or (_39018_, _39017_, _39013_);
  and (_13600_, _39018_, _43223_);
  nor (_39019_, _38912_, _38908_);
  nor (_39020_, _39019_, _38913_);
  and (_39021_, _39020_, _29828_);
  not (_39022_, _39021_);
  and (_39023_, _25499_, _24213_);
  nor (_39024_, _20910_, _19576_);
  and (_39025_, _39024_, _30319_);
  and (_39026_, _39025_, _29543_);
  and (_39027_, _38941_, _19576_);
  and (_39028_, _39027_, _30341_);
  nor (_39029_, _39028_, _39026_);
  nor (_39030_, _39029_, _29006_);
  and (_39031_, _39029_, _29006_);
  nor (_39032_, _39031_, _39030_);
  nor (_39033_, _39032_, _33383_);
  nor (_39034_, _30951_, _20561_);
  and (_39035_, _23715_, _18855_);
  nor (_39036_, _31739_, _21106_);
  nor (_39037_, _30537_, _21998_);
  or (_39038_, _39037_, _39036_);
  or (_39039_, _39038_, _39035_);
  nor (_39040_, _39039_, _39034_);
  not (_39041_, _39040_);
  nor (_39042_, _39041_, _39033_);
  not (_39043_, _39042_);
  nor (_39044_, _39043_, _39023_);
  and (_39045_, _39044_, _39022_);
  nor (_39046_, _39045_, _38886_);
  or (_39047_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_39048_, _39047_, _38886_);
  nand (_39049_, _38976_, _33090_);
  and (_39050_, _39049_, _39048_);
  or (_39051_, _39050_, _39046_);
  and (_13611_, _39051_, _43223_);
  nor (_39052_, _38917_, _38913_);
  nor (_39053_, _39052_, _38918_);
  and (_39054_, _39053_, _29828_);
  not (_39055_, _39054_);
  and (_39056_, _39027_, _20561_);
  and (_39057_, _39056_, _30341_);
  and (_39058_, _39025_, _29006_);
  and (_39059_, _39058_, _29543_);
  nor (_39060_, _39059_, _39057_);
  and (_39061_, _39060_, _19249_);
  nor (_39062_, _39060_, _19249_);
  nor (_39063_, _39062_, _39061_);
  and (_39064_, _39063_, _30254_);
  not (_39065_, _39064_);
  nor (_39066_, _30537_, _22173_);
  and (_39067_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_39068_, _39067_, _39066_);
  and (_39069_, _23747_, _18855_);
  nor (_39070_, _31739_, _20072_);
  nor (_39071_, _30951_, _19249_);
  or (_39072_, _39071_, _39070_);
  nor (_39073_, _39072_, _39069_);
  and (_39074_, _39073_, _39068_);
  and (_39075_, _39074_, _39065_);
  and (_39076_, _39075_, _39055_);
  nor (_39077_, _39076_, _38886_);
  or (_39078_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_39079_, _39078_, _38886_);
  nand (_39080_, _38976_, _33809_);
  and (_39081_, _39080_, _39079_);
  or (_39082_, _39081_, _39077_);
  and (_13622_, _39082_, _43223_);
  nor (_39083_, _38918_, _38902_);
  not (_39084_, _39083_);
  nor (_39085_, _38919_, _31326_);
  and (_39086_, _39085_, _39084_);
  not (_39087_, _39086_);
  nor (_39088_, _38936_, _29641_);
  not (_39089_, _39088_);
  and (_39090_, _39089_, _38938_);
  and (_39091_, _39056_, _19249_);
  nor (_39092_, _39091_, _20246_);
  nor (_39093_, _39092_, _38945_);
  nor (_39094_, _39093_, _29543_);
  nor (_39095_, _39094_, _39090_);
  nor (_39096_, _39095_, _33383_);
  not (_39097_, _39096_);
  and (_39098_, _23779_, _18855_);
  nor (_39099_, _30951_, _20246_);
  nor (_39100_, _30537_, _21672_);
  and (_39101_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_39102_, _39101_, _39100_);
  or (_39103_, _39102_, _31740_);
  nor (_39104_, _39103_, _39099_);
  not (_39105_, _39104_);
  nor (_39106_, _39105_, _39098_);
  and (_39107_, _39106_, _39097_);
  and (_39108_, _39107_, _39087_);
  nor (_39109_, _39108_, _38886_);
  or (_39110_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_39111_, _39110_, _38886_);
  nand (_39112_, _38976_, _34591_);
  and (_39113_, _39112_, _39111_);
  or (_39114_, _39113_, _39109_);
  and (_13633_, _39114_, _43223_);
  nor (_39115_, _38923_, _38919_);
  nor (_39116_, _39115_, _38924_);
  and (_39117_, _39116_, _29828_);
  not (_39118_, _39117_);
  and (_39119_, _23810_, _18855_);
  nor (_39120_, _38945_, _29543_);
  nor (_39121_, _39120_, _38938_);
  nor (_39122_, _39121_, _28698_);
  and (_39123_, _39121_, _28698_);
  nor (_39124_, _39123_, _39122_);
  and (_39125_, _39124_, _30254_);
  and (_39126_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_39127_, _29543_, _21300_);
  or (_39128_, _39127_, _30537_);
  nor (_39129_, _39128_, _38939_);
  nor (_39130_, _31739_, _22542_);
  nor (_39131_, _30951_, _19413_);
  or (_39132_, _39131_, _39130_);
  or (_39133_, _39132_, _39129_);
  nor (_39134_, _39133_, _39126_);
  not (_39135_, _39134_);
  nor (_39136_, _39135_, _39125_);
  not (_39137_, _39136_);
  nor (_39138_, _39137_, _39119_);
  and (_39139_, _39138_, _39118_);
  nor (_39140_, _39139_, _38886_);
  or (_39141_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_39142_, _39141_, _38886_);
  nand (_39143_, _38976_, _35277_);
  and (_39144_, _39143_, _39142_);
  or (_39145_, _39144_, _39140_);
  and (_13644_, _39145_, _43223_);
  nor (_39146_, _38924_, _38898_);
  not (_39147_, _39146_);
  nor (_39148_, _38925_, _31326_);
  and (_39149_, _39148_, _39147_);
  not (_39150_, _39149_);
  and (_39151_, _23842_, _18855_);
  and (_39152_, _38945_, _19413_);
  nor (_39153_, _39152_, _29543_);
  not (_39154_, _39153_);
  and (_39155_, _39154_, _38940_);
  and (_39156_, _39155_, _20398_);
  nor (_39157_, _39155_, _20398_);
  nor (_39158_, _39157_, _39156_);
  nor (_39159_, _39158_, _33383_);
  or (_39160_, _38949_, _30537_);
  nor (_39161_, _39160_, _36420_);
  and (_39162_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_39163_, _31739_, _21998_);
  nor (_39164_, _30951_, _20398_);
  or (_39165_, _39164_, _39163_);
  nor (_39166_, _39165_, _39162_);
  not (_39167_, _39166_);
  nor (_39168_, _39167_, _39161_);
  not (_39169_, _39168_);
  nor (_39170_, _39169_, _39159_);
  not (_39171_, _39170_);
  nor (_39172_, _39171_, _39151_);
  and (_39173_, _39172_, _39150_);
  nor (_39174_, _39173_, _38886_);
  or (_39175_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_39176_, _39175_, _38886_);
  nand (_39177_, _38976_, _36083_);
  and (_39178_, _39177_, _39176_);
  or (_39179_, _39178_, _39174_);
  and (_13655_, _39179_, _43223_);
  nor (_39180_, _38925_, _38894_);
  not (_39181_, _39180_);
  nor (_39182_, _38926_, _31326_);
  and (_39183_, _39182_, _39181_);
  not (_39184_, _39183_);
  and (_39185_, _23874_, _18855_);
  and (_39186_, _38951_, _19762_);
  nor (_39187_, _38951_, _19762_);
  nor (_39188_, _39187_, _39186_);
  nor (_39189_, _39188_, _33383_);
  and (_39190_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_39191_, _29543_, _20083_);
  or (_39192_, _39191_, _30537_);
  nor (_39193_, _39192_, _38953_);
  nor (_39194_, _31739_, _22173_);
  nor (_39195_, _30951_, _19762_);
  or (_39196_, _39195_, _39194_);
  or (_39197_, _39196_, _39193_);
  nor (_39198_, _39197_, _39190_);
  not (_39199_, _39198_);
  nor (_39200_, _39199_, _39189_);
  not (_39201_, _39200_);
  nor (_39202_, _39201_, _39185_);
  and (_39203_, _39202_, _39184_);
  nor (_39204_, _39203_, _38886_);
  or (_39205_, _38976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_39206_, _39205_, _38886_);
  nand (_39207_, _38976_, _36811_);
  and (_39208_, _39207_, _39206_);
  or (_39209_, _39208_, _39204_);
  and (_13665_, _39209_, _43223_);
  nand (_39210_, _38985_, _32393_);
  or (_39211_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_39212_, _39211_, _43223_);
  and (_13676_, _39212_, _39210_);
  nand (_39213_, _38985_, _33090_);
  or (_39214_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_39215_, _39214_, _43223_);
  and (_13687_, _39215_, _39213_);
  nand (_39216_, _38985_, _33809_);
  or (_39217_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_39218_, _39217_, _43223_);
  and (_13698_, _39218_, _39216_);
  nand (_39219_, _38985_, _34591_);
  or (_39220_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_39221_, _39220_, _43223_);
  and (_13709_, _39221_, _39219_);
  nand (_39222_, _38985_, _35277_);
  or (_39223_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_39224_, _39223_, _43223_);
  and (_13720_, _39224_, _39222_);
  nand (_39225_, _38985_, _36083_);
  or (_39226_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_39227_, _39226_, _43223_);
  and (_13731_, _39227_, _39225_);
  nand (_39228_, _38985_, _36811_);
  or (_39229_, _38985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_39230_, _39229_, _43223_);
  and (_13742_, _39230_, _39228_);
  nor (_39231_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_39232_, _39231_, _31849_);
  and (_39233_, _39231_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not (_39234_, _27953_);
  nor (_39235_, _28424_, _39234_);
  nor (_39236_, _27821_, _28128_);
  and (_39237_, _38751_, _27624_);
  and (_39238_, _39237_, _39236_);
  and (_39239_, _39238_, _39235_);
  nor (_39240_, _39234_, _27821_);
  and (_39241_, _39240_, _31926_);
  and (_39242_, _39241_, _28446_);
  or (_39243_, _39242_, _39239_);
  or (_39244_, _39243_, _39233_);
  or (_39245_, _39244_, _39232_);
  and (_39246_, _39235_, _39236_);
  and (_39247_, _39246_, _39237_);
  nand (_39250_, _39247_, _38837_);
  and (_39252_, _39250_, _43223_);
  and (_39253_, _31882_, _32481_);
  not (_39254_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_39255_, _31882_, _39254_);
  nand (_39256_, _39255_, _39242_);
  or (_39257_, _39256_, _39253_);
  and (_39258_, _39257_, _39252_);
  and (_15145_, _39258_, _39245_);
  not (_39259_, _39247_);
  not (_39260_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_39262_, _39240_, _28446_);
  and (_39271_, _39262_, _31926_);
  nand (_39277_, _39271_, _33199_);
  nand (_39283_, _39277_, _39260_);
  and (_39286_, _39283_, _39259_);
  or (_39287_, _39277_, _32481_);
  and (_39288_, _39287_, _39286_);
  nor (_39289_, _39259_, _38808_);
  or (_39290_, _39289_, _39288_);
  and (_17326_, _39290_, _43223_);
  or (_39291_, _31390_, _29740_);
  not (_39292_, _31370_);
  nand (_39293_, _39292_, _29740_);
  and (_39294_, _39293_, _28534_);
  and (_39295_, _39294_, _39291_);
  not (_39296_, _28556_);
  nand (_39297_, _30188_, _39296_);
  or (_39298_, _30188_, _28567_);
  and (_39299_, _29828_, _39298_);
  and (_39300_, _39299_, _39297_);
  and (_39301_, _38946_, _25400_);
  and (_39302_, _38944_, _24213_);
  nand (_39303_, _39302_, _39301_);
  nand (_39304_, _39303_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_39305_, _39304_, _39300_);
  or (_39306_, _39305_, _39295_);
  or (_39307_, _23978_, _23937_);
  or (_39308_, _39307_, _24000_);
  or (_39309_, _39308_, _24043_);
  or (_39312_, _39309_, _24074_);
  or (_39313_, _39312_, _24117_);
  or (_39314_, _39313_, _24148_);
  and (_39315_, _39314_, _18855_);
  or (_39316_, _39315_, _39306_);
  or (_39317_, _39316_, _28501_);
  nor (_39318_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_39319_, _39318_, _39242_);
  and (_39320_, _39319_, _39317_);
  and (_39321_, _33961_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_39322_, _39321_, _33972_);
  and (_39323_, _39322_, _39271_);
  or (_39324_, _39323_, _39247_);
  or (_39325_, _39324_, _39320_);
  nand (_39326_, _39247_, _38801_);
  and (_39327_, _39326_, _43223_);
  and (_17337_, _39327_, _39325_);
  not (_39328_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_39329_, _39271_, _34690_);
  nand (_39330_, _39329_, _39328_);
  or (_39331_, _39329_, _32481_);
  and (_39332_, _39331_, _39330_);
  and (_39333_, _39332_, _39259_);
  nor (_39334_, _39259_, _38793_);
  or (_39335_, _39334_, _39333_);
  and (_17348_, _39335_, _43223_);
  and (_39336_, _35386_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_39337_, _39336_, _35430_);
  and (_39338_, _39242_, _43223_);
  and (_39339_, _39338_, _39337_);
  and (_39340_, _39259_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_39341_, _39259_, _38786_);
  nor (_39342_, _39341_, _39340_);
  nor (_39348_, _39342_, rst);
  not (_39343_, _39242_);
  or (_39344_, _39343_, _35397_);
  and (_39345_, _39344_, _39348_);
  or (_17359_, _39345_, _39339_);
  not (_39347_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand (_39351_, _39271_, _36171_);
  nand (_39357_, _39351_, _39347_);
  and (_39362_, _39357_, _39259_);
  or (_39369_, _39351_, _32481_);
  and (_39377_, _39369_, _39362_);
  nor (_39385_, _39259_, _38778_);
  or (_39386_, _39385_, _39377_);
  and (_17370_, _39386_, _43223_);
  not (_39387_, _36909_);
  nor (_39388_, _39387_, _31849_);
  or (_39389_, _36909_, _34319_);
  nand (_39390_, _39389_, _39242_);
  or (_39391_, _39390_, _39388_);
  nand (_39392_, _39247_, _38770_);
  and (_39393_, _39392_, _43223_);
  and (_39394_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_39395_, _29828_, _30090_);
  and (_39396_, _29696_, _28534_);
  or (_39397_, _39396_, _39395_);
  and (_39398_, _39397_, _39394_);
  nand (_39399_, _39394_, _30951_);
  and (_39400_, _39399_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_39401_, _39400_, _39243_);
  or (_39402_, _39401_, _39398_);
  and (_39403_, _39402_, _39393_);
  and (_17381_, _39403_, _39391_);
  not (_39404_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39405_, _38884_, _39404_);
  not (_39406_, _39405_);
  nor (_39407_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_39408_, _39407_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39409_, _27624_, _28282_);
  and (_39410_, _28424_, _39234_);
  and (_39411_, _39410_, _39236_);
  and (_39412_, _39411_, _39409_);
  and (_39413_, _39412_, _31261_);
  nor (_39414_, _39413_, _39408_);
  nor (_39415_, _39414_, _31194_);
  and (_39416_, _28424_, _28282_);
  not (_39417_, _31926_);
  nor (_39418_, _39417_, _28128_);
  and (_39419_, _39418_, _27964_);
  and (_39420_, _39419_, _39416_);
  and (_39426_, _39420_, _31882_);
  and (_39437_, _39426_, _31849_);
  nor (_39438_, _39426_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_39439_, _39438_);
  and (_39440_, _39414_, _39406_);
  and (_39451_, _39440_, _39439_);
  not (_39457_, _39451_);
  nor (_39458_, _39457_, _39437_);
  or (_39459_, _39458_, _39415_);
  and (_39460_, _39459_, _39406_);
  nor (_39461_, _39406_, _38973_);
  or (_39462_, _39461_, _39460_);
  and (_17950_, _39462_, _43223_);
  nor (_39463_, _39406_, _39012_);
  nor (_39464_, _39414_, _32404_);
  not (_39465_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_39466_, _39416_, _28139_);
  and (_39467_, _31926_, _27964_);
  and (_39468_, _39467_, _39466_);
  nor (_39469_, _39468_, _39465_);
  not (_39470_, _39469_);
  and (_39471_, _39470_, _39414_);
  not (_39472_, _39471_);
  and (_39473_, _32481_, _27624_);
  nor (_39474_, _27624_, _39465_);
  nor (_39475_, _39474_, _39473_);
  and (_39476_, _39440_, _39468_);
  not (_39477_, _39476_);
  nor (_39478_, _39477_, _39475_);
  nor (_39479_, _39478_, _39472_);
  nor (_39480_, _39479_, _39405_);
  not (_39481_, _39480_);
  nor (_39482_, _39481_, _39464_);
  nor (_39483_, _39482_, _39463_);
  nor (_19739_, _39483_, rst);
  and (_39484_, _39405_, _39045_);
  nor (_39485_, _39414_, _33090_);
  and (_39486_, _39420_, _33199_);
  and (_39487_, _39486_, _31849_);
  nor (_39488_, _39486_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not (_39489_, _39488_);
  and (_39490_, _39489_, _39440_);
  not (_39491_, _39490_);
  nor (_39492_, _39491_, _39487_);
  nor (_39493_, _39492_, _39405_);
  not (_39494_, _39493_);
  nor (_39495_, _39494_, _39485_);
  nor (_39496_, _39495_, _39484_);
  and (_19751_, _39496_, _43223_);
  nor (_39497_, _39414_, _33809_);
  and (_39498_, _39420_, _33950_);
  and (_39499_, _39498_, _31849_);
  nor (_39500_, _39498_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_39501_, _39500_);
  and (_39502_, _39501_, _39440_);
  not (_39503_, _39502_);
  nor (_39504_, _39503_, _39499_);
  or (_39505_, _39504_, _39497_);
  and (_39506_, _39505_, _39406_);
  nor (_39507_, _39406_, _39076_);
  or (_39508_, _39507_, _39506_);
  and (_19763_, _39508_, _43223_);
  nor (_39509_, _39414_, _34591_);
  not (_39510_, _39420_);
  and (_39511_, _39440_, _39510_);
  and (_39512_, _39511_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  not (_39513_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39514_, _34690_, _39513_);
  nor (_39515_, _39514_, _34700_);
  nor (_39516_, _39515_, _39477_);
  nor (_39517_, _39516_, _39512_);
  and (_39518_, _39517_, _39406_);
  not (_39519_, _39518_);
  nor (_39520_, _39519_, _39509_);
  and (_39521_, _39405_, _39108_);
  or (_39522_, _39521_, _39520_);
  nor (_19775_, _39522_, rst);
  nor (_39523_, _39414_, _35277_);
  and (_39524_, _39420_, _35375_);
  and (_39525_, _39524_, _31849_);
  nor (_39526_, _39524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_39527_, _39526_);
  and (_39528_, _39527_, _39440_);
  not (_39529_, _39528_);
  nor (_39530_, _39529_, _39525_);
  or (_39531_, _39530_, _39523_);
  and (_39532_, _39531_, _39406_);
  nor (_39533_, _39406_, _39139_);
  or (_39534_, _39533_, _39532_);
  and (_19787_, _39534_, _43223_);
  nor (_39535_, _39414_, _36083_);
  and (_39536_, _39420_, _36171_);
  and (_39537_, _39536_, _31849_);
  nor (_39538_, _39536_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_39539_, _39538_);
  and (_39540_, _39539_, _39440_);
  not (_39541_, _39540_);
  nor (_39542_, _39541_, _39537_);
  or (_39543_, _39542_, _39535_);
  and (_39544_, _39543_, _39406_);
  nor (_39545_, _39406_, _39173_);
  or (_39546_, _39545_, _39544_);
  and (_19798_, _39546_, _43223_);
  nor (_39547_, _39414_, _36811_);
  and (_39548_, _39511_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_39549_, _39387_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_39550_, _39549_, _39388_);
  nor (_39551_, _39550_, _39477_);
  nor (_39552_, _39551_, _39548_);
  and (_39553_, _39552_, _39406_);
  not (_39554_, _39553_);
  nor (_39555_, _39554_, _39547_);
  and (_39556_, _39405_, _39203_);
  or (_39557_, _39556_, _39555_);
  nor (_19810_, _39557_, rst);
  and (_39558_, _27953_, _27821_);
  and (_39559_, _39466_, _39558_);
  and (_39560_, _39559_, _31882_);
  nand (_39561_, _39560_, _31849_);
  or (_39562_, _39560_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39563_, _39562_, _31926_);
  and (_39564_, _39563_, _39561_);
  and (_39565_, _38756_, _39409_);
  nand (_39566_, _39565_, _38837_);
  or (_39567_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39568_, _39567_, _31261_);
  and (_39569_, _39568_, _39566_);
  not (_39570_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_39571_, _31260_, _39570_);
  or (_39572_, _39571_, rst);
  or (_39573_, _39572_, _39569_);
  or (_31017_, _39573_, _39564_);
  and (_39574_, _39558_, _28446_);
  and (_39575_, _39574_, _31882_);
  nand (_39576_, _39575_, _31849_);
  or (_39577_, _39575_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39578_, _39577_, _31926_);
  and (_39579_, _39578_, _39576_);
  and (_39580_, _39235_, _38755_);
  and (_39581_, _39580_, _39409_);
  nand (_39582_, _39581_, _38837_);
  or (_39583_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39584_, _39583_, _31261_);
  and (_39585_, _39584_, _39582_);
  not (_39586_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_39587_, _31260_, _39586_);
  or (_39588_, _39587_, rst);
  or (_39589_, _39588_, _39585_);
  or (_31040_, _39589_, _39579_);
  and (_39590_, _39234_, _27821_);
  and (_39591_, _39590_, _39466_);
  and (_39592_, _39591_, _31882_);
  nand (_39593_, _39592_, _31849_);
  or (_39594_, _39592_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39595_, _39594_, _31926_);
  and (_39596_, _39595_, _39593_);
  and (_39597_, _39410_, _38755_);
  and (_39598_, _39597_, _39409_);
  not (_39599_, _39598_);
  nor (_39600_, _39599_, _38837_);
  not (_39601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_39602_, _39598_, _39601_);
  or (_39603_, _39602_, _39600_);
  and (_39604_, _39603_, _31261_);
  nor (_39605_, _31260_, _39601_);
  or (_39606_, _39605_, rst);
  or (_39607_, _39606_, _39604_);
  or (_31062_, _39607_, _39596_);
  and (_39608_, _39590_, _28446_);
  nand (_39609_, _39608_, _31882_);
  or (_39610_, _39609_, _32481_);
  not (_39611_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nand (_39612_, _39609_, _39611_);
  and (_39613_, _39612_, _31926_);
  and (_39614_, _39613_, _39610_);
  nor (_39615_, _28424_, _27953_);
  and (_39616_, _38755_, _39615_);
  and (_39617_, _39616_, _39409_);
  not (_39618_, _39617_);
  nor (_39619_, _39618_, _38837_);
  nor (_39620_, _39617_, _39611_);
  or (_39621_, _39620_, _39619_);
  and (_39622_, _39621_, _31261_);
  nor (_39623_, _31260_, _39611_);
  or (_39624_, _39623_, rst);
  or (_39625_, _39624_, _39622_);
  or (_31085_, _39625_, _39614_);
  or (_39626_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_39627_, _39626_, _31926_);
  and (_39628_, _39559_, _27624_);
  nand (_39629_, _39628_, _31849_);
  and (_39630_, _39629_, _39627_);
  nand (_39631_, _39565_, _38816_);
  and (_39632_, _39631_, _31261_);
  and (_39641_, _39632_, _39626_);
  not (_39652_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39663_, _31260_, _39652_);
  or (_39672_, _39663_, rst);
  or (_39678_, _39672_, _39641_);
  or (_40913_, _39678_, _39630_);
  and (_39699_, _33199_, _28282_);
  and (_39710_, _39699_, _38756_);
  nand (_39721_, _39710_, _31849_);
  or (_39732_, _39710_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39743_, _39732_, _31926_);
  and (_39754_, _39743_, _39721_);
  nand (_39765_, _39565_, _38808_);
  or (_39776_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39787_, _39776_, _31261_);
  and (_39798_, _39787_, _39765_);
  not (_39809_, _31260_);
  and (_39820_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39831_, _39820_, rst);
  or (_39842_, _39831_, _39798_);
  or (_40915_, _39842_, _39754_);
  not (_39846_, _34711_);
  nand (_39847_, _39559_, _39846_);
  and (_39848_, _39847_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39849_, _33983_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39850_, _39849_, _33972_);
  and (_39851_, _39850_, _39559_);
  or (_39852_, _39851_, _39848_);
  and (_39853_, _39852_, _31926_);
  nand (_39854_, _39565_, _38801_);
  or (_39855_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39856_, _39855_, _31261_);
  and (_39857_, _39856_, _39854_);
  and (_39858_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39859_, _39858_, rst);
  or (_39860_, _39859_, _39857_);
  or (_40917_, _39860_, _39853_);
  nand (_39861_, _39559_, _27361_);
  and (_39862_, _39861_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39863_, _39846_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39864_, _39863_, _34700_);
  and (_39865_, _39864_, _39559_);
  or (_39866_, _39865_, _39862_);
  and (_39867_, _39866_, _31926_);
  nand (_39868_, _39565_, _38793_);
  or (_39869_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39870_, _39869_, _31261_);
  and (_39871_, _39870_, _39868_);
  and (_39872_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39873_, _39872_, rst);
  or (_39874_, _39873_, _39871_);
  or (_40919_, _39874_, _39867_);
  not (_39875_, _39559_);
  or (_39876_, _39875_, _35397_);
  and (_39877_, _39876_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39878_, _35386_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39879_, _39878_, _35430_);
  and (_39880_, _39879_, _39559_);
  or (_39881_, _39880_, _39877_);
  and (_39882_, _39881_, _31926_);
  nand (_39883_, _39565_, _38786_);
  or (_39884_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39885_, _39884_, _31261_);
  and (_39886_, _39885_, _39883_);
  and (_39887_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39888_, _39887_, rst);
  or (_39889_, _39888_, _39886_);
  or (_40921_, _39889_, _39882_);
  and (_39890_, _39559_, _36171_);
  nand (_39891_, _39890_, _31849_);
  or (_39892_, _39890_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39893_, _39892_, _31926_);
  and (_39894_, _39893_, _39891_);
  nand (_39895_, _39565_, _38778_);
  or (_39896_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39897_, _39896_, _31261_);
  and (_39898_, _39897_, _39895_);
  and (_39899_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39900_, _39899_, rst);
  or (_39901_, _39900_, _39898_);
  or (_40923_, _39901_, _39894_);
  and (_39902_, _39559_, _36909_);
  nand (_39903_, _39902_, _31849_);
  or (_39904_, _39902_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39905_, _39904_, _31926_);
  and (_39906_, _39905_, _39903_);
  nand (_39907_, _39565_, _38770_);
  or (_39908_, _39565_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39909_, _39908_, _31261_);
  and (_39910_, _39909_, _39907_);
  and (_39911_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39912_, _39911_, rst);
  or (_39913_, _39912_, _39910_);
  or (_40925_, _39913_, _39906_);
  and (_39914_, _39574_, _27624_);
  nand (_39915_, _39914_, _31849_);
  or (_39916_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39917_, _39916_, _31926_);
  and (_39918_, _39917_, _39915_);
  nand (_39919_, _39581_, _38816_);
  and (_39920_, _39919_, _31261_);
  and (_39921_, _39920_, _39916_);
  not (_39922_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39923_, _31260_, _39922_);
  or (_39924_, _39923_, rst);
  or (_39925_, _39924_, _39921_);
  or (_40927_, _39925_, _39918_);
  and (_39926_, _39574_, _33199_);
  nand (_39927_, _39926_, _31849_);
  or (_39928_, _39926_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39929_, _39928_, _31926_);
  and (_39930_, _39929_, _39927_);
  nand (_39931_, _39581_, _38808_);
  or (_39932_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39933_, _39932_, _31261_);
  and (_39934_, _39933_, _39931_);
  and (_39935_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39936_, _39935_, rst);
  or (_39937_, _39936_, _39934_);
  or (_40929_, _39937_, _39930_);
  and (_39938_, _39574_, _33950_);
  nand (_39939_, _39938_, _31849_);
  or (_39940_, _39938_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39941_, _39940_, _31926_);
  and (_39942_, _39941_, _39939_);
  nand (_39943_, _39581_, _38801_);
  or (_39944_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39945_, _39944_, _31261_);
  and (_39946_, _39945_, _39943_);
  and (_39947_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39948_, _39947_, rst);
  or (_39949_, _39948_, _39946_);
  or (_40931_, _39949_, _39942_);
  and (_39950_, _39574_, _34690_);
  nand (_39951_, _39950_, _31849_);
  or (_39952_, _39950_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39953_, _39952_, _31926_);
  and (_39954_, _39953_, _39951_);
  nand (_39955_, _39581_, _38793_);
  or (_39956_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39957_, _39956_, _31261_);
  and (_39958_, _39957_, _39955_);
  and (_39959_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39960_, _39959_, rst);
  or (_39961_, _39960_, _39958_);
  or (_40933_, _39961_, _39954_);
  and (_39962_, _39574_, _35375_);
  nand (_39963_, _39962_, _31849_);
  or (_39964_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39965_, _39964_, _31926_);
  and (_39966_, _39965_, _39963_);
  nand (_39967_, _39581_, _38786_);
  or (_39968_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39969_, _39968_, _31261_);
  and (_39970_, _39969_, _39967_);
  and (_39971_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39972_, _39971_, rst);
  or (_39973_, _39972_, _39970_);
  or (_40935_, _39973_, _39966_);
  and (_39974_, _39574_, _36171_);
  nand (_39975_, _39974_, _31849_);
  or (_39976_, _39974_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39977_, _39976_, _31926_);
  and (_39978_, _39977_, _39975_);
  nand (_39979_, _39581_, _38778_);
  or (_39980_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39981_, _39980_, _31261_);
  and (_39982_, _39981_, _39979_);
  and (_39983_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39984_, _39983_, rst);
  or (_39985_, _39984_, _39982_);
  or (_40937_, _39985_, _39978_);
  and (_39986_, _39574_, _36909_);
  nand (_39987_, _39986_, _31849_);
  or (_39988_, _39986_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39989_, _39988_, _31926_);
  and (_39990_, _39989_, _39987_);
  nand (_39991_, _39581_, _38770_);
  or (_39992_, _39581_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39993_, _39992_, _31261_);
  and (_39994_, _39993_, _39991_);
  and (_39995_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39996_, _39995_, rst);
  or (_39997_, _39996_, _39994_);
  or (_40938_, _39997_, _39990_);
  nand (_39998_, _39598_, _31849_);
  or (_39999_, _39598_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_40000_, _39999_, _31926_);
  and (_40001_, _40000_, _39998_);
  nand (_40002_, _39598_, _38816_);
  and (_40003_, _40002_, _31261_);
  and (_40004_, _40003_, _39999_);
  not (_40005_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_40006_, _31260_, _40005_);
  or (_40007_, _40006_, rst);
  or (_40008_, _40007_, _40004_);
  or (_40940_, _40008_, _40001_);
  and (_40009_, _39591_, _33199_);
  nand (_40010_, _40009_, _31849_);
  or (_40011_, _40009_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_40012_, _40011_, _31926_);
  and (_40013_, _40012_, _40010_);
  nor (_40014_, _39599_, _38808_);
  and (_40015_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_40016_, _40015_, _40014_);
  and (_40017_, _40016_, _31261_);
  and (_40018_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_40019_, _40018_, rst);
  or (_40020_, _40019_, _40017_);
  or (_40942_, _40020_, _40013_);
  and (_40021_, _39591_, _33950_);
  nand (_40022_, _40021_, _31849_);
  or (_40023_, _40021_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_40024_, _40023_, _31926_);
  and (_40025_, _40024_, _40022_);
  nor (_40026_, _39599_, _38801_);
  and (_40027_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_40028_, _40027_, _40026_);
  and (_40029_, _40028_, _31261_);
  and (_40030_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_40031_, _40030_, rst);
  or (_40032_, _40031_, _40029_);
  or (_40944_, _40032_, _40025_);
  and (_40033_, _39591_, _34690_);
  nand (_40034_, _40033_, _31849_);
  or (_40035_, _40033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_40036_, _40035_, _31926_);
  and (_40037_, _40036_, _40034_);
  nor (_40038_, _39599_, _38793_);
  and (_40039_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_40040_, _40039_, _40038_);
  and (_40041_, _40040_, _31261_);
  and (_40042_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_40043_, _40042_, rst);
  or (_40044_, _40043_, _40041_);
  or (_40946_, _40044_, _40037_);
  and (_40045_, _39591_, _35375_);
  nand (_40046_, _40045_, _31849_);
  or (_40047_, _40045_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_40048_, _40047_, _31926_);
  and (_40049_, _40048_, _40046_);
  nor (_40050_, _39599_, _38786_);
  and (_40051_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_40052_, _40051_, _40050_);
  and (_40053_, _40052_, _31261_);
  and (_40054_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_40055_, _40054_, rst);
  or (_40056_, _40055_, _40053_);
  or (_40948_, _40056_, _40049_);
  and (_40057_, _39591_, _36171_);
  nand (_40058_, _40057_, _31849_);
  or (_40059_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_40060_, _40059_, _31926_);
  and (_40061_, _40060_, _40058_);
  nor (_40062_, _39599_, _38778_);
  and (_40067_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_40073_, _40067_, _40062_);
  and (_40074_, _40073_, _31261_);
  and (_40075_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_40076_, _40075_, rst);
  or (_40077_, _40076_, _40074_);
  or (_40950_, _40077_, _40061_);
  and (_40078_, _39591_, _36909_);
  nand (_40079_, _40078_, _31849_);
  or (_40080_, _40078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_40081_, _40080_, _31926_);
  and (_40082_, _40081_, _40079_);
  nor (_40083_, _39599_, _38770_);
  and (_40084_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_40085_, _40084_, _40083_);
  and (_40086_, _40085_, _31261_);
  and (_40087_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_40088_, _40087_, rst);
  or (_40089_, _40088_, _40086_);
  or (_40952_, _40089_, _40082_);
  and (_40090_, _39608_, _27624_);
  nand (_40091_, _40090_, _31849_);
  or (_40092_, _39617_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_40093_, _40092_, _31926_);
  and (_40094_, _40093_, _40091_);
  nand (_40095_, _39617_, _38816_);
  and (_40096_, _40095_, _31261_);
  and (_40097_, _40096_, _40092_);
  not (_40098_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_40099_, _31260_, _40098_);
  or (_40100_, _40099_, rst);
  or (_40101_, _40100_, _40097_);
  or (_40954_, _40101_, _40094_);
  and (_40102_, _39608_, _33199_);
  nand (_40103_, _40102_, _31849_);
  or (_40104_, _40102_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_40105_, _40104_, _31926_);
  and (_40106_, _40105_, _40103_);
  nor (_40107_, _39618_, _38808_);
  and (_40108_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_40109_, _40108_, _40107_);
  and (_40110_, _40109_, _31261_);
  and (_40111_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_40112_, _40111_, rst);
  or (_40113_, _40112_, _40110_);
  or (_40956_, _40113_, _40106_);
  and (_40114_, _39608_, _33950_);
  nand (_40115_, _40114_, _31849_);
  or (_40116_, _40114_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_40117_, _40116_, _31926_);
  and (_40118_, _40117_, _40115_);
  nor (_40119_, _39618_, _38801_);
  and (_40120_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_40121_, _40120_, _40119_);
  and (_40122_, _40121_, _31261_);
  and (_40123_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_40124_, _40123_, rst);
  or (_40125_, _40124_, _40122_);
  or (_40958_, _40125_, _40118_);
  and (_40126_, _39608_, _34690_);
  nand (_40127_, _40126_, _31849_);
  or (_40128_, _40126_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_40129_, _40128_, _31926_);
  and (_40130_, _40129_, _40127_);
  nor (_40131_, _39618_, _38793_);
  and (_40132_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_40133_, _40132_, _40131_);
  and (_40134_, _40133_, _31261_);
  and (_40135_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_40136_, _40135_, rst);
  or (_40137_, _40136_, _40134_);
  or (_40960_, _40137_, _40130_);
  and (_40138_, _39608_, _35375_);
  nand (_40139_, _40138_, _31849_);
  or (_40140_, _40138_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_40141_, _40140_, _31926_);
  and (_40142_, _40141_, _40139_);
  nor (_40143_, _39618_, _38786_);
  and (_40144_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_40145_, _40144_, _40143_);
  and (_40146_, _40145_, _31261_);
  and (_40147_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_40148_, _40147_, rst);
  or (_40149_, _40148_, _40146_);
  or (_40962_, _40149_, _40142_);
  and (_40150_, _39608_, _36171_);
  nand (_40151_, _40150_, _31849_);
  or (_40152_, _40150_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_40153_, _40152_, _31926_);
  and (_40154_, _40153_, _40151_);
  nor (_40155_, _39618_, _38778_);
  and (_40156_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_40157_, _40156_, _40155_);
  and (_40158_, _40157_, _31261_);
  and (_40159_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_40160_, _40159_, rst);
  or (_40161_, _40160_, _40158_);
  or (_40963_, _40161_, _40154_);
  and (_40172_, _39608_, _36909_);
  nand (_40183_, _40172_, _31849_);
  or (_40194_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_40205_, _40194_, _31926_);
  and (_40216_, _40205_, _40183_);
  nor (_40223_, _39618_, _38770_);
  and (_40224_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_40225_, _40224_, _40223_);
  and (_40226_, _40225_, _31261_);
  and (_40227_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_40228_, _40227_, rst);
  or (_40229_, _40228_, _40226_);
  or (_40965_, _40229_, _40216_);
  and (_41415_, t0_i, _43223_);
  and (_41418_, t1_i, _43223_);
  not (_40230_, _31261_);
  nor (_40231_, _40230_, _28282_);
  and (_40232_, _40231_, _34690_);
  and (_40233_, _40232_, _38756_);
  nand (_40234_, _40233_, _38837_);
  nor (_40235_, _27361_, _28282_);
  and (_40236_, _40235_, _38757_);
  and (_40237_, _40236_, _31261_);
  not (_40238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40239_, _40238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_40240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40241_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _40240_);
  nor (_40242_, _40241_, _40239_);
  or (_40243_, _40242_, _40237_);
  and (_40244_, _40243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_40245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_40246_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_40247_, t1_i);
  and (_40248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40247_);
  nor (_40249_, _40248_, _40246_);
  not (_40250_, _40249_);
  not (_40251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_40252_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _40251_);
  nor (_40253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_40254_, _40253_);
  and (_40255_, _40254_, _40252_);
  and (_40256_, _40255_, _40250_);
  not (_40257_, _40256_);
  nand (_40258_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_40259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_40260_, _40259_, _40258_);
  nor (_40261_, _40260_, _40257_);
  and (_40262_, _40261_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_40263_, _40262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand (_40264_, _40263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_40265_, _40264_, _40245_);
  not (_40266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_40267_, _40260_, _40266_);
  and (_40268_, _40267_, _40256_);
  and (_40269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_40270_, _40269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_40271_, _40270_, _40268_);
  nor (_40272_, _40271_, _40242_);
  and (_40273_, _40272_, _40265_);
  and (_40274_, _40271_, _40239_);
  and (_40275_, _40274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40276_, _40275_, _40273_);
  nor (_40277_, _40276_, _40237_);
  or (_40278_, _40277_, _40244_);
  or (_40279_, _40233_, _40278_);
  and (_40280_, _40279_, _43223_);
  and (_41421_, _40280_, _40234_);
  nand (_40281_, _40237_, _38837_);
  and (_40282_, _40231_, _38975_);
  not (_40284_, _40282_);
  and (_40290_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40291_, _40290_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40292_, _40270_, _40267_);
  and (_40293_, _40292_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_40294_, _40293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_40295_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40296_, _40295_, _40256_);
  and (_40297_, _40296_, _40291_);
  and (_40298_, _40297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40299_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40300_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40301_, _40300_, _40299_);
  and (_40302_, _40301_, _40241_);
  and (_40303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_40304_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_40305_, _40304_, _40267_);
  and (_40306_, _40305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40307_, _40306_, _40256_);
  and (_40308_, _40307_, _40291_);
  and (_40309_, _40308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40310_, _40309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_40311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_40312_, _40309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_40313_, _40312_, _40311_);
  nor (_40314_, _40313_, _40310_);
  or (_40315_, _40314_, _40303_);
  or (_40316_, _40315_, _40302_);
  or (_40317_, _40316_, _40237_);
  and (_40318_, _40317_, _40284_);
  and (_40319_, _40318_, _40281_);
  and (_40320_, _40282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_40321_, _40320_, _40319_);
  and (_41424_, _40321_, _43223_);
  and (_40322_, _40257_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_40323_, _40322_, _40299_);
  and (_40324_, _40323_, _40241_);
  or (_40325_, _40322_, _40310_);
  and (_40326_, _40325_, _40311_);
  nand (_40327_, _40256_, _40238_);
  and (_40328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_40329_, _40328_, _40327_);
  or (_40330_, _40329_, _40274_);
  or (_40331_, _40330_, _40326_);
  or (_40332_, _40331_, _40324_);
  nor (_40333_, _40233_, rst);
  nand (_40334_, _40333_, _40332_);
  nor (_41427_, _40334_, _40237_);
  and (_40335_, _40231_, _35375_);
  and (_40336_, _40335_, _38756_);
  nor (_40337_, _40336_, rst);
  not (_40338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_40339_, t0_i);
  and (_40340_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40339_);
  nor (_40341_, _40340_, _40338_);
  not (_40342_, _40341_);
  not (_40343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_40344_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_40345_, _40344_, _40343_);
  and (_40346_, _40345_, _40342_);
  not (_40347_, _40346_);
  and (_40348_, _40347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_40349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40350_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_40351_, _40350_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_40352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_40353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40354_, _40353_, _40352_);
  and (_40355_, _40354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_40356_, _40355_, _40346_);
  and (_40357_, _40356_, _40351_);
  and (_40358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40360_, _40359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40361_, _40360_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40362_, _40361_, _40358_);
  and (_40363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_40364_, _40363_, _40362_);
  or (_40365_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40366_, _40365_, _40357_);
  nor (_40367_, _40366_, _40349_);
  not (_40368_, _40349_);
  and (_40372_, _40362_, _40356_);
  and (_40380_, _40372_, _40363_);
  nor (_40381_, _40380_, _40368_);
  nor (_40382_, _40381_, _40367_);
  nor (_40383_, _40382_, _40348_);
  and (_40384_, _40231_, _33950_);
  and (_40385_, _40384_, _38756_);
  nor (_40386_, _40385_, _40383_);
  and (_41430_, _40386_, _40337_);
  and (_40387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_40388_, _40387_, _40356_);
  nor (_40389_, _40388_, _40336_);
  or (_40390_, _40389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_40391_, _40385_);
  and (_40392_, _40349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_40393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40393_);
  nor (_40395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40393_);
  or (_40396_, _40395_, _40394_);
  and (_40397_, _40356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_40398_, _40397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_40399_, _40398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_40400_, _40399_);
  and (_40401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40402_, _40401_, _40400_);
  or (_40403_, _40402_, _40396_);
  nand (_40404_, _40395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_40405_, _40404_, _40357_);
  and (_40406_, _40405_, _40403_);
  or (_40407_, _40406_, _40392_);
  or (_40408_, _40407_, _40336_);
  and (_40409_, _40408_, _40391_);
  and (_40410_, _40409_, _40390_);
  nor (_40411_, _40391_, _38837_);
  or (_40412_, _40411_, _40410_);
  and (_41433_, _40412_, _43223_);
  nand (_40413_, _40336_, _38837_);
  not (_40414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_40415_, _40355_, _40351_);
  and (_40416_, _40346_, _40393_);
  and (_40417_, _40416_, _40415_);
  and (_40418_, _40417_, _40362_);
  and (_40419_, _40418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40420_, _40419_, _40414_);
  and (_40421_, _40419_, _40414_);
  or (_40422_, _40421_, _40420_);
  and (_40423_, _40422_, _40396_);
  and (_40424_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_40425_, _40424_, _40361_);
  and (_40426_, _40425_, _40358_);
  and (_40427_, _40426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40428_, _40427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_40429_, _40424_, _40364_);
  and (_40430_, _40429_, _40428_);
  and (_40431_, _40430_, _40401_);
  and (_40432_, _40372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40433_, _40432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_40434_, _40433_, _40381_);
  or (_40435_, _40434_, _40431_);
  or (_40436_, _40435_, _40423_);
  or (_40437_, _40436_, _40336_);
  and (_40438_, _40437_, _40391_);
  and (_40439_, _40438_, _40413_);
  and (_40440_, _40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_40441_, _40440_, _40439_);
  and (_41436_, _40441_, _43223_);
  or (_40442_, _40424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_40443_, _40401_, _43223_);
  and (_40444_, _40443_, _40442_);
  not (_40445_, _40424_);
  or (_40446_, _40445_, _40364_);
  nand (_40447_, _40446_, _40444_);
  nor (_40448_, _40447_, _40336_);
  and (_41439_, _40448_, _40391_);
  nor (_40453_, _31860_, _28282_);
  and (_40454_, _40453_, _38757_);
  and (_40455_, _40454_, _31261_);
  or (_40456_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_40457_, _40456_, _43223_);
  nand (_40458_, _40455_, _38837_);
  and (_41441_, _40458_, _40457_);
  not (_40459_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_40460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_40461_, _40460_, _40237_);
  and (_40462_, _40461_, _40256_);
  nor (_40463_, _40462_, _40459_);
  and (_40464_, _40462_, _40459_);
  or (_40465_, _40464_, _40463_);
  nand (_40466_, _40293_, _40239_);
  nor (_40467_, _40466_, _40237_);
  or (_40468_, _40467_, _40233_);
  or (_40477_, _40468_, _40465_);
  nand (_40479_, _40233_, _38816_);
  and (_40480_, _40479_, _43223_);
  and (_41928_, _40480_, _40477_);
  and (_40481_, _40256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_40482_, _40481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_40483_, _40481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_40484_, _40483_, _40482_);
  nand (_40485_, _40484_, _40461_);
  or (_40486_, _40461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_40487_, _40486_, _40485_);
  nand (_40488_, _40274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_40489_, _40488_, _40237_);
  or (_40490_, _40489_, _40282_);
  or (_40491_, _40490_, _40487_);
  nand (_40492_, _40282_, _38808_);
  and (_40493_, _40492_, _43223_);
  and (_41930_, _40493_, _40491_);
  nor (_40494_, _40482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_40495_, _40482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_40496_, _40495_, _40494_);
  and (_40497_, _40496_, _40461_);
  not (_40498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_40499_, _40461_, _40498_);
  nand (_40500_, _40274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_40501_, _40500_, _40237_);
  or (_40502_, _40501_, _40499_);
  or (_40503_, _40502_, _40497_);
  and (_40504_, _40503_, _40284_);
  nor (_40505_, _40284_, _38801_);
  or (_40506_, _40505_, _40504_);
  and (_41932_, _40506_, _43223_);
  nand (_40507_, _40233_, _38793_);
  not (_40508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_40509_, _40461_, _40508_);
  or (_40510_, _40495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_40511_, _40460_, _40261_);
  and (_40512_, _40511_, _40510_);
  and (_40513_, _40274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_40514_, _40513_, _40512_);
  nor (_40515_, _40514_, _40237_);
  or (_40516_, _40515_, _40509_);
  or (_40517_, _40516_, _40233_);
  and (_40518_, _40517_, _43223_);
  and (_41934_, _40518_, _40507_);
  nor (_40519_, _40461_, _40266_);
  nand (_40520_, _40274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_40521_, _40520_, _40237_);
  or (_40522_, _40521_, _40519_);
  nor (_40523_, _40261_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_40524_, _40523_, _40268_);
  and (_40525_, _40524_, _40461_);
  or (_40526_, _40525_, _40522_);
  and (_40527_, _40526_, _40284_);
  nor (_40528_, _40284_, _38786_);
  or (_40529_, _40528_, _40527_);
  and (_41936_, _40529_, _43223_);
  nand (_40530_, _40233_, _38778_);
  and (_40531_, _40243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_40532_, _40268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_40533_, _40268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_40534_, _40533_, _40242_);
  and (_40535_, _40534_, _40532_);
  and (_40536_, _40274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_40537_, _40536_, _40535_);
  nor (_40538_, _40537_, _40237_);
  or (_40539_, _40538_, _40531_);
  or (_40540_, _40539_, _40233_);
  and (_40541_, _40540_, _43223_);
  and (_41938_, _40541_, _40530_);
  nand (_40542_, _40233_, _38770_);
  and (_40543_, _40243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_40544_, _40239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40545_, _40544_, _40256_);
  and (_40546_, _40545_, _40292_);
  nor (_40547_, _40533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_40548_, _40547_, _40242_);
  and (_40549_, _40548_, _40264_);
  nor (_40550_, _40549_, _40546_);
  nor (_40551_, _40550_, _40237_);
  or (_40552_, _40551_, _40543_);
  or (_40553_, _40552_, _40233_);
  and (_40554_, _40553_, _43223_);
  and (_41940_, _40554_, _40542_);
  nand (_40555_, _40237_, _38816_);
  not (_40556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_40557_, _40268_, _40240_);
  nor (_40558_, _40270_, _40238_);
  not (_40559_, _40558_);
  and (_40560_, _40559_, _40557_);
  nor (_40561_, _40560_, _40556_);
  and (_40562_, _40560_, _40556_);
  or (_40563_, _40562_, _40561_);
  or (_40564_, _40563_, _40237_);
  and (_40565_, _40564_, _40555_);
  or (_40566_, _40565_, _40282_);
  nand (_40567_, _40282_, _40556_);
  and (_40568_, _40567_, _43223_);
  and (_41942_, _40568_, _40566_);
  nand (_40569_, _40237_, _38808_);
  not (_40570_, _40241_);
  nor (_40571_, _40271_, _40570_);
  not (_40572_, _40571_);
  nor (_40573_, _40557_, _40241_);
  nor (_40574_, _40573_, _40556_);
  and (_40575_, _40574_, _40572_);
  or (_40576_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_40577_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_40578_, _40577_, _40576_);
  or (_40579_, _40578_, _40237_);
  and (_40580_, _40579_, _40569_);
  or (_40581_, _40580_, _40282_);
  or (_40582_, _40284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_40583_, _40582_, _43223_);
  and (_41944_, _40583_, _40581_);
  nand (_40584_, _40237_, _38801_);
  and (_40585_, _40304_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40586_, _40585_, _40268_);
  and (_40587_, _40586_, _40240_);
  nand (_40588_, _40587_, _40559_);
  and (_40589_, _40588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_40590_, _40558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_40591_, _40590_);
  not (_40592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_40593_, _40304_, _40592_);
  and (_40594_, _40593_, _40268_);
  and (_40595_, _40594_, _40591_);
  or (_40596_, _40595_, _40589_);
  or (_40597_, _40596_, _40237_);
  and (_40598_, _40597_, _40584_);
  or (_40599_, _40598_, _40282_);
  nand (_40600_, _40282_, _40592_);
  and (_40601_, _40600_, _43223_);
  and (_41946_, _40601_, _40599_);
  nand (_40602_, _40237_, _38793_);
  nor (_40603_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_40604_, _40586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_40605_, _40604_, _40270_);
  nor (_40606_, _40605_, _40603_);
  or (_40607_, _40606_, _40570_);
  not (_40608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_40609_, _40587_, _40608_);
  nor (_40610_, _40587_, _40608_);
  or (_40611_, _40610_, _40241_);
  or (_40612_, _40611_, _40609_);
  and (_40613_, _40612_, _40607_);
  or (_40614_, _40613_, _40237_);
  and (_40615_, _40614_, _40602_);
  or (_40616_, _40615_, _40282_);
  nand (_40617_, _40282_, _40608_);
  and (_40618_, _40617_, _43223_);
  and (_41948_, _40618_, _40616_);
  nand (_40619_, _40237_, _38786_);
  or (_40620_, _40605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40621_, _40605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_40622_, _40621_, _40570_);
  and (_40623_, _40622_, _40620_);
  and (_40624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40625_, _40307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_40626_, _40625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_40627_, _40625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40628_, _40627_, _40626_);
  and (_40629_, _40628_, _40311_);
  or (_40630_, _40629_, _40624_);
  or (_40631_, _40630_, _40623_);
  or (_40632_, _40631_, _40237_);
  and (_40633_, _40632_, _40619_);
  or (_40634_, _40633_, _40282_);
  or (_40635_, _40284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40636_, _40635_, _43223_);
  and (_41949_, _40636_, _40634_);
  nand (_40637_, _40237_, _38778_);
  and (_40638_, _40604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40639_, _40638_, _40311_);
  and (_40640_, _40621_, _40241_);
  nor (_40641_, _40640_, _40639_);
  and (_40642_, _40641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_40643_, _40641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_40644_, _40643_, _40642_);
  nor (_40645_, _40644_, _40237_);
  nor (_40646_, _40645_, _40233_);
  and (_40647_, _40646_, _40637_);
  and (_40648_, _40282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_40649_, _40648_, _40647_);
  and (_41951_, _40649_, _43223_);
  nand (_40650_, _40237_, _38770_);
  and (_40651_, _40638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40652_, _40591_, _40651_);
  or (_40653_, _40652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_40654_, _40652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40655_, _40654_, _40653_);
  nor (_40656_, _40655_, _40237_);
  nor (_40657_, _40656_, _40233_);
  and (_40658_, _40657_, _40650_);
  and (_40659_, _40282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_40660_, _40659_, _40658_);
  and (_41953_, _40660_, _43223_);
  nor (_40661_, _40347_, _40336_);
  or (_40662_, _40661_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40663_, _40346_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40664_, _40395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40665_, _40664_, _40415_);
  nand (_40666_, _40665_, _40663_);
  or (_40667_, _40666_, _40336_);
  and (_40668_, _40667_, _40662_);
  or (_40669_, _40668_, _40385_);
  nand (_40670_, _40385_, _38816_);
  and (_40671_, _40670_, _43223_);
  and (_41955_, _40671_, _40669_);
  nand (_40672_, _40385_, _38808_);
  and (_40673_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_40674_, _40663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_40675_, _40663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_40676_, _40675_, _40674_);
  and (_40677_, _40395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40678_, _40677_, _40357_);
  nor (_40679_, _40678_, _40676_);
  nor (_40680_, _40679_, _40336_);
  or (_40681_, _40680_, _40673_);
  or (_40682_, _40681_, _40385_);
  and (_40683_, _40682_, _43223_);
  and (_41957_, _40683_, _40672_);
  nand (_40684_, _40385_, _38801_);
  and (_40685_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_40686_, _40675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_40687_, _40663_, _40352_);
  nor (_40688_, _40687_, _40686_);
  and (_40689_, _40395_, _40357_);
  and (_40690_, _40689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_40691_, _40690_, _40688_);
  nor (_40692_, _40691_, _40336_);
  or (_40693_, _40692_, _40685_);
  or (_40694_, _40693_, _40385_);
  and (_40695_, _40694_, _43223_);
  and (_41959_, _40695_, _40684_);
  and (_40696_, _40354_, _40346_);
  nor (_40697_, _40687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_40698_, _40697_, _40696_);
  and (_40699_, _40689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_40700_, _40699_, _40698_);
  nor (_40701_, _40700_, _40336_);
  and (_40702_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_40703_, _40702_, _40701_);
  and (_40704_, _40703_, _40391_);
  nor (_40705_, _40391_, _38793_);
  or (_40706_, _40705_, _40704_);
  and (_41961_, _40706_, _43223_);
  nand (_40707_, _40385_, _38786_);
  and (_40708_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40709_, _40696_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40710_, _40709_, _40356_);
  and (_40711_, _40689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40712_, _40711_, _40710_);
  nor (_40713_, _40712_, _40336_);
  or (_40714_, _40713_, _40708_);
  or (_40715_, _40714_, _40385_);
  and (_40716_, _40715_, _43223_);
  and (_41963_, _40716_, _40707_);
  nand (_40717_, _40385_, _38778_);
  not (_40718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_40719_, _40356_, _40368_);
  and (_40720_, _40719_, _40718_);
  and (_40721_, _40689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_40722_, _40721_, _40720_);
  nor (_40723_, _40722_, _40336_);
  and (_40724_, _40719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_40725_, _40724_);
  or (_40726_, _40725_, _40336_);
  and (_40727_, _40726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_40728_, _40727_, _40723_);
  or (_40729_, _40728_, _40385_);
  and (_40730_, _40729_, _43223_);
  and (_41965_, _40730_, _40717_);
  and (_40731_, _40726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_40732_, _40395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_40733_, _40732_, _40346_);
  and (_40734_, _40733_, _40415_);
  nor (_40735_, _40725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_40736_, _40735_, _40734_);
  nor (_40737_, _40736_, _40336_);
  or (_40738_, _40737_, _40731_);
  and (_40739_, _40738_, _40391_);
  nor (_40740_, _40391_, _38770_);
  or (_40741_, _40740_, _40739_);
  and (_41967_, _40741_, _43223_);
  nor (_40742_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40743_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_40744_, _40743_, _40742_);
  and (_40745_, _40744_, _40396_);
  and (_40746_, _40424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40747_, _40424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40748_, _40747_, _40401_);
  nor (_40749_, _40748_, _40746_);
  or (_40750_, _40356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40751_, _40356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_40752_, _40751_, _40368_);
  and (_40753_, _40752_, _40750_);
  or (_40754_, _40753_, _40749_);
  or (_40755_, _40754_, _40745_);
  or (_40756_, _40755_, _40336_);
  nand (_40757_, _40336_, _38816_);
  and (_40758_, _40757_, _40756_);
  or (_40759_, _40758_, _40385_);
  or (_40760_, _40391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40761_, _40760_, _43223_);
  and (_41968_, _40761_, _40759_);
  nand (_40762_, _40336_, _38808_);
  or (_40763_, _40743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40764_, _40415_, _40346_);
  and (_40765_, _40764_, _40359_);
  not (_40766_, _40765_);
  or (_40767_, _40766_, _40395_);
  and (_40768_, _40767_, _40396_);
  and (_40769_, _40768_, _40763_);
  and (_40770_, _40424_, _40359_);
  or (_40771_, _40746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_40772_, _40771_, _40401_);
  nor (_40773_, _40772_, _40770_);
  and (_40774_, _40751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_40775_, _40751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_40776_, _40775_, _40349_);
  nor (_40777_, _40776_, _40774_);
  or (_40778_, _40777_, _40773_);
  or (_40779_, _40778_, _40769_);
  or (_40780_, _40779_, _40336_);
  and (_40781_, _40780_, _40391_);
  and (_40782_, _40781_, _40762_);
  and (_40783_, _40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_40784_, _40783_, _40782_);
  and (_41970_, _40784_, _43223_);
  nand (_40785_, _40336_, _38801_);
  and (_40786_, _40764_, _40360_);
  or (_40787_, _40765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_40788_, _40787_, _40394_);
  nor (_40789_, _40788_, _40786_);
  or (_40790_, _40774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40791_, _40360_, _40356_);
  nor (_40792_, _40791_, _40368_);
  and (_40793_, _40792_, _40790_);
  and (_40794_, _40770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40795_, _40794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40796_, _40424_, _40360_);
  nand (_40797_, _40796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40798_, _40797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40799_, _40798_, _40795_);
  or (_40800_, _40799_, _40793_);
  or (_40801_, _40800_, _40789_);
  or (_40802_, _40801_, _40336_);
  and (_40803_, _40802_, _40391_);
  and (_40804_, _40803_, _40785_);
  and (_40805_, _40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_40806_, _40805_, _40804_);
  and (_41972_, _40806_, _43223_);
  nand (_40807_, _40336_, _38793_);
  and (_40808_, _40786_, _40393_);
  not (_40809_, _40808_);
  nor (_40810_, _40809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40811_, _40809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_40812_, _40811_, _40810_);
  and (_40813_, _40812_, _40396_);
  or (_40814_, _40796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_40815_, _40425_);
  and (_40816_, _40815_, _40401_);
  and (_40817_, _40816_, _40814_);
  or (_40818_, _40791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40819_, _40361_, _40356_);
  nor (_40820_, _40819_, _40368_);
  and (_40821_, _40820_, _40818_);
  or (_40822_, _40821_, _40817_);
  or (_40823_, _40822_, _40813_);
  or (_40824_, _40823_, _40336_);
  and (_40825_, _40824_, _40391_);
  and (_40826_, _40825_, _40807_);
  and (_40827_, _40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_40828_, _40827_, _40826_);
  and (_41974_, _40828_, _43223_);
  nand (_40829_, _40336_, _38786_);
  and (_40830_, _40764_, _40361_);
  or (_40831_, _40830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40832_, _40830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40833_, _40832_, _40394_);
  and (_40834_, _40833_, _40831_);
  or (_40835_, _40819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40836_, _40819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40837_, _40836_, _40368_);
  and (_40838_, _40837_, _40835_);
  and (_40839_, _40425_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40840_, _40839_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40841_, _40840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40842_, _40425_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40843_, _40842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40844_, _40843_, _40841_);
  or (_40845_, _40844_, _40838_);
  or (_40846_, _40845_, _40834_);
  or (_40847_, _40846_, _40336_);
  and (_40848_, _40847_, _40391_);
  and (_40849_, _40848_, _40829_);
  and (_40850_, _40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_40851_, _40850_, _40849_);
  and (_41976_, _40851_, _43223_);
  nand (_40852_, _40336_, _38778_);
  nor (_40853_, _40832_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_40854_, _40853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_40855_, _40853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40856_, _40855_, _40396_);
  and (_40857_, _40856_, _40854_);
  not (_40858_, _40426_);
  and (_40859_, _40858_, _40401_);
  or (_40860_, _40842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40861_, _40860_, _40859_);
  nand (_40862_, _40836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40863_, _40836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40864_, _40863_, _40349_);
  and (_40865_, _40864_, _40862_);
  or (_40866_, _40865_, _40861_);
  or (_40867_, _40866_, _40857_);
  or (_40868_, _40867_, _40336_);
  and (_40869_, _40868_, _40391_);
  and (_40870_, _40869_, _40852_);
  and (_40871_, _40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40872_, _40871_, _40870_);
  and (_41978_, _40872_, _43223_);
  nand (_40873_, _40336_, _38770_);
  or (_40874_, _40418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_40875_, _40874_, _40396_);
  nor (_40876_, _40875_, _40419_);
  or (_40877_, _40426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_40878_, _40427_);
  and (_40879_, _40878_, _40401_);
  and (_40880_, _40879_, _40877_);
  or (_40881_, _40372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40882_, _40432_, _40368_);
  and (_40883_, _40882_, _40881_);
  or (_40884_, _40883_, _40880_);
  or (_40885_, _40884_, _40876_);
  or (_40886_, _40885_, _40336_);
  and (_40887_, _40886_, _40391_);
  and (_40888_, _40887_, _40873_);
  and (_40889_, _40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40890_, _40889_, _40888_);
  and (_41980_, _40890_, _43223_);
  nand (_40891_, _40455_, _38816_);
  or (_40892_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40893_, _40892_, _43223_);
  and (_41982_, _40893_, _40891_);
  or (_40894_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40895_, _40894_, _43223_);
  nand (_40896_, _40455_, _38808_);
  and (_41984_, _40896_, _40895_);
  or (_40897_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_40898_, _40897_, _43223_);
  nand (_40899_, _40455_, _38801_);
  and (_41985_, _40899_, _40898_);
  or (_40900_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_40901_, _40900_, _43223_);
  nand (_40902_, _40455_, _38793_);
  and (_41987_, _40902_, _40901_);
  or (_40903_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40904_, _40903_, _43223_);
  nand (_40905_, _40455_, _38786_);
  and (_41989_, _40905_, _40904_);
  or (_40906_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40907_, _40906_, _43223_);
  nand (_40908_, _40455_, _38778_);
  and (_41991_, _40908_, _40907_);
  or (_40909_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_40910_, _40909_, _43223_);
  nand (_40911_, _40455_, _38770_);
  and (_41993_, _40911_, _40910_);
  nor (_40912_, _28424_, _28282_);
  and (_40914_, _40912_, _39418_);
  and (_40916_, _40914_, _39590_);
  and (_40918_, _40916_, _31882_);
  nand (_40920_, _40918_, _31849_);
  and (_40922_, _38751_, _31882_);
  and (_40924_, _40922_, _39616_);
  not (_40926_, _40924_);
  or (_40928_, _40918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_40930_, _40928_, _40926_);
  and (_40932_, _40930_, _40920_);
  nor (_40934_, _40926_, _38837_);
  or (_40936_, _40934_, _40932_);
  and (_43160_, _40936_, _43223_);
  and (_40939_, _40231_, _27624_);
  and (_40941_, _40939_, _39597_);
  and (_40943_, _28424_, _28293_);
  and (_40945_, _40943_, _39418_);
  and (_40947_, _40945_, _39590_);
  and (_40949_, _40947_, _31882_);
  nand (_40951_, _40949_, _31849_);
  or (_40953_, _40949_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40955_, _40953_, _40951_);
  or (_40957_, _40955_, _40941_);
  nand (_40959_, _40941_, _38837_);
  and (_40961_, _40959_, _43223_);
  and (_43163_, _40961_, _40957_);
  and (_40964_, _40939_, _38756_);
  nor (_40966_, _39417_, _28282_);
  nand (_40967_, _40966_, _28424_);
  nor (_40968_, _40967_, _28128_);
  and (_40969_, _40968_, _39558_);
  nand (_40970_, _40969_, _27602_);
  and (_40971_, _40970_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40972_, _40971_, _40964_);
  or (_40973_, _27613_, _33939_);
  and (_40974_, _40973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40975_, _40974_, _39388_);
  and (_40976_, _40975_, _40969_);
  or (_40977_, _40976_, _40972_);
  nand (_40978_, _40964_, _38770_);
  and (_40979_, _40978_, _43223_);
  and (_43165_, _40979_, _40977_);
  not (_40980_, _40964_);
  nor (_40981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_40982_, _40981_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_40983_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_40984_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_40985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40985_);
  and (_40987_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40988_, _40987_, _40986_);
  nor (_40989_, _40988_, _40984_);
  or (_40990_, _40989_, _40983_);
  and (_40991_, _40985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40992_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40993_, _40992_, _40991_);
  nor (_40994_, _40993_, _40984_);
  and (_40995_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40985_);
  and (_40996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40997_, _40996_, _40995_);
  nand (_40998_, _40997_, _40994_);
  or (_40999_, _40998_, _40990_);
  and (_41000_, _40999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_41001_, _41000_, _40982_);
  and (_41002_, _38756_, _31882_);
  and (_41003_, _41002_, _40966_);
  or (_41004_, _41003_, _41001_);
  and (_41005_, _41004_, _40980_);
  nand (_41006_, _41003_, _31849_);
  and (_41007_, _41006_, _41005_);
  nor (_41008_, _40980_, _38837_);
  or (_41009_, _41008_, _41007_);
  and (_43168_, _41009_, _43223_);
  and (_41010_, _40236_, _31926_);
  nand (_41011_, _41010_, _31849_);
  not (_41012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_41013_, _41012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_41014_, _40997_, _40984_);
  not (_41015_, _41014_);
  or (_41016_, _41015_, _40994_);
  or (_41017_, _41016_, _40990_);
  and (_41018_, _41017_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_41019_, _41018_, _41013_);
  or (_41020_, _41019_, _41010_);
  and (_41021_, _41020_, _40980_);
  and (_41022_, _41021_, _41011_);
  nor (_41023_, _40980_, _38778_);
  or (_41024_, _41023_, _41022_);
  and (_43170_, _41024_, _43223_);
  not (_41025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_41026_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _41025_);
  nand (_41027_, _40989_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_41028_, _41014_, _40994_);
  or (_41029_, _41028_, _41027_);
  and (_41030_, _41029_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_41031_, _41030_, _41026_);
  and (_41032_, _40454_, _31926_);
  or (_41033_, _41032_, _41031_);
  and (_41034_, _41033_, _40980_);
  nand (_41035_, _41032_, _31849_);
  and (_41036_, _41035_, _41034_);
  nor (_41037_, _40980_, _38808_);
  or (_41038_, _41037_, _41036_);
  and (_43172_, _41038_, _43223_);
  and (_41039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_41040_, _41027_, _41016_);
  and (_41041_, _41040_, _41039_);
  and (_41042_, _40966_, _38975_);
  or (_41043_, _41042_, _41041_);
  and (_41044_, _41043_, _40980_);
  nand (_41045_, _41042_, _31849_);
  and (_41046_, _41045_, _41044_);
  nor (_41047_, _40980_, _38793_);
  or (_41048_, _41047_, _41046_);
  and (_43174_, _41048_, _43223_);
  nand (_41049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_41050_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40985_);
  and (_41051_, _41050_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_41052_, _41051_, _41049_);
  or (_41053_, _41052_, _40984_);
  and (_41054_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_41055_, _41054_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_41056_, _41055_);
  and (_41057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_41058_, _41057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_41059_, _41058_);
  and (_41060_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_41061_, _41060_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_41062_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_41063_, _41062_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_41064_, _41063_, _41061_);
  and (_41065_, _41064_, _41059_);
  and (_41066_, _41065_, _41056_);
  not (_41067_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_41068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_41069_, _41068_, _41067_);
  nand (_41070_, _41069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_41071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_41072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_41073_, _41072_, _41071_);
  and (_41074_, _41073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_41075_, _41074_);
  and (_41076_, _41075_, _41070_);
  nand (_41077_, _41076_, _41066_);
  and (_41078_, _41077_, _41053_);
  and (_41079_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_41080_, _41079_, _40985_);
  and (_41081_, _41080_, _41078_);
  not (_41082_, _41081_);
  not (_41083_, _41080_);
  and (_41084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40984_);
  not (_41085_, _41084_);
  not (_41086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_41087_, _41057_, _41086_);
  not (_41088_, _41087_);
  not (_41089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_41090_, _41060_, _41089_);
  not (_41091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_41092_, _41062_, _41091_);
  nor (_41093_, _41092_, _41090_);
  and (_41094_, _41093_, _41088_);
  or (_41095_, _41094_, _41085_);
  not (_41096_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_41097_, _41069_, _41096_);
  not (_41098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_41099_, _41073_, _41098_);
  nor (_41100_, _41099_, _41097_);
  not (_41101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_41102_, _41054_, _41101_);
  not (_41103_, _41102_);
  and (_41104_, _41103_, _41100_);
  nor (_41105_, _41104_, _41085_);
  not (_41106_, _41105_);
  and (_41107_, _41106_, _41095_);
  or (_41108_, _41107_, _41083_);
  and (_41109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43223_);
  and (_41110_, _41109_, _41108_);
  and (_43210_, _41110_, _41082_);
  nor (_41111_, _41079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_41112_, _41111_);
  not (_41113_, _41078_);
  and (_41114_, _41107_, _41113_);
  nor (_41115_, _41114_, _41112_);
  nand (_41116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43223_);
  nor (_43212_, _41116_, _41115_);
  and (_41117_, _41076_, _41056_);
  nand (_41118_, _41117_, _41078_);
  or (_41119_, _41105_, _41078_);
  and (_41120_, _41119_, _41080_);
  and (_41121_, _41120_, _41118_);
  or (_41122_, _41121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_41123_, _41082_, _41065_);
  nor (_41124_, _41083_, _41078_);
  not (_41125_, _41124_);
  or (_41126_, _41125_, _41095_);
  and (_41127_, _41126_, _43223_);
  and (_41128_, _41127_, _41123_);
  and (_43214_, _41128_, _41122_);
  and (_41129_, _41118_, _41111_);
  or (_41130_, _41129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_41131_, _41111_, _41078_);
  not (_41132_, _41131_);
  or (_41133_, _41132_, _41065_);
  or (_41134_, _41105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_41135_, _41112_, _41095_);
  and (_41136_, _41135_, _41134_);
  or (_41137_, _41136_, _41078_);
  and (_41138_, _41137_, _43223_);
  and (_41139_, _41138_, _41133_);
  and (_43216_, _41139_, _41130_);
  nand (_41140_, _41114_, _40984_);
  nor (_41141_, _40985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_41142_, _41141_, _41079_);
  and (_41143_, _41142_, _43223_);
  and (_43218_, _41143_, _41140_);
  and (_41144_, _41114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_41145_, _40985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_41146_, _41145_, _41141_);
  nor (_41147_, _41146_, _41113_);
  or (_41148_, _41147_, _41079_);
  or (_41149_, _41148_, _41144_);
  not (_41150_, _41079_);
  or (_41151_, _41146_, _41150_);
  and (_41152_, _41151_, _43223_);
  and (_43220_, _41152_, _41149_);
  and (_41153_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43223_);
  and (_43221_, _41153_, _41079_);
  nor (_43226_, _40981_, rst);
  and (_43228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _43223_);
  nor (_41154_, _41114_, _41079_);
  and (_41155_, _41079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_41156_, _41155_, _41154_);
  and (_00137_, _41156_, _43223_);
  and (_41157_, _41079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_41158_, _41157_, _41154_);
  and (_00139_, _41158_, _43223_);
  and (_41159_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _43223_);
  and (_00141_, _41159_, _41079_);
  not (_41160_, _41092_);
  nor (_41161_, _41099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_41162_, _41161_, _41097_);
  or (_41163_, _41162_, _41102_);
  and (_41164_, _41163_, _41160_);
  or (_41165_, _41164_, _41090_);
  nor (_41166_, _41107_, _41078_);
  and (_41167_, _41166_, _41088_);
  and (_41168_, _41167_, _41165_);
  not (_41169_, _41063_);
  or (_41170_, _41074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_41171_, _41170_, _41070_);
  or (_41172_, _41171_, _41055_);
  and (_41173_, _41172_, _41169_);
  or (_41174_, _41173_, _41061_);
  and (_41175_, _41078_, _41059_);
  and (_41176_, _41175_, _41174_);
  or (_41183_, _41176_, _41079_);
  or (_41184_, _41183_, _41168_);
  or (_41190_, _41150_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_41196_, _41190_, _43223_);
  and (_00143_, _41196_, _41184_);
  nor (_41204_, _41090_, _41087_);
  or (_41205_, _41102_, _41092_);
  and (_41206_, _41100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_41207_, _41206_, _41205_);
  and (_41208_, _41207_, _41204_);
  and (_41209_, _41208_, _41166_);
  not (_41210_, _41061_);
  or (_41211_, _41063_, _41055_);
  and (_41212_, _41076_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_41213_, _41212_, _41211_);
  and (_41214_, _41213_, _41210_);
  and (_41215_, _41214_, _41175_);
  or (_41216_, _41215_, _41079_);
  or (_41217_, _41216_, _41209_);
  or (_41218_, _41150_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_41224_, _41218_, _43223_);
  and (_00144_, _41224_, _41217_);
  and (_41228_, _41103_, _41084_);
  nand (_41229_, _41228_, _41094_);
  or (_41231_, _41229_, _41100_);
  nor (_41232_, _41231_, _41078_);
  nand (_41238_, _41066_, _41053_);
  nor (_41241_, _41238_, _41076_);
  or (_41242_, _41241_, _41079_);
  or (_41243_, _41242_, _41232_);
  or (_41246_, _41150_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_41252_, _41246_, _43223_);
  and (_00146_, _41252_, _41243_);
  and (_41254_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _43223_);
  and (_00148_, _41254_, _41079_);
  and (_41261_, _41079_, _40985_);
  or (_41264_, _41261_, _41115_);
  or (_41265_, _41264_, _41124_);
  and (_00150_, _41265_, _43223_);
  not (_41268_, _41154_);
  and (_41274_, _41268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_41276_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_41279_, _41074_, _40985_);
  or (_41280_, _41279_, _41276_);
  nor (_41286_, _41070_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_41288_, _41286_, _41055_);
  nand (_41290_, _41288_, _41280_);
  or (_41291_, _41056_, _40987_);
  and (_41297_, _41291_, _41290_);
  or (_41300_, _41297_, _41063_);
  or (_41301_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40985_);
  or (_41303_, _41301_, _41169_);
  and (_41309_, _41303_, _41210_);
  and (_41312_, _41309_, _41300_);
  and (_41313_, _41061_, _40987_);
  or (_41314_, _41313_, _41058_);
  or (_41317_, _41314_, _41312_);
  or (_41323_, _41301_, _41059_);
  and (_41325_, _41323_, _41078_);
  and (_41326_, _41325_, _41317_);
  and (_41329_, _41099_, _40985_);
  or (_41335_, _41329_, _41276_);
  and (_41337_, _41097_, _40985_);
  nor (_41338_, _41337_, _41102_);
  nand (_41340_, _41338_, _41335_);
  or (_41346_, _41103_, _40987_);
  and (_41349_, _41346_, _41340_);
  or (_41350_, _41349_, _41092_);
  not (_41352_, _41090_);
  or (_41358_, _41301_, _41160_);
  and (_41361_, _41358_, _41352_);
  and (_41362_, _41361_, _41350_);
  and (_41363_, _41090_, _40987_);
  or (_41368_, _41363_, _41087_);
  or (_41373_, _41368_, _41362_);
  and (_41374_, _41301_, _41166_);
  or (_41375_, _41374_, _41167_);
  and (_41380_, _41375_, _41373_);
  or (_41385_, _41380_, _41326_);
  and (_41386_, _41385_, _41150_);
  or (_41387_, _41386_, _41274_);
  and (_00152_, _41387_, _43223_);
  and (_41396_, _41268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_41397_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40985_);
  and (_41398_, _41397_, _41059_);
  or (_41402_, _41398_, _41065_);
  or (_41407_, _41279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_41408_, _41407_, _41288_);
  nand (_41409_, _41055_, _40996_);
  nand (_41410_, _41409_, _41064_);
  or (_41411_, _41410_, _41408_);
  and (_41412_, _41411_, _41402_);
  and (_41413_, _41058_, _40996_);
  or (_41414_, _41413_, _41412_);
  and (_41416_, _41414_, _41078_);
  and (_41417_, _41102_, _41093_);
  or (_41419_, _41417_, _41087_);
  and (_41420_, _41419_, _40996_);
  or (_41422_, _41329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_41423_, _41338_, _41093_);
  and (_41425_, _41423_, _41422_);
  not (_41426_, _41093_);
  and (_41428_, _41397_, _41426_);
  or (_41429_, _41428_, _41425_);
  and (_41431_, _41429_, _41088_);
  or (_41432_, _41431_, _41420_);
  and (_41434_, _41432_, _41166_);
  or (_41435_, _41434_, _41416_);
  and (_41437_, _41435_, _41150_);
  or (_41438_, _41437_, _41396_);
  and (_00154_, _41438_, _43223_);
  and (_41440_, _41268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_41442_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41443_, _41442_, _41059_);
  and (_41444_, _41443_, _41078_);
  not (_41445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_41446_, _41074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41447_, _41446_, _41445_);
  nor (_41448_, _41070_, _40985_);
  nor (_41449_, _41448_, _41055_);
  nand (_41450_, _41449_, _41447_);
  or (_41451_, _41056_, _40986_);
  and (_41452_, _41451_, _41450_);
  or (_41453_, _41452_, _41063_);
  or (_41454_, _41442_, _41169_);
  and (_41455_, _41454_, _41210_);
  and (_41456_, _41455_, _41453_);
  and (_41457_, _41061_, _40986_);
  or (_41458_, _41457_, _41058_);
  or (_41459_, _41458_, _41456_);
  and (_41460_, _41459_, _41444_);
  or (_41461_, _41442_, _41088_);
  and (_41462_, _41099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_41463_, _41462_, _41445_);
  and (_41464_, _41097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_41465_, _41464_, _41102_);
  nand (_41466_, _41465_, _41463_);
  or (_41467_, _41103_, _40986_);
  and (_41468_, _41467_, _41466_);
  or (_41469_, _41468_, _41092_);
  or (_41470_, _41442_, _41160_);
  and (_41471_, _41470_, _41352_);
  and (_41472_, _41471_, _41469_);
  and (_41473_, _41090_, _40986_);
  or (_41474_, _41473_, _41087_);
  or (_41475_, _41474_, _41472_);
  and (_41476_, _41475_, _41166_);
  and (_41477_, _41476_, _41461_);
  or (_41478_, _41477_, _41460_);
  and (_41479_, _41478_, _41150_);
  or (_41480_, _41479_, _41440_);
  and (_00155_, _41480_, _43223_);
  or (_41481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_41482_, _41481_, _41059_);
  or (_41483_, _41482_, _41065_);
  or (_41484_, _41446_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_41485_, _41484_, _41449_);
  nand (_41486_, _41055_, _40995_);
  nand (_41487_, _41486_, _41064_);
  or (_41488_, _41487_, _41485_);
  and (_41489_, _41488_, _41483_);
  nand (_41490_, _41058_, _40995_);
  nand (_41491_, _41490_, _41078_);
  or (_41492_, _41491_, _41489_);
  and (_41493_, _41481_, _41426_);
  or (_41494_, _41462_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_41495_, _41465_, _41093_);
  and (_41496_, _41495_, _41494_);
  or (_41497_, _41496_, _41493_);
  and (_41498_, _41497_, _41088_);
  and (_41499_, _41419_, _40995_);
  or (_41500_, _41499_, _41107_);
  or (_41501_, _41500_, _41078_);
  or (_41502_, _41501_, _41498_);
  and (_41503_, _41502_, _41492_);
  or (_41504_, _41503_, _41079_);
  or (_41505_, _41154_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_41506_, _41505_, _43223_);
  and (_00157_, _41506_, _41504_);
  or (_41507_, _41112_, _41107_);
  and (_41508_, _41507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_41509_, _41508_, _41131_);
  and (_00159_, _41509_, _43223_);
  and (_41510_, _41108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_41511_, _41510_, _41081_);
  and (_00161_, _41511_, _43223_);
  and (_41512_, _40969_, _27624_);
  or (_41513_, _41512_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_41514_, _41513_, _40980_);
  nand (_41515_, _41512_, _31849_);
  and (_41516_, _41515_, _41514_);
  and (_41517_, _40964_, _38817_);
  or (_41518_, _41517_, _41516_);
  and (_00163_, _41518_, _43223_);
  and (_41519_, _40969_, _33950_);
  or (_41520_, _41519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_41521_, _41520_, _40980_);
  nand (_41522_, _41519_, _31849_);
  and (_41523_, _41522_, _41521_);
  nor (_41524_, _40980_, _38801_);
  or (_41525_, _41524_, _41523_);
  and (_00165_, _41525_, _43223_);
  nand (_41526_, _40969_, _35375_);
  nor (_41527_, _41526_, _31849_);
  and (_41528_, _41526_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_41529_, _41528_, _40964_);
  or (_41530_, _41529_, _41527_);
  nand (_41531_, _40964_, _38786_);
  and (_41532_, _41531_, _43223_);
  and (_00166_, _41532_, _41530_);
  not (_41533_, _40941_);
  and (_41534_, _40947_, _27624_);
  or (_41535_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_41536_, _41535_, _41533_);
  nand (_41537_, _41534_, _31849_);
  and (_41538_, _41537_, _41536_);
  and (_41539_, _40941_, _38817_);
  or (_41540_, _41539_, _41538_);
  and (_00168_, _41540_, _43223_);
  and (_41541_, _40947_, _33199_);
  or (_41542_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_41543_, _41542_, _41533_);
  nand (_41544_, _41541_, _31849_);
  and (_41545_, _41544_, _41543_);
  nor (_41546_, _41533_, _38808_);
  or (_41547_, _41546_, _41545_);
  and (_00170_, _41547_, _43223_);
  nand (_41548_, _40947_, _39846_);
  and (_41549_, _41548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_41550_, _41549_, _40941_);
  and (_41551_, _33983_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_41552_, _41551_, _33972_);
  and (_41553_, _41552_, _40947_);
  or (_41554_, _41553_, _41550_);
  nand (_41555_, _40941_, _38801_);
  and (_41556_, _41555_, _43223_);
  and (_00172_, _41556_, _41554_);
  and (_41557_, _40947_, _34690_);
  or (_41558_, _41557_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_41559_, _41558_, _41533_);
  nand (_41560_, _41557_, _31849_);
  and (_41561_, _41560_, _41559_);
  nor (_41562_, _41533_, _38793_);
  or (_41563_, _41562_, _41561_);
  and (_00174_, _41563_, _43223_);
  and (_41564_, _40947_, _35375_);
  nand (_41565_, _41564_, _31849_);
  or (_41566_, _41564_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_41567_, _41566_, _41565_);
  or (_41568_, _41567_, _40941_);
  nand (_41569_, _40941_, _38786_);
  and (_41570_, _41569_, _43223_);
  and (_00176_, _41570_, _41568_);
  and (_41571_, _40947_, _36171_);
  or (_41572_, _41571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_41573_, _41572_, _41533_);
  nand (_41574_, _41571_, _31849_);
  and (_41575_, _41574_, _41573_);
  nor (_41576_, _41533_, _38778_);
  or (_41577_, _41576_, _41575_);
  and (_00177_, _41577_, _43223_);
  and (_41578_, _40947_, _36909_);
  or (_41579_, _41578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_41580_, _41579_, _41533_);
  nand (_41581_, _41578_, _31849_);
  and (_41582_, _41581_, _41580_);
  nor (_41583_, _41533_, _38770_);
  or (_41584_, _41583_, _41582_);
  and (_00179_, _41584_, _43223_);
  and (_41585_, _40916_, _27624_);
  nand (_41586_, _41585_, _31849_);
  or (_41587_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_41588_, _41587_, _41586_);
  or (_41589_, _41588_, _40924_);
  nand (_41590_, _40924_, _38816_);
  and (_41591_, _41590_, _43223_);
  and (_00181_, _41591_, _41589_);
  and (_41592_, _40916_, _33199_);
  nand (_41593_, _41592_, _31849_);
  or (_41594_, _41592_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_41595_, _41594_, _40926_);
  and (_41596_, _41595_, _41593_);
  nor (_41597_, _40926_, _38808_);
  or (_41598_, _41597_, _41596_);
  and (_00183_, _41598_, _43223_);
  and (_41599_, _33983_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_41600_, _41599_, _33972_);
  and (_41601_, _41600_, _40916_);
  nand (_41602_, _40916_, _39846_);
  and (_41603_, _41602_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_41604_, _41603_, _40924_);
  or (_41605_, _41604_, _41601_);
  nand (_41606_, _40924_, _38801_);
  and (_41607_, _41606_, _43223_);
  and (_00185_, _41607_, _41605_);
  and (_41608_, _40916_, _34690_);
  nand (_41609_, _41608_, _31849_);
  or (_41610_, _41608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_41611_, _41610_, _41609_);
  or (_41612_, _41611_, _40924_);
  nand (_41613_, _40924_, _38793_);
  and (_41614_, _41613_, _43223_);
  and (_00187_, _41614_, _41612_);
  and (_41615_, _40916_, _35375_);
  nand (_41616_, _41615_, _31849_);
  or (_41617_, _41615_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_41618_, _41617_, _40926_);
  and (_41619_, _41618_, _41616_);
  nor (_41620_, _40926_, _38786_);
  or (_41621_, _41620_, _41619_);
  and (_00188_, _41621_, _43223_);
  and (_41622_, _40916_, _36171_);
  nand (_41623_, _41622_, _31849_);
  or (_41624_, _41622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_41625_, _41624_, _41623_);
  or (_41626_, _41625_, _40924_);
  nand (_41627_, _40924_, _38778_);
  and (_41628_, _41627_, _43223_);
  and (_00190_, _41628_, _41626_);
  and (_41629_, _40916_, _36909_);
  nand (_41630_, _41629_, _31849_);
  or (_41631_, _41629_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_41632_, _41631_, _40926_);
  and (_41633_, _41632_, _41630_);
  nor (_41634_, _40926_, _38770_);
  or (_41635_, _41634_, _41633_);
  and (_00192_, _41635_, _43223_);
  and (_41636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_41638_, _40981_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_41639_, _41638_, _41637_);
  not (_41640_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_41641_, _41640_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_41642_, _41641_, _41639_);
  nor (_41643_, _41642_, _41636_);
  or (_41644_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41645_, _41644_, _43223_);
  nor (_00552_, _41645_, _41643_);
  nor (_41646_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41647_, _41646_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41648_, _41646_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_41649_, _41648_, _43223_);
  and (_00555_, _41649_, _41647_);
  not (_41650_, rxd_i);
  and (_41651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _41650_);
  nor (_41652_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_41653_, _41652_);
  and (_41654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_41655_, _41654_, _41653_);
  and (_41656_, _41655_, _41651_);
  not (_41657_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_41658_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _41657_);
  and (_41659_, _41658_, _41652_);
  or (_41660_, _41659_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_41661_, _41660_, _41656_);
  and (_41662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _43223_);
  and (_00558_, _41662_, _41661_);
  and (_41663_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_41664_, _41663_, _41653_);
  not (_41665_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_41666_, _41652_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41667_, _41666_, _41665_);
  nor (_41668_, _41667_, _41664_);
  not (_41669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_41670_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _41669_);
  not (_41671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_41672_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _41671_);
  and (_41673_, _41672_, _41670_);
  not (_41674_, _41673_);
  or (_41675_, _41674_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_41676_, _41673_, _41664_);
  and (_41677_, _41664_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41678_, _41677_, _41676_);
  and (_41679_, _41678_, _41675_);
  or (_41680_, _41679_, _41668_);
  and (_41681_, _41652_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_41682_, _41681_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not (_41683_, _41682_);
  or (_41684_, _41683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_41685_, _41684_, _41680_);
  nand (_00560_, _41685_, _41662_);
  not (_41686_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_41687_, _41664_);
  nor (_41688_, _41665_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_41689_, _41688_);
  not (_41690_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41691_, _41652_, _41690_);
  and (_41692_, _41691_, _41689_);
  and (_41693_, _41692_, _41687_);
  nor (_41694_, _41693_, _41686_);
  and (_41695_, _41693_, rxd_i);
  or (_41696_, _41695_, rst);
  or (_00563_, _41696_, _41694_);
  nor (_41697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41698_, _41697_, _41670_);
  and (_41699_, _41698_, _41677_);
  nand (_41700_, _41699_, _41650_);
  or (_41701_, _41699_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_41702_, _41701_, _43223_);
  and (_00566_, _41702_, _41700_);
  and (_41703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41704_, _41703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41705_, _41704_, _41669_);
  and (_41706_, _41705_, _41677_);
  and (_41707_, _41655_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41708_, _41707_, _41677_);
  nor (_41709_, _41704_, _41687_);
  or (_41710_, _41709_, _41708_);
  and (_41711_, _41710_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_41712_, _41711_, _41706_);
  and (_00568_, _41712_, _43223_);
  and (_41713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _43223_);
  nand (_41714_, _41713_, _41690_);
  nand (_41715_, _41662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_00571_, _41715_, _41714_);
  and (_41716_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41690_);
  not (_41717_, _41655_);
  not (_41718_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_41719_, _41659_, _41718_);
  and (_41720_, _41719_, _41717_);
  and (_41721_, _41720_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_41722_, _41721_, _41664_);
  or (_41723_, _41673_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_41724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41725_, _41724_, _41676_);
  and (_41726_, _41725_, _41723_);
  and (_41727_, _41726_, _41722_);
  or (_41728_, _41727_, _41682_);
  nand (_41729_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41730_, _41729_, _41664_);
  or (_41731_, _41730_, _41674_);
  and (_41732_, _41731_, _41683_);
  or (_41733_, _41732_, rxd_i);
  and (_41734_, _41733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41735_, _41734_, _41728_);
  or (_41736_, _41735_, _41716_);
  and (_00574_, _41736_, _43223_);
  and (_41737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41738_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41739_, _41638_, _41738_);
  or (_41740_, _41739_, _41641_);
  nor (_41741_, _41740_, _41737_);
  or (_41742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41743_, _41742_, _43223_);
  nor (_00576_, _41743_, _41741_);
  nor (_41744_, _41741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41745_, _41744_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41746_, _41744_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_41747_, _41746_, _43223_);
  and (_00579_, _41747_, _41745_);
  and (_41748_, _41681_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_41749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_41750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_41751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41752_, _41751_, _41750_);
  and (_41753_, _41752_, _41749_);
  not (_41754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_41755_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_41756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41757_, _41756_, _41755_);
  and (_41758_, _41757_, _41754_);
  and (_41759_, _41758_, _41753_);
  or (_41760_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_41761_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41762_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41763_, _41762_, _41761_);
  and (_41764_, _41653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_41765_, _41764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41766_, _41765_, _41763_);
  not (_41767_, _41766_);
  or (_41768_, _41767_, _41760_);
  and (_41769_, _41763_, _41764_);
  not (_41770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or (_41771_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41770_);
  or (_41772_, _41771_, _41769_);
  and (_41773_, _41772_, _41768_);
  or (_41774_, _41773_, _41748_);
  not (_41775_, _41748_);
  not (_41776_, _41759_);
  or (_41777_, _41776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_41778_, _41777_, _41760_);
  or (_41779_, _41778_, _41775_);
  nand (_41780_, _41779_, _41774_);
  and (_41781_, _40453_, _33188_);
  and (_41782_, _41781_, _31261_);
  and (_41783_, _41782_, _39580_);
  nor (_41784_, _41783_, rst);
  nand (_41785_, _41784_, _41780_);
  not (_41786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_41787_, _41783_, _43223_);
  nand (_41788_, _41787_, _41786_);
  and (_00582_, _41788_, _41785_);
  nor (_41789_, _41776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_41790_, _41769_, _41789_);
  and (_41791_, _41759_, _41748_);
  or (_41792_, _41770_, rst);
  nor (_41793_, _41792_, _41791_);
  and (_41794_, _41793_, _41790_);
  or (_00584_, _41794_, _41787_);
  or (_41795_, _41767_, _41789_);
  or (_41796_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_41797_, _41681_, _41770_);
  and (_41798_, _41797_, _41796_);
  and (_41799_, _41798_, _41795_);
  or (_41800_, _41799_, _41791_);
  and (_00587_, _41800_, _41784_);
  and (_41801_, _41765_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_41802_, _41801_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_41803_, _41802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_41804_, _41803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_41805_, _41803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41806_, _41805_, _41804_);
  and (_00590_, _41806_, _41784_);
  and (_41807_, _41787_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_41808_, _41766_, _41748_);
  and (_41809_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41810_, _41809_, _41784_);
  or (_00592_, _41810_, _41807_);
  and (_41811_, _40922_, _38756_);
  or (_41812_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_41813_, _41812_, _43223_);
  nand (_41814_, _41811_, _38837_);
  and (_00595_, _41814_, _41813_);
  and (_41815_, _40939_, _39580_);
  and (_41816_, _40914_, _39558_);
  and (_41817_, _41816_, _31882_);
  nand (_41818_, _41817_, _31849_);
  or (_41819_, _41817_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_41820_, _41819_, _41818_);
  or (_41821_, _41820_, _41815_);
  nand (_41822_, _41815_, _38837_);
  and (_41823_, _41822_, _43223_);
  and (_00598_, _41823_, _41821_);
  nor (_41824_, _41682_, _41676_);
  not (_41825_, _41824_);
  nor (_41826_, _41720_, _41664_);
  nor (_41827_, _41826_, _41825_);
  nor (_41828_, _41827_, _41690_);
  or (_41829_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_41830_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _41690_);
  or (_41831_, _41830_, _41824_);
  and (_41832_, _41831_, _43223_);
  and (_01215_, _41832_, _41829_);
  or (_41833_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_41834_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _41690_);
  or (_41835_, _41834_, _41824_);
  and (_41836_, _41835_, _43223_);
  and (_01217_, _41836_, _41833_);
  or (_41837_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_41838_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41690_);
  or (_41839_, _41838_, _41824_);
  and (_41840_, _41839_, _43223_);
  and (_01219_, _41840_, _41837_);
  or (_41841_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_41842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41690_);
  or (_41843_, _41842_, _41824_);
  and (_41844_, _41843_, _43223_);
  and (_01221_, _41844_, _41841_);
  or (_41845_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_41846_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41690_);
  or (_41847_, _41846_, _41824_);
  and (_41848_, _41847_, _43223_);
  and (_01223_, _41848_, _41845_);
  or (_41849_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_41850_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41690_);
  or (_41851_, _41850_, _41824_);
  and (_41852_, _41851_, _43223_);
  and (_01225_, _41852_, _41849_);
  or (_41853_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_41854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41690_);
  or (_41855_, _41854_, _41824_);
  and (_41856_, _41855_, _43223_);
  and (_01226_, _41856_, _41853_);
  or (_41857_, _41828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_41858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _41690_);
  or (_41859_, _41858_, _41824_);
  and (_41860_, _41859_, _43223_);
  and (_01228_, _41860_, _41857_);
  nor (_41861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_41862_, _41861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_41863_, _41674_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_41864_, _41673_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41865_, _41864_, _41664_);
  and (_41866_, _41865_, _41863_);
  or (_41867_, _41655_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41868_, _41867_, _41719_);
  and (_41869_, _41868_, _41687_);
  or (_41870_, _41869_, _41866_);
  or (_41871_, _41870_, _41682_);
  or (_41872_, _41683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41873_, _41872_, _41662_);
  and (_41874_, _41873_, _41871_);
  or (_01230_, _41874_, _41862_);
  and (_41875_, _41673_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_41876_, _41875_, _41720_);
  or (_41877_, _41876_, _41827_);
  and (_41878_, _41877_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41879_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _41690_);
  nand (_41880_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41881_, _41880_, _41824_);
  or (_41882_, _41881_, _41879_);
  or (_41883_, _41882_, _41878_);
  and (_01232_, _41883_, _43223_);
  not (_41884_, _41828_);
  and (_41885_, _41884_, _41713_);
  or (_41886_, _41876_, _41825_);
  and (_41887_, _41662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_41888_, _41887_, _41886_);
  or (_01234_, _41888_, _41885_);
  or (_41889_, _41706_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_41890_, _41706_, _41650_);
  and (_41891_, _41890_, _43223_);
  and (_01236_, _41891_, _41889_);
  or (_41892_, _41708_, _41671_);
  or (_41893_, _41677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41894_, _41893_, _43223_);
  and (_01238_, _41894_, _41892_);
  and (_41895_, _41708_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_41896_, _41697_, _41703_);
  and (_41897_, _41896_, _41677_);
  or (_41898_, _41897_, _41895_);
  and (_01240_, _41898_, _43223_);
  and (_41899_, _41710_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41900_, _41703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41901_, _41900_, _41709_);
  or (_41902_, _41901_, _41899_);
  and (_01242_, _41902_, _43223_);
  and (_41903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41690_);
  and (_41904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41905_, _41904_, _41903_);
  and (_01244_, _41905_, _43223_);
  and (_41906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41690_);
  and (_41907_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41908_, _41907_, _41906_);
  and (_01246_, _41908_, _43223_);
  and (_41909_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41690_);
  and (_41910_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41911_, _41910_, _41909_);
  and (_01248_, _41911_, _43223_);
  and (_41912_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41690_);
  and (_41913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41914_, _41913_, _41912_);
  and (_01250_, _41914_, _43223_);
  and (_41915_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41690_);
  and (_41916_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41917_, _41916_, _41915_);
  and (_01252_, _41917_, _43223_);
  and (_41918_, _41662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01254_, _41918_, _41862_);
  and (_41919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41920_, _41919_, _41879_);
  and (_01256_, _41920_, _43223_);
  nor (_41921_, _41765_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41922_, _41921_, _41801_);
  and (_01258_, _41922_, _41784_);
  nor (_41923_, _41801_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_41924_, _41923_, _41802_);
  and (_01260_, _41924_, _41784_);
  nor (_41925_, _41802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_41926_, _41925_, _41803_);
  and (_01262_, _41926_, _41784_);
  or (_41927_, _41766_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41929_, _41767_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41931_, _41929_, _41927_);
  and (_41933_, _41931_, _41775_);
  and (_41935_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41937_, _41935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41939_, _41937_, _41748_);
  or (_41941_, _41939_, _41933_);
  and (_41943_, _41941_, _41784_);
  nor (_41945_, _41653_, _38816_);
  and (_41947_, _41945_, _41787_);
  or (_01264_, _41947_, _41943_);
  not (_41950_, _41808_);
  and (_41952_, _41950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_41954_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_41956_, _41954_, _41952_);
  and (_41958_, _41956_, _41784_);
  nand (_41960_, _41652_, _38808_);
  nand (_41962_, _41653_, _38816_);
  and (_41964_, _41962_, _41787_);
  and (_41966_, _41964_, _41960_);
  or (_01266_, _41966_, _41958_);
  nor (_41969_, _41808_, _41754_);
  and (_41971_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_41973_, _41971_, _41969_);
  and (_41975_, _41973_, _41784_);
  nand (_41977_, _41652_, _38801_);
  nand (_41979_, _41653_, _38808_);
  and (_41981_, _41979_, _41787_);
  and (_41983_, _41981_, _41977_);
  or (_01268_, _41983_, _41975_);
  nor (_41986_, _41808_, _41750_);
  and (_41988_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_41990_, _41988_, _41986_);
  and (_41992_, _41990_, _41784_);
  nand (_41994_, _41653_, _38801_);
  nand (_41995_, _41652_, _38793_);
  and (_41996_, _41995_, _41787_);
  and (_41997_, _41996_, _41994_);
  or (_01269_, _41997_, _41992_);
  and (_41998_, _41950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41999_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or (_42000_, _41999_, _41998_);
  and (_42001_, _42000_, _41784_);
  nand (_42002_, _41653_, _38793_);
  nand (_42003_, _41652_, _38786_);
  and (_42004_, _42003_, _41787_);
  and (_42005_, _42004_, _42002_);
  or (_01271_, _42005_, _42001_);
  and (_42006_, _41950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_42007_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_42008_, _42007_, _42006_);
  and (_42009_, _42008_, _41784_);
  nand (_42010_, _41652_, _38778_);
  nand (_42011_, _41653_, _38786_);
  and (_42012_, _42011_, _41787_);
  and (_42013_, _42012_, _42010_);
  or (_01273_, _42013_, _42009_);
  and (_42014_, _41950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_42015_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_42016_, _42015_, _42014_);
  and (_42017_, _42016_, _41784_);
  nand (_42018_, _41652_, _38770_);
  nand (_42019_, _41653_, _38778_);
  and (_42020_, _42019_, _41787_);
  and (_42021_, _42020_, _42018_);
  or (_01275_, _42021_, _42017_);
  and (_42022_, _41950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_42023_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_42024_, _42023_, _42022_);
  and (_42025_, _42024_, _41784_);
  nand (_42026_, _41652_, _38837_);
  nand (_42027_, _41653_, _38770_);
  and (_42028_, _42027_, _41787_);
  and (_42029_, _42028_, _42026_);
  or (_01277_, _42029_, _42025_);
  and (_42030_, _41783_, _41653_);
  nand (_42031_, _42030_, _38837_);
  and (_42032_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_42033_, _41950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_42034_, _42033_, _42032_);
  or (_42035_, _42034_, _41783_);
  and (_42036_, _42035_, _43223_);
  and (_01279_, _42036_, _42031_);
  and (_42037_, _41950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_42038_, _41808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_42039_, _42038_, _42037_);
  and (_42040_, _42039_, _41784_);
  or (_42041_, _41640_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_42042_, _42041_, _41653_);
  and (_42043_, _42042_, _41787_);
  or (_01281_, _42043_, _42040_);
  nand (_42044_, _41811_, _38816_);
  or (_42045_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_42046_, _42045_, _43223_);
  and (_01283_, _42046_, _42044_);
  or (_42047_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_42048_, _42047_, _43223_);
  nand (_42049_, _41811_, _38808_);
  and (_01285_, _42049_, _42048_);
  or (_42050_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_42051_, _42050_, _43223_);
  nand (_42052_, _41811_, _38801_);
  and (_01287_, _42052_, _42051_);
  or (_42053_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_42054_, _42053_, _43223_);
  nand (_42055_, _41811_, _38793_);
  and (_01289_, _42055_, _42054_);
  or (_42056_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_42057_, _42056_, _43223_);
  nand (_42058_, _41811_, _38786_);
  and (_01291_, _42058_, _42057_);
  or (_42059_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_42060_, _42059_, _43223_);
  nand (_42061_, _41811_, _38778_);
  and (_01293_, _42061_, _42060_);
  or (_42062_, _41811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_42063_, _42062_, _43223_);
  nand (_42064_, _41811_, _38770_);
  and (_01295_, _42064_, _42063_);
  not (_42065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_42066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _42065_);
  or (_42067_, _42066_, _41652_);
  nor (_42068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_42069_, _42068_, _42067_);
  or (_42070_, _42069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_42071_, _42070_, _41816_);
  or (_42072_, _27624_, _41657_);
  nand (_42073_, _42072_, _41816_);
  or (_42074_, _42073_, _39473_);
  and (_42075_, _42074_, _42071_);
  or (_42076_, _42075_, _41815_);
  nand (_42077_, _41815_, _38816_);
  and (_42078_, _42077_, _43223_);
  and (_01297_, _42078_, _42076_);
  or (_42079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_42080_, _42079_, _41816_);
  not (_42081_, _33199_);
  nor (_42082_, _42081_, _31849_);
  nand (_42083_, _42081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_42084_, _42083_, _41816_);
  or (_42085_, _42084_, _42082_);
  and (_42086_, _42085_, _42080_);
  or (_42087_, _42086_, _41815_);
  nand (_42088_, _41815_, _38808_);
  and (_42089_, _42088_, _43223_);
  and (_01298_, _42089_, _42087_);
  not (_42090_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not (_42091_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_42092_, _41666_, _42091_);
  nor (_42093_, _42092_, _42090_);
  and (_42094_, _42092_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_42095_, _42094_, _42093_);
  or (_42096_, _42095_, _41816_);
  or (_42097_, _33950_, _42090_);
  nand (_42098_, _42097_, _41816_);
  or (_42099_, _42098_, _33972_);
  and (_42100_, _42099_, _42096_);
  or (_42101_, _42100_, _41815_);
  nand (_42102_, _41815_, _38801_);
  and (_42103_, _42102_, _43223_);
  and (_01300_, _42103_, _42101_);
  and (_42104_, _41816_, _34690_);
  nand (_42105_, _42104_, _31849_);
  not (_42106_, _41815_);
  or (_42107_, _42104_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_42108_, _42107_, _42106_);
  and (_42109_, _42108_, _42105_);
  nor (_42110_, _42106_, _38793_);
  or (_42111_, _42110_, _42109_);
  and (_01302_, _42111_, _43223_);
  and (_42112_, _41816_, _35375_);
  nand (_42113_, _42112_, _31849_);
  or (_42114_, _42112_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_42115_, _42114_, _42106_);
  and (_42116_, _42115_, _42113_);
  nor (_42117_, _42106_, _38786_);
  or (_42118_, _42117_, _42116_);
  and (_01304_, _42118_, _43223_);
  and (_42119_, _41816_, _36171_);
  nand (_42120_, _42119_, _31849_);
  or (_42121_, _42119_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_42122_, _42121_, _42120_);
  or (_42123_, _42122_, _41815_);
  nand (_42124_, _41815_, _38778_);
  and (_42125_, _42124_, _43223_);
  and (_01306_, _42125_, _42123_);
  and (_42126_, _41816_, _36909_);
  nand (_42127_, _42126_, _31849_);
  or (_42128_, _42126_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_42129_, _42128_, _42106_);
  and (_42130_, _42129_, _42127_);
  nor (_42131_, _42106_, _38770_);
  or (_42132_, _42131_, _42130_);
  and (_01308_, _42132_, _43223_);
  and (_01612_, t2_i, _43223_);
  nor (_42133_, t2_i, rst);
  and (_01615_, _42133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_42134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _43223_);
  nor (_01618_, _42134_, t2ex_i);
  and (_01621_, t2ex_i, _43223_);
  and (_42135_, _38753_, _39236_);
  and (_42136_, _42135_, _40384_);
  nand (_42137_, _42136_, _38837_);
  and (_42138_, _42135_, _40232_);
  not (_42139_, _42138_);
  not (_42140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_42141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_42142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_42143_, _42142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_42144_, _42143_, _42141_);
  nor (_42145_, _42144_, _42140_);
  and (_42146_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_42147_, _42146_, _42145_);
  or (_42148_, _42136_, _42147_);
  and (_42149_, _42148_, _42139_);
  and (_42150_, _42149_, _42137_);
  and (_42151_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_42152_, _42151_, _42150_);
  and (_01624_, _42152_, _43223_);
  nand (_42153_, _42138_, _38837_);
  not (_42154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_42155_, _42144_);
  nor (_42156_, _42136_, _42155_);
  nor (_42157_, _42156_, _42154_);
  and (_42158_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_42159_, _42158_, _42157_);
  or (_42160_, _42159_, _42138_);
  and (_42161_, _42160_, _43223_);
  and (_01627_, _42161_, _42153_);
  not (_42162_, _42142_);
  or (_42163_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_42164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_42165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _42164_);
  and (_42166_, _42165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_42167_, _42166_, _42163_);
  and (_42168_, _42167_, _42162_);
  and (_42169_, _42135_, _40335_);
  and (_42170_, _40231_, _36171_);
  and (_42171_, _42170_, _42135_);
  nor (_42172_, _42171_, _42169_);
  and (_42173_, _42172_, _42168_);
  or (_42174_, _42173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_42175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_42176_, _42175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_42177_, _42176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_42178_, _42177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_42179_, _42178_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_42180_, _42179_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_42181_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_42182_, _42181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_42183_, _42182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_42184_, _42183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_42185_, _42184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_42186_, _42185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_42187_, _42186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_42188_, _42187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_42189_, _42188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_42190_, _42189_);
  nand (_42191_, _42190_, _42173_);
  and (_42192_, _42191_, _43223_);
  and (_01630_, _42192_, _42174_);
  nand (_42193_, _42169_, _38837_);
  and (_42194_, _42135_, _36171_);
  and (_42195_, _42194_, _40231_);
  not (_42196_, _42195_);
  not (_42197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_42198_, _42141_, _42197_);
  and (_42199_, _42198_, _42142_);
  and (_42200_, _42199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not (_42201_, _42199_);
  nor (_42202_, _42143_, _42140_);
  and (_42203_, _42189_, _42167_);
  and (_42204_, _42203_, _42202_);
  and (_42205_, _42180_, _42167_);
  or (_42206_, _42205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_42207_, _42205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_42208_, _42207_, _42206_);
  or (_42209_, _42208_, _42204_);
  and (_42210_, _42209_, _42201_);
  or (_42211_, _42210_, _42200_);
  or (_42212_, _42211_, _42169_);
  and (_42213_, _42212_, _42196_);
  and (_42214_, _42213_, _42193_);
  and (_42215_, _42195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_42216_, _42215_, _42214_);
  and (_01633_, _42216_, _43223_);
  and (_42217_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_42218_, _42188_, _42167_);
  or (_42219_, _42218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_42220_, _42143_, _42154_);
  nand (_42221_, _42220_, _42203_);
  and (_42222_, _42221_, _42219_);
  or (_42223_, _42222_, _42199_);
  nand (_42224_, _42199_, _42154_);
  and (_42225_, _42224_, _42172_);
  and (_42226_, _42225_, _42223_);
  nor (_42227_, _42196_, _38837_);
  or (_42228_, _42227_, _42226_);
  or (_42229_, _42228_, _42217_);
  and (_01636_, _42229_, _43223_);
  and (_42230_, _42201_, _42167_);
  and (_42231_, _42230_, _42142_);
  nand (_42232_, _42231_, _42189_);
  nand (_42233_, _42232_, _42172_);
  or (_42234_, _42172_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42235_, _42234_, _43223_);
  and (_01639_, _42235_, _42233_);
  or (_42236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42237_, _40945_, _39240_);
  or (_42238_, _42237_, _42236_);
  not (_42239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_42240_, _31882_, _42239_);
  nand (_42241_, _42240_, _42237_);
  or (_42242_, _42241_, _39253_);
  and (_42243_, _42242_, _42238_);
  and (_42244_, _42135_, _40939_);
  or (_42245_, _42244_, _42243_);
  nand (_42246_, _42244_, _38837_);
  and (_42247_, _42246_, _43223_);
  and (_01642_, _42247_, _42245_);
  nand (_42248_, _42136_, _38816_);
  or (_42249_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not (_42250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_42251_, _42144_, _42250_);
  and (_42252_, _42251_, _42249_);
  or (_42253_, _42252_, _42136_);
  and (_42254_, _42253_, _42248_);
  or (_42255_, _42254_, _42138_);
  not (_42256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_42257_, _42138_, _42256_);
  and (_42258_, _42257_, _43223_);
  and (_02128_, _42258_, _42255_);
  nand (_42259_, _42136_, _38808_);
  and (_42260_, _42155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_42261_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_42262_, _42261_, _42260_);
  or (_42263_, _42262_, _42136_);
  and (_42264_, _42263_, _42139_);
  and (_42265_, _42264_, _42259_);
  and (_42266_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_42267_, _42266_, _42265_);
  and (_02129_, _42267_, _43223_);
  nand (_42268_, _42136_, _38801_);
  and (_42269_, _42155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_42270_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_42271_, _42270_, _42269_);
  or (_42272_, _42271_, _42136_);
  and (_42273_, _42272_, _42139_);
  and (_42274_, _42273_, _42268_);
  and (_42275_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_42276_, _42275_, _42274_);
  and (_02131_, _42276_, _43223_);
  nand (_42277_, _42136_, _38793_);
  and (_42278_, _42155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42279_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_42280_, _42279_, _42278_);
  or (_42281_, _42280_, _42136_);
  and (_42282_, _42281_, _42139_);
  and (_42283_, _42282_, _42277_);
  and (_42284_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_42285_, _42284_, _42283_);
  and (_02133_, _42285_, _43223_);
  nand (_42286_, _42136_, _38786_);
  and (_42287_, _42155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_42288_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_42289_, _42288_, _42287_);
  or (_42290_, _42289_, _42136_);
  and (_42291_, _42290_, _42139_);
  and (_42292_, _42291_, _42286_);
  and (_42293_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_42294_, _42293_, _42292_);
  and (_02135_, _42294_, _43223_);
  nand (_42295_, _42136_, _38778_);
  and (_42296_, _42155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_42297_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_42298_, _42297_, _42296_);
  or (_42299_, _42298_, _42136_);
  and (_42300_, _42299_, _42139_);
  and (_42301_, _42300_, _42295_);
  and (_42302_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_42303_, _42302_, _42301_);
  and (_02136_, _42303_, _43223_);
  nand (_42304_, _42136_, _38770_);
  and (_42305_, _42155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_42306_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_42307_, _42306_, _42305_);
  or (_42308_, _42307_, _42136_);
  and (_42309_, _42308_, _42139_);
  and (_42310_, _42309_, _42304_);
  and (_42311_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_42312_, _42311_, _42310_);
  and (_02138_, _42312_, _43223_);
  or (_42313_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_42314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_42315_, _42156_, _42314_);
  and (_42316_, _42315_, _42313_);
  or (_42317_, _42316_, _42138_);
  nand (_42318_, _42138_, _38816_);
  and (_42319_, _42318_, _43223_);
  and (_02140_, _42319_, _42317_);
  nand (_42320_, _42138_, _38808_);
  or (_42321_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  not (_42322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_42323_, _42156_, _42322_);
  and (_42324_, _42323_, _42321_);
  or (_42325_, _42324_, _42138_);
  and (_42326_, _42325_, _43223_);
  and (_02142_, _42326_, _42320_);
  nand (_42327_, _42138_, _38801_);
  not (_42328_, _42156_);
  and (_42329_, _42328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_42330_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_42331_, _42330_, _42329_);
  or (_42332_, _42331_, _42138_);
  and (_42333_, _42332_, _43223_);
  and (_02143_, _42333_, _42327_);
  nand (_42334_, _42138_, _38793_);
  and (_42335_, _42328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_42336_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42337_, _42336_, _42335_);
  or (_42338_, _42337_, _42138_);
  and (_42339_, _42338_, _43223_);
  and (_02145_, _42339_, _42334_);
  nand (_42340_, _42138_, _38786_);
  and (_42341_, _42328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_42342_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42343_, _42342_, _42341_);
  or (_42344_, _42343_, _42138_);
  and (_42345_, _42344_, _43223_);
  and (_02147_, _42345_, _42340_);
  nand (_42346_, _42138_, _38778_);
  and (_42347_, _42328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_42348_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_42349_, _42348_, _42347_);
  or (_42350_, _42349_, _42138_);
  and (_42351_, _42350_, _43223_);
  and (_02149_, _42351_, _42346_);
  nand (_42352_, _42138_, _38770_);
  and (_42353_, _42328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_42354_, _42156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_42355_, _42354_, _42353_);
  or (_42356_, _42355_, _42138_);
  and (_42357_, _42356_, _43223_);
  and (_02150_, _42357_, _42352_);
  or (_42358_, _42167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_42359_, _42167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_42360_, _42143_, _42256_);
  nand (_42361_, _42360_, _42189_);
  nand (_42362_, _42361_, _42359_);
  and (_42363_, _42362_, _42358_);
  or (_42364_, _42363_, _42199_);
  and (_42365_, _42199_, _42256_);
  nor (_42366_, _42365_, _42169_);
  and (_42367_, _42366_, _42364_);
  and (_42368_, _42169_, _38817_);
  or (_42369_, _42368_, _42195_);
  or (_42370_, _42369_, _42367_);
  nand (_42371_, _42171_, _42250_);
  and (_42372_, _42371_, _43223_);
  and (_02152_, _42372_, _42370_);
  not (_42373_, _42143_);
  and (_42374_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_42375_, _42374_, _42230_);
  and (_42376_, _42375_, _42189_);
  and (_42377_, _42199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  not (_42378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor (_42379_, _42359_, _42378_);
  and (_42380_, _42359_, _42378_);
  or (_42381_, _42380_, _42379_);
  and (_42382_, _42381_, _42201_);
  nor (_42383_, _42382_, _42377_);
  nand (_42384_, _42383_, _42172_);
  or (_42385_, _42384_, _42376_);
  nand (_42386_, _42169_, _38808_);
  nand (_42387_, _42171_, _42378_);
  and (_42388_, _42387_, _43223_);
  and (_42389_, _42388_, _42386_);
  and (_02154_, _42389_, _42385_);
  not (_42390_, _42169_);
  or (_42391_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_42392_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_42393_, _42392_, _42203_);
  nand (_42394_, _42175_, _42167_);
  and (_42395_, _42394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_42396_, _42394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_42397_, _42396_, _42199_);
  or (_42398_, _42397_, _42395_);
  or (_42399_, _42398_, _42393_);
  nand (_42400_, _42399_, _42391_);
  nand (_42401_, _42400_, _42390_);
  nand (_42402_, _42169_, _38801_);
  and (_42403_, _42402_, _42401_);
  or (_42404_, _42403_, _42171_);
  or (_42405_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_42406_, _42405_, _43223_);
  and (_02156_, _42406_, _42404_);
  and (_42407_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_42408_, _42407_, _42203_);
  nand (_42409_, _42176_, _42167_);
  and (_42410_, _42409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_42411_, _42409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_42412_, _42411_, _42199_);
  or (_42413_, _42412_, _42410_);
  or (_42414_, _42413_, _42408_);
  nor (_42415_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor (_42416_, _42415_, _42169_);
  and (_42417_, _42416_, _42414_);
  nor (_42418_, _42390_, _38793_);
  or (_42419_, _42418_, _42417_);
  or (_42420_, _42419_, _42195_);
  or (_42421_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_42422_, _42421_, _43223_);
  and (_02157_, _42422_, _42420_);
  or (_42423_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_42424_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_42425_, _42424_, _42203_);
  nand (_42426_, _42177_, _42167_);
  and (_42427_, _42426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_42428_, _42426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_42429_, _42428_, _42199_);
  or (_42430_, _42429_, _42427_);
  or (_42431_, _42430_, _42425_);
  nand (_42432_, _42431_, _42423_);
  nand (_42433_, _42432_, _42390_);
  nand (_42434_, _42169_, _38786_);
  and (_42435_, _42434_, _42433_);
  or (_42436_, _42435_, _42171_);
  or (_42437_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_42438_, _42437_, _43223_);
  and (_02159_, _42438_, _42436_);
  and (_42439_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_42440_, _42439_, _42203_);
  nand (_42441_, _42178_, _42167_);
  and (_42442_, _42441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_42443_, _42441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_42444_, _42443_, _42199_);
  or (_42445_, _42444_, _42442_);
  or (_42446_, _42445_, _42440_);
  nor (_42447_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_42448_, _42447_, _42169_);
  and (_42449_, _42448_, _42446_);
  nor (_42450_, _42390_, _38778_);
  or (_42451_, _42450_, _42449_);
  or (_42452_, _42451_, _42195_);
  or (_42453_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_42454_, _42453_, _43223_);
  and (_02161_, _42454_, _42452_);
  nor (_42455_, _42390_, _38770_);
  and (_42456_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_42457_, _42456_, _42203_);
  and (_42458_, _42179_, _42167_);
  nor (_42459_, _42458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_42460_, _42459_, _42205_);
  or (_42461_, _42460_, _42199_);
  or (_42462_, _42461_, _42457_);
  nor (_42463_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_42464_, _42463_, _42169_);
  and (_42465_, _42464_, _42462_);
  or (_42466_, _42465_, _42195_);
  or (_42467_, _42466_, _42455_);
  or (_42468_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_42469_, _42468_, _43223_);
  and (_02163_, _42469_, _42467_);
  not (_42470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_42471_, _42143_, _42470_);
  and (_42472_, _42471_, _42203_);
  nand (_42473_, _42207_, _42314_);
  or (_42474_, _42207_, _42314_);
  and (_42475_, _42474_, _42473_);
  or (_42476_, _42475_, _42199_);
  or (_42477_, _42476_, _42472_);
  and (_42478_, _42199_, _42470_);
  nor (_42479_, _42478_, _42169_);
  and (_42480_, _42479_, _42477_);
  and (_42481_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_42482_, _42481_, _42195_);
  or (_42483_, _42482_, _42480_);
  nand (_42484_, _42171_, _38816_);
  and (_42485_, _42484_, _43223_);
  and (_02164_, _42485_, _42483_);
  and (_42486_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_42487_, _42486_, _42203_);
  nand (_42488_, _42474_, _42322_);
  or (_42489_, _42474_, _42322_);
  and (_42490_, _42489_, _42488_);
  or (_42491_, _42490_, _42199_);
  or (_42492_, _42491_, _42487_);
  nor (_42493_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_42494_, _42493_, _42169_);
  and (_42495_, _42494_, _42492_);
  and (_42496_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_42497_, _42496_, _42195_);
  or (_42498_, _42497_, _42495_);
  nand (_42499_, _42195_, _38808_);
  and (_42500_, _42499_, _43223_);
  and (_02166_, _42500_, _42498_);
  and (_42501_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_42502_, _42501_, _42203_);
  nand (_42503_, _42183_, _42167_);
  and (_42504_, _42503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_42505_, _42503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_42506_, _42505_, _42199_);
  or (_42507_, _42506_, _42504_);
  or (_42508_, _42507_, _42502_);
  nor (_42509_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_42510_, _42509_, _42169_);
  and (_42511_, _42510_, _42508_);
  and (_42512_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_42513_, _42512_, _42195_);
  or (_42514_, _42513_, _42511_);
  nand (_42515_, _42195_, _38801_);
  and (_42516_, _42515_, _43223_);
  and (_02168_, _42516_, _42514_);
  and (_42517_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_42518_, _42517_, _42203_);
  nand (_42519_, _42184_, _42167_);
  and (_42520_, _42519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_42521_, _42519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42522_, _42521_, _42199_);
  or (_42523_, _42522_, _42520_);
  or (_42524_, _42523_, _42518_);
  nor (_42525_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_42526_, _42525_, _42169_);
  and (_42527_, _42526_, _42524_);
  and (_42528_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_42529_, _42528_, _42195_);
  or (_42530_, _42529_, _42527_);
  nand (_42531_, _42195_, _38793_);
  and (_42532_, _42531_, _43223_);
  and (_02170_, _42532_, _42530_);
  and (_42533_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_42534_, _42533_, _42203_);
  nand (_42535_, _42185_, _42167_);
  and (_42536_, _42535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_42537_, _42535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42538_, _42537_, _42199_);
  or (_42539_, _42538_, _42536_);
  or (_42540_, _42539_, _42534_);
  nor (_42541_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_42542_, _42541_, _42169_);
  and (_42543_, _42542_, _42540_);
  and (_42544_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_42545_, _42544_, _42195_);
  or (_42546_, _42545_, _42543_);
  nand (_42547_, _42195_, _38786_);
  and (_42548_, _42547_, _43223_);
  and (_02171_, _42548_, _42546_);
  and (_42549_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_42550_, _42549_, _42203_);
  nand (_42551_, _42186_, _42167_);
  and (_42552_, _42551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_42553_, _42551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_42554_, _42553_, _42199_);
  or (_42555_, _42554_, _42552_);
  or (_42556_, _42555_, _42550_);
  nor (_42557_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_42558_, _42557_, _42169_);
  and (_42559_, _42558_, _42556_);
  and (_42560_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_42561_, _42560_, _42195_);
  or (_42562_, _42561_, _42559_);
  nand (_42563_, _42195_, _38778_);
  and (_42564_, _42563_, _43223_);
  and (_02173_, _42564_, _42562_);
  and (_42565_, _42373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_42566_, _42565_, _42203_);
  and (_42567_, _42187_, _42167_);
  nor (_42568_, _42567_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_42569_, _42568_, _42218_);
  or (_42570_, _42569_, _42199_);
  or (_42571_, _42570_, _42566_);
  nor (_42572_, _42201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_42573_, _42572_, _42169_);
  and (_42574_, _42573_, _42571_);
  and (_42575_, _42169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_42576_, _42575_, _42195_);
  or (_42577_, _42576_, _42574_);
  nand (_42578_, _42195_, _38770_);
  and (_42579_, _42578_, _43223_);
  and (_02175_, _42579_, _42577_);
  not (_42580_, _42244_);
  and (_42581_, _42237_, _27624_);
  or (_42582_, _42581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_42583_, _42582_, _42580_);
  nand (_42584_, _42581_, _31849_);
  and (_42585_, _42584_, _42583_);
  and (_42586_, _42244_, _38817_);
  or (_42587_, _42586_, _42585_);
  and (_02177_, _42587_, _43223_);
  and (_42588_, _42237_, _33199_);
  or (_42589_, _42588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_42590_, _42589_, _42580_);
  nand (_42591_, _42588_, _31849_);
  and (_42592_, _42591_, _42590_);
  nor (_42593_, _42580_, _38808_);
  or (_42594_, _42593_, _42592_);
  and (_02178_, _42594_, _43223_);
  nand (_42595_, _42237_, _39846_);
  and (_42596_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_42597_, _42596_, _42244_);
  and (_42598_, _33983_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_42599_, _42598_, _33972_);
  and (_42600_, _42599_, _42237_);
  or (_42601_, _42600_, _42597_);
  nand (_42602_, _42244_, _38801_);
  and (_42603_, _42602_, _43223_);
  and (_02179_, _42603_, _42601_);
  and (_42604_, _42237_, _34690_);
  or (_42605_, _42604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_42606_, _42605_, _42580_);
  nand (_42607_, _42604_, _31849_);
  and (_42608_, _42607_, _42606_);
  nor (_42609_, _42580_, _38793_);
  or (_42610_, _42609_, _42608_);
  and (_02180_, _42610_, _43223_);
  and (_42611_, _42237_, _35375_);
  or (_42612_, _42611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_42613_, _42612_, _42580_);
  nand (_42614_, _42611_, _31849_);
  and (_42615_, _42614_, _42613_);
  nor (_42616_, _42580_, _38786_);
  or (_42617_, _42616_, _42615_);
  and (_02181_, _42617_, _43223_);
  and (_42618_, _42237_, _36171_);
  or (_42619_, _42618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_42620_, _42619_, _42580_);
  nand (_42621_, _42618_, _31849_);
  and (_42622_, _42621_, _42620_);
  nor (_42623_, _42580_, _38778_);
  or (_42624_, _42623_, _42622_);
  and (_02182_, _42624_, _43223_);
  not (_42625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42626_, _42141_, _42625_);
  or (_42627_, _42626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_42628_, _42627_, _42237_);
  nand (_42629_, _39387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_42630_, _42629_, _42237_);
  or (_42631_, _42630_, _39388_);
  and (_42632_, _42631_, _42628_);
  or (_42633_, _42632_, _42244_);
  nand (_42634_, _42244_, _38770_);
  and (_42635_, _42634_, _43223_);
  and (_02184_, _42635_, _42633_);
  and (_42636_, _31238_, _28106_);
  and (_42637_, _38839_, _38749_);
  not (_42638_, _42637_);
  not (_42639_, _38612_);
  not (_42640_, _38748_);
  nor (_42641_, _42640_, _38714_);
  not (_42642_, _37083_);
  and (_42643_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_42644_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42645_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_42646_, _42645_, _42644_);
  and (_42647_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_42648_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_42649_, _42648_, _42647_);
  and (_42650_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_42651_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42652_, _42651_, _42650_);
  and (_42653_, _42652_, _42649_);
  and (_42654_, _42653_, _42646_);
  nor (_42655_, _37269_, _42642_);
  not (_42656_, _42655_);
  nor (_42657_, _42656_, _42654_);
  nor (_42658_, _42657_, _42643_);
  not (_42659_, _42658_);
  and (_42660_, _42659_, _42641_);
  nor (_42661_, _42660_, _42639_);
  and (_42662_, _42640_, _38714_);
  nor (_42663_, _39239_, _39328_);
  nor (_42664_, _42663_, _39334_);
  nor (_42665_, _42664_, _28293_);
  and (_42666_, _42664_, _28293_);
  or (_42667_, _42666_, _42665_);
  not (_42668_, _42667_);
  nor (_42669_, _38504_, _27602_);
  and (_42670_, _38504_, _27602_);
  nor (_42671_, _42670_, _42669_);
  and (_42672_, _27821_, _28128_);
  not (_42673_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_42674_, _31238_, _42673_);
  and (_42675_, _42674_, _33983_);
  and (_42676_, _42675_, _42672_);
  and (_42677_, _42676_, _42671_);
  and (_42678_, _42677_, _27953_);
  not (_42679_, _28424_);
  and (_42680_, _39342_, _42679_);
  nor (_42681_, _39342_, _42679_);
  nor (_42682_, _42681_, _42680_);
  and (_42683_, _42682_, _42678_);
  and (_42684_, _42683_, _42668_);
  not (_42685_, _39342_);
  nor (_42686_, _42664_, _38639_);
  and (_42687_, _42686_, _42685_);
  and (_42688_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor (_42689_, _42664_, _38504_);
  and (_42690_, _42689_, _42685_);
  and (_42691_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_42692_, _42691_, _42688_);
  and (_42693_, _42664_, _38504_);
  and (_42694_, _42693_, _39342_);
  and (_42695_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_42696_, _42693_, _42685_);
  and (_42697_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_42698_, _42697_, _42695_);
  and (_42699_, _42698_, _42692_);
  and (_42700_, _42664_, _38639_);
  and (_42701_, _42700_, _39342_);
  and (_42702_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_42703_, _42686_, _39342_);
  and (_42704_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_42705_, _42704_, _42702_);
  and (_42706_, _42689_, _39342_);
  and (_42707_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_42708_, _42700_, _42685_);
  and (_42709_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_42710_, _42709_, _42707_);
  and (_42711_, _42710_, _42705_);
  and (_42712_, _42711_, _42699_);
  nor (_42713_, _42712_, _42684_);
  not (_42714_, _38837_);
  and (_42715_, _42684_, _42714_);
  nor (_42716_, _42715_, _42713_);
  not (_42717_, _42716_);
  and (_42718_, _42717_, _42662_);
  not (_42719_, _42718_);
  and (_42720_, _42719_, _42661_);
  and (_42721_, _42720_, _42638_);
  not (_42722_, _38688_);
  and (_42723_, _42722_, _38682_);
  nor (_42724_, _38677_, _38673_);
  nor (_42725_, _38685_, _38670_);
  and (_42726_, _42725_, _38660_);
  and (_42727_, _42726_, _42724_);
  and (_42728_, _42727_, _42723_);
  nor (_42729_, _42728_, _37039_);
  not (_42730_, _42729_);
  or (_42731_, _38692_, _38667_);
  and (_42732_, _42731_, _38602_);
  and (_42733_, _38600_, _42732_);
  nor (_42734_, _38699_, _37039_);
  nor (_42735_, _42734_, _42733_);
  and (_42736_, _42735_, _42730_);
  not (_42737_, _42736_);
  and (_42738_, _42737_, _42721_);
  and (_42739_, _42641_, _38612_);
  and (_42740_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_42741_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42742_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_42743_, _42742_, _42741_);
  and (_42744_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_42745_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42746_, _42745_, _42744_);
  and (_42747_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_42748_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_42749_, _42748_, _42747_);
  and (_42750_, _42749_, _42746_);
  and (_42751_, _42750_, _42743_);
  nor (_42752_, _42751_, _42656_);
  nor (_42753_, _42752_, _42740_);
  not (_42754_, _42753_);
  and (_42755_, _42754_, _42739_);
  and (_42756_, _38748_, _38714_);
  and (_42757_, _42756_, _38612_);
  and (_42758_, _42757_, _42685_);
  nor (_42759_, _42758_, _42755_);
  and (_42760_, _42662_, _38612_);
  and (_42761_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_42762_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_42763_, _42762_, _42761_);
  and (_42764_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_42765_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_42766_, _42765_, _42764_);
  and (_42767_, _42766_, _42763_);
  and (_42768_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_42769_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_42770_, _42769_, _42768_);
  and (_42771_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_42772_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_42773_, _42772_, _42771_);
  and (_42774_, _42773_, _42770_);
  and (_42775_, _42774_, _42767_);
  nor (_42776_, _42775_, _42684_);
  not (_42777_, _38786_);
  and (_42778_, _42684_, _42777_);
  nor (_42779_, _42778_, _42776_);
  not (_42780_, _42779_);
  and (_42781_, _42780_, _42760_);
  not (_42782_, _42781_);
  not (_42783_, _38871_);
  and (_42784_, _42783_, _38750_);
  and (_42785_, _42639_, _38748_);
  nor (_42786_, _42785_, _42784_);
  and (_42787_, _42786_, _42782_);
  and (_42788_, _42787_, _42759_);
  not (_42789_, _42788_);
  and (_42790_, _42789_, _42738_);
  and (_42791_, _42662_, _42639_);
  and (_42792_, _42757_, _38527_);
  or (_42793_, _42792_, _42791_);
  and (_42794_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_42795_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_42796_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_42797_, _42796_, _42795_);
  and (_42798_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42799_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42800_, _42799_, _42798_);
  and (_42801_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_42802_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_42803_, _42802_, _42801_);
  and (_42804_, _42803_, _42800_);
  and (_42805_, _42804_, _42797_);
  nor (_42806_, _42805_, _42656_);
  nor (_42807_, _42806_, _42794_);
  not (_42808_, _42807_);
  and (_42809_, _42808_, _42739_);
  not (_42810_, _38853_);
  and (_42811_, _42810_, _38750_);
  and (_42812_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_42813_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_42814_, _42813_, _42812_);
  and (_42815_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_42816_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_42817_, _42816_, _42815_);
  and (_42818_, _42817_, _42814_);
  and (_42819_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_42820_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_42821_, _42820_, _42819_);
  and (_42822_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_42823_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_42824_, _42823_, _42822_);
  and (_42825_, _42824_, _42821_);
  and (_42826_, _42825_, _42818_);
  nor (_42827_, _42826_, _42684_);
  not (_42828_, _38808_);
  and (_42829_, _42684_, _42828_);
  nor (_42830_, _42829_, _42827_);
  not (_42831_, _42830_);
  and (_42832_, _42831_, _42760_);
  or (_42833_, _42832_, _42811_);
  or (_42834_, _42833_, _42809_);
  nor (_42835_, _42834_, _42793_);
  nor (_42836_, _42835_, _42737_);
  nor (_42837_, _42836_, _42790_);
  and (_42838_, _28128_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42839_, _42838_, _42679_);
  nor (_42840_, _27481_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42841_, _42840_, _42839_);
  nand (_42842_, _42841_, _42837_);
  or (_42843_, _42841_, _42837_);
  and (_42844_, _42843_, _42842_);
  and (_42845_, _42838_, _28293_);
  nor (_42846_, _27602_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42847_, _42846_, _42845_);
  not (_42848_, _42847_);
  not (_42849_, _38865_);
  and (_42850_, _42849_, _38750_);
  and (_42851_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_42852_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_42853_, _42852_, _42851_);
  and (_42854_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_42855_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_42856_, _42855_, _42854_);
  and (_42857_, _42856_, _42853_);
  and (_42858_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_42859_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_42860_, _42859_, _42858_);
  and (_42861_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_42862_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_42863_, _42862_, _42861_);
  and (_42864_, _42863_, _42860_);
  and (_42865_, _42864_, _42857_);
  nor (_42866_, _42865_, _42684_);
  not (_42867_, _38793_);
  and (_42868_, _42684_, _42867_);
  nor (_42869_, _42868_, _42866_);
  not (_42870_, _42869_);
  and (_42871_, _42870_, _42760_);
  nor (_42872_, _42871_, _42850_);
  not (_42873_, _42664_);
  and (_42874_, _42757_, _42873_);
  and (_42875_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_42876_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42877_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_42878_, _42877_, _42876_);
  and (_42879_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_42880_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_42881_, _42880_, _42879_);
  and (_42882_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_42883_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42884_, _42883_, _42882_);
  and (_42885_, _42884_, _42881_);
  and (_42886_, _42885_, _42878_);
  nor (_42887_, _42886_, _42656_);
  nor (_42888_, _42887_, _42875_);
  not (_42889_, _42888_);
  and (_42890_, _42889_, _42739_);
  nor (_42891_, _42890_, _42874_);
  and (_42892_, _42891_, _42872_);
  not (_42893_, _42892_);
  and (_42894_, _42893_, _42738_);
  not (_42895_, _38847_);
  and (_42896_, _42895_, _38750_);
  and (_42897_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_42898_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_42899_, _42898_, _42897_);
  and (_42900_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_42901_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_42902_, _42901_, _42900_);
  and (_42903_, _42902_, _42899_);
  and (_42904_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_42905_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_42906_, _42905_, _42904_);
  and (_42907_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_42908_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_42909_, _42908_, _42907_);
  and (_42910_, _42909_, _42906_);
  and (_42911_, _42910_, _42903_);
  nor (_42912_, _42911_, _42684_);
  and (_42913_, _42684_, _38817_);
  nor (_42914_, _42913_, _42912_);
  not (_42915_, _42914_);
  and (_42916_, _42915_, _42760_);
  nor (_42917_, _42916_, _42896_);
  and (_42918_, _42757_, _38504_);
  and (_42919_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_42920_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42921_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_42922_, _42921_, _42920_);
  and (_42923_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_42924_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_42925_, _42924_, _42923_);
  and (_42926_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_42927_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42928_, _42927_, _42926_);
  and (_42929_, _42928_, _42925_);
  and (_42930_, _42929_, _42922_);
  nor (_42931_, _42930_, _42656_);
  nor (_42932_, _42931_, _42919_);
  not (_42933_, _42932_);
  and (_42934_, _42933_, _42739_);
  nor (_42935_, _42934_, _42918_);
  and (_42936_, _42935_, _42917_);
  nor (_42937_, _42936_, _42737_);
  nor (_42938_, _42937_, _42894_);
  and (_42939_, _42938_, _42848_);
  nor (_42940_, _42938_, _42848_);
  nor (_42941_, _42940_, _42939_);
  not (_42942_, _42941_);
  nor (_42943_, _42942_, _42844_);
  and (_42944_, _42838_, _38754_);
  nor (_42945_, _42838_, _28282_);
  nor (_42946_, _42945_, _42944_);
  nor (_42947_, _42662_, _38612_);
  and (_42948_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_42949_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_42950_, _42949_, _42948_);
  and (_42951_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_42952_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_42953_, _42952_, _42951_);
  and (_42954_, _42953_, _42950_);
  and (_42955_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_42956_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_42957_, _42956_, _42955_);
  and (_42958_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_42959_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_42960_, _42959_, _42958_);
  and (_42961_, _42960_, _42957_);
  and (_42962_, _42961_, _42954_);
  nor (_42963_, _42962_, _42684_);
  not (_42964_, _38770_);
  and (_42965_, _42684_, _42964_);
  nor (_42966_, _42965_, _42963_);
  not (_42967_, _42966_);
  and (_42968_, _42967_, _42760_);
  nor (_42969_, _42968_, _42947_);
  not (_42970_, _38883_);
  and (_42971_, _42970_, _38750_);
  and (_42972_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_42973_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42974_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_42975_, _42974_, _42973_);
  and (_42976_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_42977_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_42978_, _42977_, _42976_);
  and (_42979_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_42980_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42981_, _42980_, _42979_);
  and (_42982_, _42981_, _42978_);
  and (_42983_, _42982_, _42975_);
  nor (_42984_, _42983_, _42656_);
  nor (_42985_, _42984_, _42972_);
  not (_42986_, _42985_);
  and (_42987_, _42986_, _42739_);
  nor (_42988_, _42987_, _42971_);
  and (_42989_, _42988_, _42969_);
  and (_42990_, _42989_, _42738_);
  nor (_42991_, _42893_, _42738_);
  nor (_42992_, _42991_, _42990_);
  nor (_42993_, _42992_, _42946_);
  and (_42994_, _42992_, _42946_);
  nor (_42995_, _42994_, _42993_);
  and (_42996_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_42997_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42998_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_42999_, _42998_, _42997_);
  and (_43000_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_43001_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_43002_, _43001_, _43000_);
  and (_43003_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_43004_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_43005_, _43004_, _43003_);
  and (_43006_, _43005_, _43002_);
  and (_43007_, _43006_, _42999_);
  nor (_43008_, _43007_, _42656_);
  nor (_43009_, _43008_, _42996_);
  not (_43010_, _43009_);
  and (_43011_, _43010_, _42739_);
  and (_43012_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_43013_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_43014_, _43013_, _43012_);
  and (_43015_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_43016_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_43017_, _43016_, _43015_);
  and (_43018_, _43017_, _43014_);
  and (_43019_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_43020_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_43021_, _43020_, _43019_);
  and (_43022_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_43023_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_43024_, _43023_, _43022_);
  and (_43025_, _43024_, _43021_);
  and (_43026_, _43025_, _43018_);
  nor (_43027_, _43026_, _42684_);
  not (_43028_, _38778_);
  and (_43029_, _42684_, _43028_);
  nor (_43030_, _43029_, _43027_);
  not (_43031_, _43030_);
  and (_43032_, _43031_, _42760_);
  nor (_43033_, _43032_, _43011_);
  nor (_43034_, _38877_, _38748_);
  nor (_43035_, _43034_, _42639_);
  or (_43036_, _42641_, _42662_);
  nor (_43037_, _43036_, _43035_);
  not (_43038_, _43037_);
  and (_43039_, _43038_, _43033_);
  not (_43040_, _43039_);
  and (_43041_, _43040_, _42738_);
  and (_43042_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_43043_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_43044_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_43045_, _43044_, _43043_);
  and (_43046_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_43047_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_43048_, _43047_, _43046_);
  and (_43049_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_43050_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_43051_, _43050_, _43049_);
  and (_43052_, _43051_, _43048_);
  and (_43053_, _43052_, _43045_);
  nor (_43054_, _43053_, _42656_);
  nor (_43055_, _43054_, _43042_);
  not (_43056_, _43055_);
  and (_43057_, _43056_, _42739_);
  and (_43058_, _42706_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_43059_, _42701_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_43060_, _43059_, _43058_);
  and (_43061_, _42696_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_43062_, _42687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_43063_, _43062_, _43061_);
  and (_43064_, _43063_, _43060_);
  and (_43065_, _42703_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_43066_, _42708_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_43067_, _43066_, _43065_);
  and (_43068_, _42690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_43069_, _42694_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_43070_, _43069_, _43068_);
  and (_43071_, _43070_, _43067_);
  and (_43072_, _43071_, _43064_);
  nor (_43073_, _43072_, _42684_);
  not (_43074_, _38801_);
  and (_43075_, _42684_, _43074_);
  nor (_43076_, _43075_, _43073_);
  not (_43077_, _43076_);
  and (_43078_, _43077_, _42760_);
  nor (_43079_, _43078_, _43057_);
  not (_43080_, _38859_);
  and (_43081_, _43080_, _38750_);
  and (_43082_, _42757_, _38548_);
  nor (_43083_, _43082_, _43081_);
  and (_43084_, _43083_, _43079_);
  nor (_43085_, _43084_, _42737_);
  nor (_43086_, _43085_, _43041_);
  and (_43087_, _42838_, _39234_);
  nor (_43088_, _27361_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_43089_, _43088_, _43087_);
  not (_43090_, _43089_);
  nor (_43091_, _43090_, _43086_);
  and (_43092_, _43090_, _43086_);
  nor (_43093_, _43092_, _43091_);
  and (_43094_, _43093_, _42995_);
  and (_43095_, _43094_, _42943_);
  and (_43096_, _43095_, _42636_);
  nor (_43097_, _42989_, _42738_);
  nor (_43098_, _42838_, _27821_);
  not (_43099_, _43098_);
  nor (_43100_, _43099_, _43097_);
  nor (_43101_, _43040_, _42738_);
  nor (_43102_, _42838_, _39234_);
  not (_43103_, _43102_);
  and (_43104_, _43103_, _43101_);
  and (_43105_, _43099_, _43097_);
  or (_43106_, _43105_, _43104_);
  or (_43107_, _43106_, _43100_);
  nor (_43108_, _42788_, _42738_);
  nor (_43109_, _42838_, _28424_);
  not (_43110_, _43109_);
  and (_43111_, _43110_, _43108_);
  nor (_43112_, _43110_, _43108_);
  nor (_43113_, _43112_, _43111_);
  nor (_43114_, _43103_, _43101_);
  nor (_43115_, _42721_, _28128_);
  and (_43116_, _42721_, _28128_);
  nor (_43117_, _43116_, _43115_);
  nor (_43118_, _43117_, _43114_);
  nand (_43119_, _43118_, _43113_);
  nor (_43120_, _43119_, _43107_);
  and (_43121_, _43120_, _43096_);
  not (_43122_, _43086_);
  not (_43123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_43124_, _42938_, _43123_);
  and (_43125_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_43126_, _43125_, _42837_);
  or (_43127_, _43126_, _43124_);
  and (_43128_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_43129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_43130_, _42938_, _43129_);
  nand (_43131_, _43130_, _42837_);
  or (_43132_, _43131_, _43128_);
  and (_43133_, _43132_, _43127_);
  or (_43134_, _43133_, _43122_);
  not (_43135_, _42992_);
  not (_43136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_43137_, _42938_, _43136_);
  and (_43138_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_43139_, _43138_, _42837_);
  or (_43140_, _43139_, _43137_);
  and (_43141_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_43142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_43143_, _42938_, _43142_);
  nand (_43144_, _43143_, _42837_);
  or (_43145_, _43144_, _43141_);
  and (_43146_, _43145_, _43140_);
  or (_43147_, _43146_, _43086_);
  and (_43148_, _43147_, _43135_);
  and (_43149_, _43148_, _43134_);
  not (_43150_, _42837_);
  not (_43151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_43152_, _42938_, _43151_);
  or (_43153_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_43154_, _43153_, _43152_);
  or (_43155_, _43154_, _43150_);
  or (_43156_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_43157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_43158_, _42938_, _43157_);
  and (_43159_, _43158_, _43156_);
  or (_43161_, _43159_, _42837_);
  and (_43162_, _43161_, _43155_);
  or (_43164_, _43162_, _43122_);
  not (_43166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_43167_, _42938_, _43166_);
  or (_43169_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_43171_, _43169_, _43167_);
  or (_43173_, _43171_, _43150_);
  or (_43175_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_43176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_43177_, _42938_, _43176_);
  and (_43178_, _43177_, _43175_);
  or (_43179_, _43178_, _42837_);
  and (_43180_, _43179_, _43173_);
  or (_43181_, _43180_, _43086_);
  and (_43182_, _43181_, _42992_);
  and (_43183_, _43182_, _43164_);
  or (_43184_, _43183_, _43149_);
  or (_43185_, _43184_, _43121_);
  not (_43186_, _43121_);
  or (_43187_, _43186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_43188_, _43096_);
  nor (_43189_, _43121_, _43188_);
  nor (_43190_, _43189_, rst);
  and (_43191_, _43190_, _43187_);
  and (_43192_, _43191_, _43185_);
  and (_43193_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_43194_, _43193_, _29269_);
  nor (_43195_, _43194_, _31849_);
  nor (_43196_, _38837_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43197_, _29269_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_43198_, _20627_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43199_, _43198_, _43197_);
  or (_43200_, _43199_, _43196_);
  or (_43201_, _43200_, _43195_);
  and (_40450_, _43201_, _43223_);
  and (_43202_, _40450_, _43189_);
  or (_02560_, _43202_, _43192_);
  not (_43203_, _42636_);
  nor (_43204_, _42847_, _43203_);
  nor (_43205_, _43203_, _42841_);
  and (_43206_, _43205_, _43204_);
  nor (_43207_, _42946_, _43203_);
  nor (_43208_, _43203_, _43089_);
  and (_43209_, _43208_, _43207_);
  and (_43211_, _43209_, _43206_);
  and (_43213_, _43201_, _42636_);
  and (_43215_, _43213_, _43211_);
  not (_43217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_43219_, _43211_, _43217_);
  or (_02571_, _43219_, _43215_);
  nor (_43222_, _43208_, _43207_);
  nor (_43224_, _43205_, _43204_);
  and (_43225_, _43224_, _42636_);
  and (_43227_, _43225_, _43222_);
  and (_43229_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _29345_);
  and (_43230_, _43229_, _29291_);
  nand (_43231_, _43230_, _31849_);
  not (_43232_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43233_, _38816_, _43232_);
  or (_43234_, _19467_, _43232_);
  and (_43235_, _43234_, _43233_);
  or (_43236_, _43235_, _43230_);
  and (_43237_, _43236_, _43231_);
  and (_43238_, _43237_, _43227_);
  not (_43239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_43240_, _43227_, _43239_);
  or (_02806_, _43240_, _43238_);
  nand (_43241_, _43229_, _29236_);
  nor (_43242_, _43241_, _31849_);
  nor (_43243_, _38808_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43244_, _43229_, _29181_);
  and (_43245_, _43229_, _29269_);
  or (_43246_, _43245_, _43193_);
  or (_43247_, _43246_, _43244_);
  and (_43248_, _43247_, _20453_);
  or (_43249_, _43248_, _43243_);
  or (_43250_, _43249_, _43242_);
  and (_43251_, _43250_, _43227_);
  not (_43252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_43253_, _43227_, _43252_);
  or (_02811_, _43253_, _43251_);
  not (_43254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_43255_, _43227_, _43254_);
  nand (_43256_, _43229_, _29192_);
  nor (_43257_, _43256_, _31849_);
  nor (_43258_, _38801_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43259_, _43229_, _29225_);
  or (_43260_, _43259_, _43246_);
  and (_43261_, _43260_, _19106_);
  or (_43262_, _43261_, _43258_);
  or (_43263_, _43262_, _43257_);
  and (_43264_, _43263_, _43227_);
  or (_02816_, _43264_, _43255_);
  and (_43265_, _43245_, _32481_);
  nor (_43266_, _38793_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_43267_, _43244_, _43193_);
  or (_43268_, _43267_, _43259_);
  and (_43269_, _43268_, _20137_);
  or (_43270_, _43269_, _43266_);
  or (_43271_, _43270_, _43265_);
  and (_43272_, _43271_, _43227_);
  not (_43273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_43274_, _43227_, _43273_);
  or (_02820_, _43274_, _43272_);
  nand (_43275_, _43193_, _29291_);
  nor (_43276_, _43275_, _31849_);
  nor (_43277_, _38786_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43278_, _29291_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_43279_, _19304_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43280_, _43279_, _43278_);
  or (_43281_, _43280_, _43277_);
  or (_43282_, _43281_, _43276_);
  and (_43283_, _43282_, _43227_);
  not (_43284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_43285_, _43227_, _43284_);
  or (_02825_, _43285_, _43283_);
  not (_43286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_43287_, _43227_, _43286_);
  nand (_43288_, _43193_, _29236_);
  nor (_43289_, _43288_, _31849_);
  nor (_43290_, _38778_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43291_, _29236_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_43292_, _20290_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43293_, _43292_, _43291_);
  or (_43294_, _43293_, _43290_);
  or (_43295_, _43294_, _43289_);
  and (_43296_, _43295_, _43227_);
  or (_02830_, _43296_, _43287_);
  nand (_43297_, _43193_, _29192_);
  nor (_43298_, _43297_, _31849_);
  nor (_43299_, _38770_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_43300_, _29192_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_43301_, _19641_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_43302_, _43301_, _43300_);
  or (_43303_, _43302_, _43299_);
  or (_43304_, _43303_, _43298_);
  and (_43305_, _43304_, _43227_);
  not (_43306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_43307_, _43227_, _43306_);
  or (_02835_, _43307_, _43305_);
  not (_43308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_43309_, _43227_, _43308_);
  and (_43310_, _43227_, _43201_);
  or (_02837_, _43310_, _43309_);
  and (_43311_, _43237_, _42636_);
  and (_43312_, _43204_, _42841_);
  and (_43313_, _43312_, _43222_);
  and (_43314_, _43313_, _43311_);
  not (_43315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_43316_, _43313_, _43315_);
  or (_02844_, _43316_, _43314_);
  and (_43317_, _43250_, _42636_);
  and (_43318_, _43313_, _43317_);
  not (_43319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_43320_, _43313_, _43319_);
  or (_02848_, _43320_, _43318_);
  and (_43321_, _43263_, _42636_);
  and (_43322_, _43313_, _43321_);
  not (_43323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_43324_, _43313_, _43323_);
  or (_02851_, _43324_, _43322_);
  and (_43325_, _43271_, _42636_);
  and (_43326_, _43313_, _43325_);
  not (_43327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_43328_, _43313_, _43327_);
  or (_02855_, _43328_, _43326_);
  and (_43329_, _43282_, _42636_);
  and (_43330_, _43313_, _43329_);
  not (_43331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_43332_, _43313_, _43331_);
  or (_02858_, _43332_, _43330_);
  and (_43333_, _43295_, _42636_);
  and (_43334_, _43313_, _43333_);
  not (_43335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_43336_, _43313_, _43335_);
  or (_02862_, _43336_, _43334_);
  and (_43337_, _43304_, _42636_);
  and (_43338_, _43313_, _43337_);
  not (_43339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_43340_, _43313_, _43339_);
  or (_02865_, _43340_, _43338_);
  and (_43341_, _43313_, _43213_);
  nor (_43342_, _43313_, _43129_);
  or (_02867_, _43342_, _43341_);
  and (_43343_, _43205_, _42847_);
  and (_43344_, _43343_, _43222_);
  and (_43345_, _43344_, _43311_);
  not (_43346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_43347_, _43344_, _43346_);
  or (_02874_, _43347_, _43345_);
  and (_43348_, _43344_, _43317_);
  not (_43349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_43350_, _43344_, _43349_);
  or (_02878_, _43350_, _43348_);
  and (_43351_, _43344_, _43321_);
  not (_43352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_43353_, _43344_, _43352_);
  or (_02882_, _43353_, _43351_);
  and (_43354_, _43344_, _43325_);
  not (_43355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_43356_, _43344_, _43355_);
  or (_02885_, _43356_, _43354_);
  and (_43357_, _43344_, _43329_);
  not (_43358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_43359_, _43344_, _43358_);
  or (_02890_, _43359_, _43357_);
  and (_43360_, _43344_, _43333_);
  not (_43361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_43362_, _43344_, _43361_);
  or (_02893_, _43362_, _43360_);
  and (_43363_, _43344_, _43337_);
  not (_43364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_43365_, _43344_, _43364_);
  or (_02897_, _43365_, _43363_);
  and (_43366_, _43344_, _43213_);
  not (_43367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_43368_, _43344_, _43367_);
  or (_02900_, _43368_, _43366_);
  and (_43369_, _43222_, _43206_);
  and (_43370_, _43369_, _43311_);
  not (_43371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_43372_, _43369_, _43371_);
  or (_02906_, _43372_, _43370_);
  and (_43373_, _43369_, _43317_);
  not (_43374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_43375_, _43369_, _43374_);
  or (_02910_, _43375_, _43373_);
  and (_43376_, _43369_, _43321_);
  not (_43377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_43378_, _43369_, _43377_);
  or (_02913_, _43378_, _43376_);
  and (_43379_, _43369_, _43325_);
  not (_43380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_43381_, _43369_, _43380_);
  or (_02917_, _43381_, _43379_);
  and (_43382_, _43369_, _43329_);
  not (_43383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_43384_, _43369_, _43383_);
  or (_02920_, _43384_, _43382_);
  and (_43385_, _43369_, _43333_);
  not (_43386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_43387_, _43369_, _43386_);
  or (_02924_, _43387_, _43385_);
  and (_43388_, _43369_, _43337_);
  not (_43389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_43390_, _43369_, _43389_);
  or (_02928_, _43390_, _43388_);
  and (_43391_, _43369_, _43213_);
  nor (_43392_, _43369_, _43123_);
  or (_02931_, _43392_, _43391_);
  and (_43393_, _43208_, _42946_);
  and (_43394_, _43393_, _43224_);
  and (_43395_, _43394_, _43311_);
  not (_43396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_43397_, _43394_, _43396_);
  or (_02939_, _43397_, _43395_);
  and (_43398_, _43394_, _43317_);
  not (_43399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_43400_, _43394_, _43399_);
  or (_02943_, _43400_, _43398_);
  and (_43401_, _43394_, _43321_);
  not (_43402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_43403_, _43394_, _43402_);
  or (_02946_, _43403_, _43401_);
  and (_43404_, _43394_, _43325_);
  not (_43405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_43406_, _43394_, _43405_);
  or (_02950_, _43406_, _43404_);
  and (_43407_, _43394_, _43329_);
  not (_43408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_43409_, _43394_, _43408_);
  or (_02954_, _43409_, _43407_);
  and (_43410_, _43394_, _43333_);
  not (_43411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_43412_, _43394_, _43411_);
  or (_02957_, _43412_, _43410_);
  and (_43413_, _43394_, _43337_);
  not (_43414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_43415_, _43394_, _43414_);
  or (_02961_, _43415_, _43413_);
  and (_43416_, _43394_, _43213_);
  not (_43417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_43418_, _43394_, _43417_);
  or (_02964_, _43418_, _43416_);
  and (_43419_, _43393_, _43312_);
  and (_43420_, _43419_, _43311_);
  not (_43421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_43422_, _43419_, _43421_);
  or (_02969_, _43422_, _43420_);
  and (_43423_, _43419_, _43317_);
  not (_43424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_43425_, _43419_, _43424_);
  or (_02972_, _43425_, _43423_);
  and (_43426_, _43419_, _43321_);
  not (_43427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_43428_, _43419_, _43427_);
  or (_02976_, _43428_, _43426_);
  and (_43429_, _43419_, _43325_);
  not (_43430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_43431_, _43419_, _43430_);
  or (_02980_, _43431_, _43429_);
  and (_43432_, _43419_, _43329_);
  not (_43433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_43434_, _43419_, _43433_);
  or (_02983_, _43434_, _43432_);
  and (_43435_, _43419_, _43333_);
  not (_43436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_43437_, _43419_, _43436_);
  or (_02987_, _43437_, _43435_);
  and (_43438_, _43419_, _43337_);
  not (_43439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_43440_, _43419_, _43439_);
  or (_02991_, _43440_, _43438_);
  and (_43441_, _43419_, _43213_);
  nor (_43442_, _43419_, _43142_);
  or (_02993_, _43442_, _43441_);
  and (_43443_, _43393_, _43343_);
  and (_43444_, _43443_, _43311_);
  not (_43445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_43446_, _43443_, _43445_);
  or (_02997_, _43446_, _43444_);
  and (_43447_, _43443_, _43317_);
  not (_43448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_43449_, _43443_, _43448_);
  or (_03002_, _43449_, _43447_);
  and (_43450_, _43443_, _43321_);
  not (_43451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_43452_, _43443_, _43451_);
  or (_03005_, _43452_, _43450_);
  and (_43453_, _43443_, _43325_);
  not (_43454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_43455_, _43443_, _43454_);
  or (_03008_, _43455_, _43453_);
  and (_43456_, _43443_, _43329_);
  not (_43457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_43458_, _43443_, _43457_);
  or (_03012_, _43458_, _43456_);
  and (_43459_, _43443_, _43333_);
  not (_43460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_43461_, _43443_, _43460_);
  or (_03016_, _43461_, _43459_);
  and (_43462_, _43443_, _43337_);
  not (_43463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_43464_, _43443_, _43463_);
  or (_03019_, _43464_, _43462_);
  and (_43465_, _43443_, _43213_);
  not (_43466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_43467_, _43443_, _43466_);
  or (_03021_, _43467_, _43465_);
  and (_43468_, _43393_, _43206_);
  and (_43469_, _43468_, _43311_);
  not (_43470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_43471_, _43468_, _43470_);
  or (_03026_, _43471_, _43469_);
  and (_43472_, _43468_, _43317_);
  not (_43473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_43474_, _43468_, _43473_);
  or (_03030_, _43474_, _43472_);
  and (_43475_, _43468_, _43321_);
  not (_43476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_43477_, _43468_, _43476_);
  or (_03033_, _43477_, _43475_);
  and (_43478_, _43468_, _43325_);
  not (_43479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_43480_, _43468_, _43479_);
  or (_03036_, _43480_, _43478_);
  and (_43481_, _43468_, _43329_);
  not (_43482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_43483_, _43468_, _43482_);
  or (_03039_, _43483_, _43481_);
  and (_43484_, _43468_, _43333_);
  not (_43485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_43486_, _43468_, _43485_);
  or (_03043_, _43486_, _43484_);
  and (_43487_, _43468_, _43337_);
  not (_43488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_43489_, _43468_, _43488_);
  or (_03046_, _43489_, _43487_);
  and (_43490_, _43468_, _43213_);
  nor (_43491_, _43468_, _43136_);
  or (_03048_, _43491_, _43490_);
  and (_43492_, _43207_, _43089_);
  and (_43493_, _43492_, _43224_);
  and (_43494_, _43493_, _43311_);
  not (_43495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_43496_, _43493_, _43495_);
  or (_03055_, _43496_, _43494_);
  and (_43497_, _43493_, _43317_);
  not (_43498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_43499_, _43493_, _43498_);
  or (_03057_, _43499_, _43497_);
  and (_43500_, _43493_, _43321_);
  not (_43501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_43502_, _43493_, _43501_);
  or (_03061_, _43502_, _43500_);
  and (_43503_, _43493_, _43325_);
  not (_43504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_43505_, _43493_, _43504_);
  or (_03064_, _43505_, _43503_);
  and (_43506_, _43493_, _43329_);
  not (_43507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_43508_, _43493_, _43507_);
  or (_03068_, _43508_, _43506_);
  and (_43509_, _43493_, _43333_);
  not (_43510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_43511_, _43493_, _43510_);
  or (_03072_, _43511_, _43509_);
  and (_43512_, _43493_, _43337_);
  not (_43513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_43514_, _43493_, _43513_);
  or (_03076_, _43514_, _43512_);
  and (_43515_, _43493_, _43213_);
  nor (_43516_, _43493_, _43151_);
  or (_03078_, _43516_, _43515_);
  and (_43517_, _43492_, _43312_);
  and (_43518_, _43517_, _43311_);
  not (_43519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_43520_, _43517_, _43519_);
  or (_03083_, _43520_, _43518_);
  and (_43521_, _43517_, _43317_);
  not (_43522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_43523_, _43517_, _43522_);
  or (_03086_, _43523_, _43521_);
  and (_43524_, _43517_, _43321_);
  not (_43525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_43526_, _43517_, _43525_);
  or (_03090_, _43526_, _43524_);
  and (_43527_, _43517_, _43325_);
  not (_43528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_43529_, _43517_, _43528_);
  or (_03093_, _43529_, _43527_);
  and (_43530_, _43517_, _43329_);
  not (_43531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_43532_, _43517_, _43531_);
  or (_03097_, _43532_, _43530_);
  and (_43533_, _43517_, _43333_);
  not (_43534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_43535_, _43517_, _43534_);
  or (_03101_, _43535_, _43533_);
  and (_43536_, _43517_, _43337_);
  not (_43537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_43538_, _43517_, _43537_);
  or (_03104_, _43538_, _43536_);
  and (_43539_, _43517_, _43213_);
  not (_43540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_43541_, _43517_, _43540_);
  or (_03107_, _43541_, _43539_);
  and (_43542_, _43492_, _43343_);
  and (_43543_, _43542_, _43311_);
  not (_43544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_43545_, _43542_, _43544_);
  or (_03112_, _43545_, _43543_);
  and (_43546_, _43542_, _43317_);
  not (_43547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_43548_, _43542_, _43547_);
  or (_03116_, _43548_, _43546_);
  and (_43549_, _43542_, _43321_);
  not (_43550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_43551_, _43542_, _43550_);
  or (_03120_, _43551_, _43549_);
  and (_43552_, _43542_, _43325_);
  not (_43553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_43554_, _43542_, _43553_);
  or (_03124_, _43554_, _43552_);
  and (_43555_, _43542_, _43329_);
  not (_43556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_43557_, _43542_, _43556_);
  or (_03127_, _43557_, _43555_);
  and (_43558_, _43542_, _43333_);
  not (_43559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_43560_, _43542_, _43559_);
  or (_03132_, _43560_, _43558_);
  and (_43561_, _43542_, _43337_);
  not (_43562_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_43563_, _43542_, _43562_);
  or (_03136_, _43563_, _43561_);
  and (_43564_, _43542_, _43213_);
  nor (_43565_, _43542_, _43157_);
  or (_03139_, _43565_, _43564_);
  and (_43566_, _43492_, _43206_);
  and (_43567_, _43566_, _43311_);
  not (_43568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_43569_, _43566_, _43568_);
  or (_03144_, _43569_, _43567_);
  and (_43570_, _43566_, _43317_);
  not (_43571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_43572_, _43566_, _43571_);
  or (_03147_, _43572_, _43570_);
  and (_43573_, _43566_, _43321_);
  not (_43574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_43575_, _43566_, _43574_);
  or (_03151_, _43575_, _43573_);
  and (_43576_, _43566_, _43325_);
  not (_43577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_43578_, _43566_, _43577_);
  or (_03155_, _43578_, _43576_);
  and (_43579_, _43566_, _43329_);
  not (_43580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_43581_, _43566_, _43580_);
  or (_03159_, _43581_, _43579_);
  and (_43582_, _43566_, _43333_);
  not (_43583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_43584_, _43566_, _43583_);
  or (_03163_, _43584_, _43582_);
  and (_43585_, _43566_, _43337_);
  not (_43586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_43587_, _43566_, _43586_);
  or (_03166_, _43587_, _43585_);
  and (_43588_, _43566_, _43213_);
  not (_43589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_43590_, _43566_, _43589_);
  or (_03169_, _43590_, _43588_);
  and (_43591_, _43224_, _43209_);
  and (_43592_, _43591_, _43311_);
  not (_43593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_43594_, _43591_, _43593_);
  or (_03173_, _43594_, _43592_);
  and (_43595_, _43591_, _43317_);
  not (_43596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_43597_, _43591_, _43596_);
  or (_03177_, _43597_, _43595_);
  and (_43598_, _43591_, _43321_);
  not (_43599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_43600_, _43591_, _43599_);
  or (_03180_, _43600_, _43598_);
  and (_43601_, _43591_, _43325_);
  not (_43602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_43603_, _43591_, _43602_);
  or (_03183_, _43603_, _43601_);
  and (_43604_, _43591_, _43329_);
  not (_43605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_43606_, _43591_, _43605_);
  or (_03186_, _43606_, _43604_);
  and (_43607_, _43591_, _43333_);
  not (_43608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_43609_, _43591_, _43608_);
  or (_03190_, _43609_, _43607_);
  and (_43610_, _43591_, _43337_);
  not (_43611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_43612_, _43591_, _43611_);
  or (_03193_, _43612_, _43610_);
  and (_43613_, _43591_, _43213_);
  nor (_43614_, _43591_, _43166_);
  or (_03195_, _43614_, _43613_);
  and (_43615_, _43312_, _43209_);
  and (_43616_, _43615_, _43311_);
  not (_43617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_43618_, _43615_, _43617_);
  or (_03200_, _43618_, _43616_);
  and (_43619_, _43615_, _43317_);
  not (_43620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_43621_, _43615_, _43620_);
  or (_03203_, _43621_, _43619_);
  and (_43622_, _43615_, _43321_);
  not (_43623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_43624_, _43615_, _43623_);
  or (_03207_, _43624_, _43622_);
  and (_43625_, _43615_, _43325_);
  not (_43626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_43627_, _43615_, _43626_);
  or (_03211_, _43627_, _43625_);
  and (_43628_, _43615_, _43329_);
  not (_43629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_43630_, _43615_, _43629_);
  or (_03214_, _43630_, _43628_);
  and (_43631_, _43615_, _43333_);
  not (_43632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_43633_, _43615_, _43632_);
  or (_03218_, _43633_, _43631_);
  and (_43634_, _43615_, _43337_);
  not (_43635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_43636_, _43615_, _43635_);
  or (_03221_, _43636_, _43634_);
  and (_43637_, _43615_, _43213_);
  not (_43638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_43639_, _43615_, _43638_);
  or (_03224_, _43639_, _43637_);
  and (_43640_, _43343_, _43209_);
  and (_43641_, _43640_, _43311_);
  not (_43642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_43643_, _43640_, _43642_);
  or (_03228_, _43643_, _43641_);
  and (_43644_, _43640_, _43317_);
  not (_43645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_43646_, _43640_, _43645_);
  or (_03232_, _43646_, _43644_);
  and (_43647_, _43640_, _43321_);
  not (_43648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_43649_, _43640_, _43648_);
  or (_03236_, _43649_, _43647_);
  and (_43650_, _43640_, _43325_);
  not (_43651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_43652_, _43640_, _43651_);
  or (_03239_, _43652_, _43650_);
  and (_43653_, _43640_, _43329_);
  not (_43654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_43655_, _43640_, _43654_);
  or (_03243_, _43655_, _43653_);
  and (_43656_, _43640_, _43333_);
  not (_43657_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_43658_, _43640_, _43657_);
  or (_03246_, _43658_, _43656_);
  and (_43659_, _43640_, _43337_);
  not (_43660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_43661_, _43640_, _43660_);
  or (_03250_, _43661_, _43659_);
  and (_43662_, _43640_, _43213_);
  nor (_43663_, _43640_, _43176_);
  or (_03253_, _43663_, _43662_);
  and (_43664_, _43311_, _43211_);
  not (_43665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_43666_, _43211_, _43665_);
  or (_03257_, _43666_, _43664_);
  and (_43667_, _43317_, _43211_);
  not (_43668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_43669_, _43211_, _43668_);
  or (_03260_, _43669_, _43667_);
  and (_43670_, _43321_, _43211_);
  not (_43671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_43672_, _43211_, _43671_);
  or (_03263_, _43672_, _43670_);
  and (_43673_, _43325_, _43211_);
  not (_43674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_43675_, _43211_, _43674_);
  or (_03267_, _43675_, _43673_);
  and (_43676_, _43329_, _43211_);
  not (_43677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_43678_, _43211_, _43677_);
  or (_03270_, _43678_, _43676_);
  and (_43679_, _43333_, _43211_);
  not (_43680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_43681_, _43211_, _43680_);
  or (_03273_, _43681_, _43679_);
  and (_43682_, _43337_, _43211_);
  not (_43683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_43684_, _43211_, _43683_);
  or (_03276_, _43684_, _43682_);
  nor (_43685_, _42938_, _43371_);
  and (_43686_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_43687_, _43686_, _42837_);
  or (_43688_, _43687_, _43685_);
  and (_43689_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_43690_, _42938_, _43315_);
  nand (_43691_, _43690_, _42837_);
  or (_43692_, _43691_, _43689_);
  and (_43693_, _43692_, _43688_);
  or (_43694_, _43693_, _43122_);
  nor (_43695_, _42938_, _43470_);
  and (_43696_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_43697_, _43696_, _42837_);
  or (_43698_, _43697_, _43695_);
  and (_43699_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_43700_, _42938_, _43421_);
  nand (_43701_, _43700_, _42837_);
  or (_43702_, _43701_, _43699_);
  and (_43703_, _43702_, _43698_);
  or (_43704_, _43703_, _43086_);
  and (_43705_, _43704_, _43135_);
  and (_43706_, _43705_, _43694_);
  nand (_43707_, _42938_, _43495_);
  or (_43708_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_43709_, _43708_, _43707_);
  or (_43710_, _43709_, _43150_);
  or (_43711_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_43712_, _42938_, _43544_);
  and (_43713_, _43712_, _43711_);
  or (_43714_, _43713_, _42837_);
  and (_43715_, _43714_, _43710_);
  or (_43716_, _43715_, _43122_);
  nand (_43717_, _42938_, _43593_);
  or (_43718_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_43719_, _43718_, _43717_);
  or (_43720_, _43719_, _43150_);
  or (_43721_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_43722_, _42938_, _43642_);
  and (_43723_, _43722_, _43721_);
  or (_43724_, _43723_, _42837_);
  and (_43725_, _43724_, _43720_);
  or (_43726_, _43725_, _43086_);
  and (_43727_, _43726_, _42992_);
  and (_43728_, _43727_, _43716_);
  or (_43729_, _43728_, _43706_);
  or (_43730_, _43729_, _43121_);
  or (_43731_, _43186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_43732_, _43731_, _43190_);
  and (_43733_, _43732_, _43730_);
  and (_40469_, _43237_, _43223_);
  and (_43734_, _40469_, _43189_);
  or (_05039_, _43734_, _43733_);
  nor (_43735_, _42938_, _43374_);
  and (_43736_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_43737_, _43736_, _42837_);
  or (_43738_, _43737_, _43735_);
  and (_43739_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_43740_, _42938_, _43319_);
  nand (_43741_, _43740_, _42837_);
  or (_43742_, _43741_, _43739_);
  and (_43743_, _43742_, _43738_);
  or (_43744_, _43743_, _43122_);
  nor (_43745_, _42938_, _43473_);
  and (_43746_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_43747_, _43746_, _42837_);
  or (_43748_, _43747_, _43745_);
  and (_43749_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_43750_, _42938_, _43424_);
  nand (_43751_, _43750_, _42837_);
  or (_43752_, _43751_, _43749_);
  and (_43753_, _43752_, _43748_);
  or (_43754_, _43753_, _43086_);
  and (_43755_, _43754_, _43135_);
  and (_43756_, _43755_, _43744_);
  nand (_43757_, _42938_, _43498_);
  or (_43758_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_43759_, _43758_, _43757_);
  or (_43760_, _43759_, _43150_);
  or (_43766_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand (_43770_, _42938_, _43547_);
  and (_43777_, _43770_, _43766_);
  or (_43785_, _43777_, _42837_);
  and (_43789_, _43785_, _43760_);
  or (_43794_, _43789_, _43122_);
  nand (_43802_, _42938_, _43596_);
  or (_43808_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_43812_, _43808_, _43802_);
  or (_43819_, _43812_, _43150_);
  or (_43827_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand (_43831_, _42938_, _43645_);
  and (_43836_, _43831_, _43827_);
  or (_43844_, _43836_, _42837_);
  and (_43850_, _43844_, _43819_);
  or (_43853_, _43850_, _43086_);
  and (_43857_, _43853_, _42992_);
  and (_43868_, _43857_, _43794_);
  or (_43872_, _43868_, _43756_);
  or (_43879_, _43872_, _43121_);
  or (_43887_, _43186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_43891_, _43887_, _43190_);
  and (_43896_, _43891_, _43879_);
  and (_40470_, _43250_, _43223_);
  and (_43909_, _40470_, _43189_);
  or (_05041_, _43909_, _43896_);
  nor (_43919_, _42938_, _43377_);
  and (_43927_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_43931_, _43927_, _42837_);
  or (_43936_, _43931_, _43919_);
  and (_43944_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_43950_, _42938_, _43323_);
  nand (_43953_, _43950_, _42837_);
  or (_43954_, _43953_, _43944_);
  and (_43955_, _43954_, _43936_);
  or (_43956_, _43955_, _43122_);
  nor (_43957_, _42938_, _43476_);
  and (_43958_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_43959_, _43958_, _42837_);
  or (_43960_, _43959_, _43957_);
  and (_43961_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_43962_, _42938_, _43427_);
  nand (_43963_, _43962_, _42837_);
  or (_43964_, _43963_, _43961_);
  and (_43965_, _43964_, _43960_);
  or (_43966_, _43965_, _43086_);
  and (_43967_, _43966_, _43135_);
  and (_43968_, _43967_, _43956_);
  nand (_43969_, _42938_, _43501_);
  or (_43970_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_43971_, _43970_, _43969_);
  or (_43972_, _43971_, _43150_);
  or (_43973_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_43974_, _42938_, _43550_);
  and (_43975_, _43974_, _43973_);
  or (_43976_, _43975_, _42837_);
  and (_43977_, _43976_, _43972_);
  or (_43978_, _43977_, _43122_);
  nand (_43979_, _42938_, _43599_);
  or (_43980_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_43981_, _43980_, _43979_);
  or (_43982_, _43981_, _43150_);
  or (_43983_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_43984_, _42938_, _43648_);
  and (_43985_, _43984_, _43983_);
  or (_43986_, _43985_, _42837_);
  and (_43987_, _43986_, _43982_);
  or (_43988_, _43987_, _43086_);
  and (_43989_, _43988_, _42992_);
  and (_43990_, _43989_, _43978_);
  or (_43991_, _43990_, _43968_);
  or (_43992_, _43991_, _43121_);
  or (_43993_, _43186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_43994_, _43993_, _43190_);
  and (_43995_, _43994_, _43992_);
  and (_40471_, _43263_, _43223_);
  and (_43996_, _40471_, _43189_);
  or (_05043_, _43996_, _43995_);
  nor (_43997_, _42938_, _43380_);
  and (_43998_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_43999_, _43998_, _42837_);
  or (_44000_, _43999_, _43997_);
  and (_44001_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_44002_, _42938_, _43327_);
  nand (_44003_, _44002_, _42837_);
  or (_44004_, _44003_, _44001_);
  and (_44005_, _44004_, _44000_);
  or (_44006_, _44005_, _43122_);
  nor (_44007_, _42938_, _43479_);
  and (_44008_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_44009_, _44008_, _42837_);
  or (_44010_, _44009_, _44007_);
  and (_44011_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_44012_, _42938_, _43430_);
  nand (_44013_, _44012_, _42837_);
  or (_44014_, _44013_, _44011_);
  and (_44015_, _44014_, _44010_);
  or (_44016_, _44015_, _43086_);
  and (_44017_, _44016_, _43135_);
  and (_44018_, _44017_, _44006_);
  nand (_44019_, _42938_, _43504_);
  or (_44020_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_44021_, _44020_, _44019_);
  or (_44022_, _44021_, _43150_);
  or (_44023_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_44024_, _42938_, _43553_);
  and (_44025_, _44024_, _44023_);
  or (_44026_, _44025_, _42837_);
  and (_44027_, _44026_, _44022_);
  or (_44028_, _44027_, _43122_);
  nand (_44029_, _42938_, _43602_);
  or (_44030_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_44031_, _44030_, _44029_);
  or (_44032_, _44031_, _43150_);
  or (_44033_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_44034_, _42938_, _43651_);
  and (_44035_, _44034_, _44033_);
  or (_44036_, _44035_, _42837_);
  and (_44037_, _44036_, _44032_);
  or (_44038_, _44037_, _43086_);
  and (_44039_, _44038_, _42992_);
  and (_44040_, _44039_, _44028_);
  nor (_44041_, _44040_, _44018_);
  nor (_44042_, _44041_, _43121_);
  and (_44043_, _43121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_44044_, _44043_, _43189_);
  or (_44045_, _44044_, _44042_);
  and (_40472_, _43271_, _43223_);
  or (_44046_, _40472_, _43190_);
  and (_05045_, _44046_, _44045_);
  and (_44047_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_44048_, _42938_, _43331_);
  nand (_44049_, _44048_, _42837_);
  or (_44050_, _44049_, _44047_);
  nor (_44051_, _42938_, _43383_);
  and (_44052_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_44053_, _44052_, _42837_);
  or (_44054_, _44053_, _44051_);
  and (_44055_, _44054_, _44050_);
  or (_44056_, _44055_, _43122_);
  nor (_44057_, _42938_, _43482_);
  and (_44058_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_44059_, _44058_, _42837_);
  or (_44060_, _44059_, _44057_);
  and (_44061_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_44062_, _42938_, _43433_);
  nand (_44063_, _44062_, _42837_);
  or (_44064_, _44063_, _44061_);
  and (_44065_, _44064_, _44060_);
  or (_44066_, _44065_, _43086_);
  and (_44067_, _44066_, _43135_);
  and (_44068_, _44067_, _44056_);
  nor (_44069_, _42938_, _43580_);
  and (_44070_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_44071_, _44070_, _42837_);
  or (_44072_, _44071_, _44069_);
  and (_44073_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_44074_, _42938_, _43531_);
  nand (_44075_, _44074_, _42837_);
  or (_44076_, _44075_, _44073_);
  and (_44077_, _44076_, _44072_);
  or (_44078_, _44077_, _43122_);
  nor (_44079_, _42938_, _43677_);
  and (_44080_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_44081_, _44080_, _42837_);
  or (_44082_, _44081_, _44079_);
  and (_44083_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_44084_, _42938_, _43629_);
  nand (_44085_, _44084_, _42837_);
  or (_44086_, _44085_, _44083_);
  and (_44087_, _44086_, _44082_);
  or (_44088_, _44087_, _43086_);
  and (_44089_, _44088_, _42992_);
  and (_44090_, _44089_, _44078_);
  or (_44091_, _44090_, _44068_);
  and (_44092_, _44091_, _43188_);
  and (_44093_, _43282_, _43189_);
  and (_44094_, _43121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_44095_, _44094_, _44093_);
  or (_44096_, _44095_, _44092_);
  and (_05047_, _44096_, _43223_);
  nor (_44097_, _42938_, _43386_);
  and (_44098_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_44099_, _44098_, _42837_);
  or (_44100_, _44099_, _44097_);
  and (_44101_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_44102_, _42938_, _43335_);
  nand (_44103_, _44102_, _42837_);
  or (_44104_, _44103_, _44101_);
  and (_44105_, _44104_, _44100_);
  or (_44106_, _44105_, _43122_);
  nor (_44107_, _42938_, _43485_);
  and (_44108_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_44109_, _44108_, _42837_);
  or (_44110_, _44109_, _44107_);
  and (_44111_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_44112_, _42938_, _43436_);
  nand (_44113_, _44112_, _42837_);
  or (_44114_, _44113_, _44111_);
  and (_44115_, _44114_, _44110_);
  or (_44116_, _44115_, _43086_);
  and (_44117_, _44116_, _43135_);
  and (_44118_, _44117_, _44106_);
  nand (_44119_, _42938_, _43510_);
  or (_44120_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_44121_, _44120_, _44119_);
  or (_44122_, _44121_, _43150_);
  or (_44123_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_44124_, _42938_, _43559_);
  and (_44125_, _44124_, _44123_);
  or (_44126_, _44125_, _42837_);
  and (_44127_, _44126_, _44122_);
  or (_44128_, _44127_, _43122_);
  nand (_44129_, _42938_, _43608_);
  or (_44130_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_44131_, _44130_, _44129_);
  or (_44132_, _44131_, _43150_);
  or (_44133_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_44134_, _42938_, _43657_);
  and (_44135_, _44134_, _44133_);
  or (_44136_, _44135_, _42837_);
  and (_44137_, _44136_, _44132_);
  or (_44138_, _44137_, _43086_);
  and (_44139_, _44138_, _42992_);
  and (_44140_, _44139_, _44128_);
  or (_44141_, _44140_, _44118_);
  or (_44142_, _44141_, _43121_);
  or (_44143_, _43186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_44144_, _44143_, _43190_);
  and (_44145_, _44144_, _44142_);
  and (_40474_, _43295_, _43223_);
  and (_44146_, _40474_, _43189_);
  or (_05049_, _44146_, _44145_);
  or (_44147_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_44148_, _42938_, _43660_);
  and (_44149_, _44148_, _44147_);
  or (_44150_, _44149_, _42837_);
  nand (_00002_, _42938_, _43611_);
  or (_00003_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_00004_, _00003_, _00002_);
  or (_00005_, _00004_, _43150_);
  and (_00006_, _00005_, _42992_);
  and (_00007_, _00006_, _44150_);
  and (_00008_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_00009_, _42938_, _43439_);
  nand (_00010_, _00009_, _42837_);
  or (_00011_, _00010_, _00008_);
  nor (_00012_, _42938_, _43488_);
  and (_00013_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_00014_, _00013_, _42837_);
  or (_00015_, _00014_, _00012_);
  and (_00016_, _00015_, _43135_);
  and (_00017_, _00016_, _00011_);
  or (_00018_, _00017_, _00007_);
  and (_00019_, _00018_, _43122_);
  or (_00020_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_00021_, _42938_, _43562_);
  and (_00022_, _00021_, _00020_);
  or (_00023_, _00022_, _42837_);
  nand (_00024_, _42938_, _43513_);
  or (_00025_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_00026_, _00025_, _00024_);
  or (_00027_, _00026_, _43150_);
  and (_00028_, _00027_, _42992_);
  and (_00029_, _00028_, _00023_);
  and (_00030_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_00031_, _42938_, _43339_);
  nand (_00032_, _00031_, _42837_);
  or (_00033_, _00032_, _00030_);
  nor (_00034_, _42938_, _43389_);
  and (_00035_, _42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_00036_, _00035_, _42837_);
  or (_00037_, _00036_, _00034_);
  and (_00038_, _00037_, _43135_);
  and (_00039_, _00038_, _00033_);
  or (_00040_, _00039_, _00029_);
  and (_00041_, _00040_, _43086_);
  or (_00042_, _00041_, _43096_);
  or (_00043_, _00042_, _00019_);
  or (_00044_, _43186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_40475_, _43304_, _43223_);
  or (_00045_, _40475_, _43190_);
  and (_00046_, _00045_, _00044_);
  and (_05051_, _00046_, _00043_);
  or (_00047_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_00048_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_00049_, _00048_, \oc8051_gm_cxrom_1.cell0.data [7]);
  and (_00050_, _00049_, _00047_);
  or (_00051_, _00050_, rst);
  or (_00052_, \oc8051_gm_cxrom_1.cell0.data [7], _43223_);
  and (_05059_, _00052_, _00051_);
  or (_00053_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_00054_, \oc8051_gm_cxrom_1.cell0.data [0], _00048_);
  and (_00055_, _00054_, _00053_);
  or (_00056_, _00055_, rst);
  or (_00057_, \oc8051_gm_cxrom_1.cell0.data [0], _43223_);
  and (_05066_, _00057_, _00056_);
  or (_00058_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_00059_, \oc8051_gm_cxrom_1.cell0.data [1], _00048_);
  and (_00060_, _00059_, _00058_);
  or (_00061_, _00060_, rst);
  or (_00062_, \oc8051_gm_cxrom_1.cell0.data [1], _43223_);
  and (_05070_, _00062_, _00061_);
  or (_00063_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_00064_, \oc8051_gm_cxrom_1.cell0.data [2], _00048_);
  and (_00065_, _00064_, _00063_);
  or (_00066_, _00065_, rst);
  or (_00067_, \oc8051_gm_cxrom_1.cell0.data [2], _43223_);
  and (_05074_, _00067_, _00066_);
  or (_00068_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_00069_, \oc8051_gm_cxrom_1.cell0.data [3], _00048_);
  and (_00070_, _00069_, _00068_);
  or (_00071_, _00070_, rst);
  or (_00072_, \oc8051_gm_cxrom_1.cell0.data [3], _43223_);
  and (_05077_, _00072_, _00071_);
  or (_00073_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_00074_, \oc8051_gm_cxrom_1.cell0.data [4], _00048_);
  and (_00075_, _00074_, _00073_);
  or (_00076_, _00075_, rst);
  or (_00077_, \oc8051_gm_cxrom_1.cell0.data [4], _43223_);
  and (_05081_, _00077_, _00076_);
  or (_00078_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_00079_, \oc8051_gm_cxrom_1.cell0.data [5], _00048_);
  and (_00080_, _00079_, _00078_);
  or (_00081_, _00080_, rst);
  or (_00082_, \oc8051_gm_cxrom_1.cell0.data [5], _43223_);
  and (_05085_, _00082_, _00081_);
  or (_00083_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_00084_, \oc8051_gm_cxrom_1.cell0.data [6], _00048_);
  and (_00085_, _00084_, _00083_);
  or (_00086_, _00085_, rst);
  or (_00087_, \oc8051_gm_cxrom_1.cell0.data [6], _43223_);
  and (_05089_, _00087_, _00086_);
  or (_00088_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_00089_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_00090_, _00089_, \oc8051_gm_cxrom_1.cell1.data [7]);
  and (_00091_, _00090_, _00088_);
  or (_00092_, _00091_, rst);
  or (_00093_, \oc8051_gm_cxrom_1.cell1.data [7], _43223_);
  and (_05110_, _00093_, _00092_);
  or (_00094_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00095_, \oc8051_gm_cxrom_1.cell1.data [0], _00089_);
  and (_00096_, _00095_, _00094_);
  or (_00097_, _00096_, rst);
  or (_00098_, \oc8051_gm_cxrom_1.cell1.data [0], _43223_);
  and (_05117_, _00098_, _00097_);
  or (_00099_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00100_, \oc8051_gm_cxrom_1.cell1.data [1], _00089_);
  and (_00101_, _00100_, _00099_);
  or (_00102_, _00101_, rst);
  or (_00103_, \oc8051_gm_cxrom_1.cell1.data [1], _43223_);
  and (_05121_, _00103_, _00102_);
  or (_00104_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00105_, \oc8051_gm_cxrom_1.cell1.data [2], _00089_);
  and (_00106_, _00105_, _00104_);
  or (_00107_, _00106_, rst);
  or (_00108_, \oc8051_gm_cxrom_1.cell1.data [2], _43223_);
  and (_05125_, _00108_, _00107_);
  or (_00109_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00110_, \oc8051_gm_cxrom_1.cell1.data [3], _00089_);
  and (_00111_, _00110_, _00109_);
  or (_00112_, _00111_, rst);
  or (_00113_, \oc8051_gm_cxrom_1.cell1.data [3], _43223_);
  and (_05129_, _00113_, _00112_);
  or (_00114_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00115_, \oc8051_gm_cxrom_1.cell1.data [4], _00089_);
  and (_00116_, _00115_, _00114_);
  or (_00117_, _00116_, rst);
  or (_00118_, \oc8051_gm_cxrom_1.cell1.data [4], _43223_);
  and (_05133_, _00118_, _00117_);
  or (_00119_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00120_, \oc8051_gm_cxrom_1.cell1.data [5], _00089_);
  and (_00121_, _00120_, _00119_);
  or (_00122_, _00121_, rst);
  or (_00123_, \oc8051_gm_cxrom_1.cell1.data [5], _43223_);
  and (_05137_, _00123_, _00122_);
  or (_00124_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00125_, \oc8051_gm_cxrom_1.cell1.data [6], _00089_);
  and (_00126_, _00125_, _00124_);
  or (_00127_, _00126_, rst);
  or (_00128_, \oc8051_gm_cxrom_1.cell1.data [6], _43223_);
  and (_05141_, _00128_, _00127_);
  or (_00129_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_00130_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_00131_, _00130_, \oc8051_gm_cxrom_1.cell2.data [7]);
  and (_00132_, _00131_, _00129_);
  or (_00133_, _00132_, rst);
  or (_00134_, \oc8051_gm_cxrom_1.cell2.data [7], _43223_);
  and (_05162_, _00134_, _00133_);
  or (_00135_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00136_, \oc8051_gm_cxrom_1.cell2.data [0], _00130_);
  and (_00138_, _00136_, _00135_);
  or (_00140_, _00138_, rst);
  or (_00142_, \oc8051_gm_cxrom_1.cell2.data [0], _43223_);
  and (_05169_, _00142_, _00140_);
  or (_00145_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00147_, \oc8051_gm_cxrom_1.cell2.data [1], _00130_);
  and (_00149_, _00147_, _00145_);
  or (_00151_, _00149_, rst);
  or (_00153_, \oc8051_gm_cxrom_1.cell2.data [1], _43223_);
  and (_05173_, _00153_, _00151_);
  or (_00156_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00158_, \oc8051_gm_cxrom_1.cell2.data [2], _00130_);
  and (_00160_, _00158_, _00156_);
  or (_00162_, _00160_, rst);
  or (_00164_, \oc8051_gm_cxrom_1.cell2.data [2], _43223_);
  and (_05177_, _00164_, _00162_);
  or (_00167_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00169_, \oc8051_gm_cxrom_1.cell2.data [3], _00130_);
  and (_00171_, _00169_, _00167_);
  or (_00173_, _00171_, rst);
  or (_00175_, \oc8051_gm_cxrom_1.cell2.data [3], _43223_);
  and (_05181_, _00175_, _00173_);
  or (_00178_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00180_, \oc8051_gm_cxrom_1.cell2.data [4], _00130_);
  and (_00182_, _00180_, _00178_);
  or (_00184_, _00182_, rst);
  or (_00186_, \oc8051_gm_cxrom_1.cell2.data [4], _43223_);
  and (_05185_, _00186_, _00184_);
  or (_00189_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00191_, \oc8051_gm_cxrom_1.cell2.data [5], _00130_);
  and (_00193_, _00191_, _00189_);
  or (_00194_, _00193_, rst);
  or (_00195_, \oc8051_gm_cxrom_1.cell2.data [5], _43223_);
  and (_05188_, _00195_, _00194_);
  or (_00196_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00197_, \oc8051_gm_cxrom_1.cell2.data [6], _00130_);
  and (_00198_, _00197_, _00196_);
  or (_00199_, _00198_, rst);
  or (_00200_, \oc8051_gm_cxrom_1.cell2.data [6], _43223_);
  and (_05192_, _00200_, _00199_);
  or (_00201_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_00202_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_00203_, _00202_, \oc8051_gm_cxrom_1.cell3.data [7]);
  and (_00204_, _00203_, _00201_);
  or (_00205_, _00204_, rst);
  or (_00206_, \oc8051_gm_cxrom_1.cell3.data [7], _43223_);
  and (_05214_, _00206_, _00205_);
  or (_00207_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00208_, \oc8051_gm_cxrom_1.cell3.data [0], _00202_);
  and (_00209_, _00208_, _00207_);
  or (_00210_, _00209_, rst);
  or (_00211_, \oc8051_gm_cxrom_1.cell3.data [0], _43223_);
  and (_05220_, _00211_, _00210_);
  or (_00212_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00213_, \oc8051_gm_cxrom_1.cell3.data [1], _00202_);
  and (_00214_, _00213_, _00212_);
  or (_00215_, _00214_, rst);
  or (_00216_, \oc8051_gm_cxrom_1.cell3.data [1], _43223_);
  and (_05224_, _00216_, _00215_);
  or (_00217_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00218_, \oc8051_gm_cxrom_1.cell3.data [2], _00202_);
  and (_00219_, _00218_, _00217_);
  or (_00220_, _00219_, rst);
  or (_00221_, \oc8051_gm_cxrom_1.cell3.data [2], _43223_);
  and (_05228_, _00221_, _00220_);
  or (_00222_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00223_, \oc8051_gm_cxrom_1.cell3.data [3], _00202_);
  and (_00224_, _00223_, _00222_);
  or (_00225_, _00224_, rst);
  or (_00226_, \oc8051_gm_cxrom_1.cell3.data [3], _43223_);
  and (_05232_, _00226_, _00225_);
  or (_00227_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00228_, \oc8051_gm_cxrom_1.cell3.data [4], _00202_);
  and (_00229_, _00228_, _00227_);
  or (_00230_, _00229_, rst);
  or (_00231_, \oc8051_gm_cxrom_1.cell3.data [4], _43223_);
  and (_05236_, _00231_, _00230_);
  or (_00232_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00233_, \oc8051_gm_cxrom_1.cell3.data [5], _00202_);
  and (_00234_, _00233_, _00232_);
  or (_00235_, _00234_, rst);
  or (_00236_, \oc8051_gm_cxrom_1.cell3.data [5], _43223_);
  and (_05240_, _00236_, _00235_);
  or (_00237_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00238_, \oc8051_gm_cxrom_1.cell3.data [6], _00202_);
  and (_00239_, _00238_, _00237_);
  or (_00240_, _00239_, rst);
  or (_00241_, \oc8051_gm_cxrom_1.cell3.data [6], _43223_);
  and (_05244_, _00241_, _00240_);
  or (_00242_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_00243_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_00244_, _00243_, \oc8051_gm_cxrom_1.cell4.data [7]);
  and (_00245_, _00244_, _00242_);
  or (_00246_, _00245_, rst);
  or (_00247_, \oc8051_gm_cxrom_1.cell4.data [7], _43223_);
  and (_05265_, _00247_, _00246_);
  or (_00248_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00249_, \oc8051_gm_cxrom_1.cell4.data [0], _00243_);
  and (_00250_, _00249_, _00248_);
  or (_00251_, _00250_, rst);
  or (_00252_, \oc8051_gm_cxrom_1.cell4.data [0], _43223_);
  and (_05272_, _00252_, _00251_);
  or (_00253_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00254_, \oc8051_gm_cxrom_1.cell4.data [1], _00243_);
  and (_00255_, _00254_, _00253_);
  or (_00256_, _00255_, rst);
  or (_00257_, \oc8051_gm_cxrom_1.cell4.data [1], _43223_);
  and (_05276_, _00257_, _00256_);
  or (_00258_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00259_, \oc8051_gm_cxrom_1.cell4.data [2], _00243_);
  and (_00260_, _00259_, _00258_);
  or (_00261_, _00260_, rst);
  or (_00262_, \oc8051_gm_cxrom_1.cell4.data [2], _43223_);
  and (_05280_, _00262_, _00261_);
  or (_00263_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00264_, \oc8051_gm_cxrom_1.cell4.data [3], _00243_);
  and (_00265_, _00264_, _00263_);
  or (_00266_, _00265_, rst);
  or (_00267_, \oc8051_gm_cxrom_1.cell4.data [3], _43223_);
  and (_05284_, _00267_, _00266_);
  or (_00268_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00269_, \oc8051_gm_cxrom_1.cell4.data [4], _00243_);
  and (_00270_, _00269_, _00268_);
  or (_00271_, _00270_, rst);
  or (_00272_, \oc8051_gm_cxrom_1.cell4.data [4], _43223_);
  and (_05288_, _00272_, _00271_);
  or (_00273_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00274_, \oc8051_gm_cxrom_1.cell4.data [5], _00243_);
  and (_00275_, _00274_, _00273_);
  or (_00276_, _00275_, rst);
  or (_00277_, \oc8051_gm_cxrom_1.cell4.data [5], _43223_);
  and (_05292_, _00277_, _00276_);
  or (_00278_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00279_, \oc8051_gm_cxrom_1.cell4.data [6], _00243_);
  and (_00280_, _00279_, _00278_);
  or (_00281_, _00280_, rst);
  or (_00282_, \oc8051_gm_cxrom_1.cell4.data [6], _43223_);
  and (_05295_, _00282_, _00281_);
  or (_00283_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_00284_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_00285_, _00284_, \oc8051_gm_cxrom_1.cell5.data [7]);
  and (_00286_, _00285_, _00283_);
  or (_00287_, _00286_, rst);
  or (_00288_, \oc8051_gm_cxrom_1.cell5.data [7], _43223_);
  and (_05317_, _00288_, _00287_);
  or (_00289_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00290_, \oc8051_gm_cxrom_1.cell5.data [0], _00284_);
  and (_00291_, _00290_, _00289_);
  or (_00292_, _00291_, rst);
  or (_00293_, \oc8051_gm_cxrom_1.cell5.data [0], _43223_);
  and (_05324_, _00293_, _00292_);
  or (_00294_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00295_, \oc8051_gm_cxrom_1.cell5.data [1], _00284_);
  and (_00296_, _00295_, _00294_);
  or (_00297_, _00296_, rst);
  or (_00298_, \oc8051_gm_cxrom_1.cell5.data [1], _43223_);
  and (_05328_, _00298_, _00297_);
  or (_00299_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00300_, \oc8051_gm_cxrom_1.cell5.data [2], _00284_);
  and (_00301_, _00300_, _00299_);
  or (_00302_, _00301_, rst);
  or (_00303_, \oc8051_gm_cxrom_1.cell5.data [2], _43223_);
  and (_05331_, _00303_, _00302_);
  or (_00304_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00305_, \oc8051_gm_cxrom_1.cell5.data [3], _00284_);
  and (_00306_, _00305_, _00304_);
  or (_00307_, _00306_, rst);
  or (_00308_, \oc8051_gm_cxrom_1.cell5.data [3], _43223_);
  and (_05335_, _00308_, _00307_);
  or (_00309_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00310_, \oc8051_gm_cxrom_1.cell5.data [4], _00284_);
  and (_00311_, _00310_, _00309_);
  or (_00312_, _00311_, rst);
  or (_00313_, \oc8051_gm_cxrom_1.cell5.data [4], _43223_);
  and (_05339_, _00313_, _00312_);
  or (_00314_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00315_, \oc8051_gm_cxrom_1.cell5.data [5], _00284_);
  and (_00316_, _00315_, _00314_);
  or (_00317_, _00316_, rst);
  or (_00318_, \oc8051_gm_cxrom_1.cell5.data [5], _43223_);
  and (_05343_, _00318_, _00317_);
  or (_00319_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00320_, \oc8051_gm_cxrom_1.cell5.data [6], _00284_);
  and (_00321_, _00320_, _00319_);
  or (_00322_, _00321_, rst);
  or (_00323_, \oc8051_gm_cxrom_1.cell5.data [6], _43223_);
  and (_05347_, _00323_, _00322_);
  or (_00324_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_00325_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_00326_, _00325_, \oc8051_gm_cxrom_1.cell6.data [7]);
  and (_00327_, _00326_, _00324_);
  or (_00328_, _00327_, rst);
  or (_00329_, \oc8051_gm_cxrom_1.cell6.data [7], _43223_);
  and (_05368_, _00329_, _00328_);
  or (_00330_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00331_, \oc8051_gm_cxrom_1.cell6.data [0], _00325_);
  and (_00332_, _00331_, _00330_);
  or (_00333_, _00332_, rst);
  or (_00334_, \oc8051_gm_cxrom_1.cell6.data [0], _43223_);
  and (_05375_, _00334_, _00333_);
  or (_00335_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00336_, \oc8051_gm_cxrom_1.cell6.data [1], _00325_);
  and (_00337_, _00336_, _00335_);
  or (_00338_, _00337_, rst);
  or (_00339_, \oc8051_gm_cxrom_1.cell6.data [1], _43223_);
  and (_05379_, _00339_, _00338_);
  or (_00340_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00341_, \oc8051_gm_cxrom_1.cell6.data [2], _00325_);
  and (_00342_, _00341_, _00340_);
  or (_00343_, _00342_, rst);
  or (_00344_, \oc8051_gm_cxrom_1.cell6.data [2], _43223_);
  and (_05383_, _00344_, _00343_);
  or (_00345_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00346_, \oc8051_gm_cxrom_1.cell6.data [3], _00325_);
  and (_00347_, _00346_, _00345_);
  or (_00348_, _00347_, rst);
  or (_00349_, \oc8051_gm_cxrom_1.cell6.data [3], _43223_);
  and (_05387_, _00349_, _00348_);
  or (_00350_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00351_, \oc8051_gm_cxrom_1.cell6.data [4], _00325_);
  and (_00352_, _00351_, _00350_);
  or (_00353_, _00352_, rst);
  or (_00354_, \oc8051_gm_cxrom_1.cell6.data [4], _43223_);
  and (_05391_, _00354_, _00353_);
  or (_00355_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00356_, \oc8051_gm_cxrom_1.cell6.data [5], _00325_);
  and (_00357_, _00356_, _00355_);
  or (_00358_, _00357_, rst);
  or (_00359_, \oc8051_gm_cxrom_1.cell6.data [5], _43223_);
  and (_05395_, _00359_, _00358_);
  or (_00360_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00361_, \oc8051_gm_cxrom_1.cell6.data [6], _00325_);
  and (_00362_, _00361_, _00360_);
  or (_00363_, _00362_, rst);
  or (_00364_, \oc8051_gm_cxrom_1.cell6.data [6], _43223_);
  and (_05399_, _00364_, _00363_);
  or (_00365_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_00366_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_00367_, _00366_, \oc8051_gm_cxrom_1.cell7.data [7]);
  and (_00368_, _00367_, _00365_);
  or (_00369_, _00368_, rst);
  or (_00370_, \oc8051_gm_cxrom_1.cell7.data [7], _43223_);
  and (_05420_, _00370_, _00369_);
  or (_00371_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00372_, \oc8051_gm_cxrom_1.cell7.data [0], _00366_);
  and (_00373_, _00372_, _00371_);
  or (_00374_, _00373_, rst);
  or (_00375_, \oc8051_gm_cxrom_1.cell7.data [0], _43223_);
  and (_05427_, _00375_, _00374_);
  or (_00376_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00377_, \oc8051_gm_cxrom_1.cell7.data [1], _00366_);
  and (_00378_, _00377_, _00376_);
  or (_00379_, _00378_, rst);
  or (_00380_, \oc8051_gm_cxrom_1.cell7.data [1], _43223_);
  and (_05431_, _00380_, _00379_);
  or (_00381_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00382_, \oc8051_gm_cxrom_1.cell7.data [2], _00366_);
  and (_00383_, _00382_, _00381_);
  or (_00384_, _00383_, rst);
  or (_00385_, \oc8051_gm_cxrom_1.cell7.data [2], _43223_);
  and (_05435_, _00385_, _00384_);
  or (_00386_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00387_, \oc8051_gm_cxrom_1.cell7.data [3], _00366_);
  and (_00388_, _00387_, _00386_);
  or (_00389_, _00388_, rst);
  or (_00390_, \oc8051_gm_cxrom_1.cell7.data [3], _43223_);
  and (_05439_, _00390_, _00389_);
  or (_00391_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00392_, \oc8051_gm_cxrom_1.cell7.data [4], _00366_);
  and (_00393_, _00392_, _00391_);
  or (_00394_, _00393_, rst);
  or (_00395_, \oc8051_gm_cxrom_1.cell7.data [4], _43223_);
  and (_05442_, _00395_, _00394_);
  or (_00396_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00397_, \oc8051_gm_cxrom_1.cell7.data [5], _00366_);
  and (_00398_, _00397_, _00396_);
  or (_00399_, _00398_, rst);
  or (_00400_, \oc8051_gm_cxrom_1.cell7.data [5], _43223_);
  and (_05446_, _00400_, _00399_);
  or (_00401_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00402_, \oc8051_gm_cxrom_1.cell7.data [6], _00366_);
  and (_00403_, _00402_, _00401_);
  or (_00404_, _00403_, rst);
  or (_00405_, \oc8051_gm_cxrom_1.cell7.data [6], _43223_);
  and (_05450_, _00405_, _00404_);
  or (_00406_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_00407_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_00408_, _00407_, \oc8051_gm_cxrom_1.cell8.data [7]);
  and (_00409_, _00408_, _00406_);
  or (_00410_, _00409_, rst);
  or (_00411_, \oc8051_gm_cxrom_1.cell8.data [7], _43223_);
  and (_05472_, _00411_, _00410_);
  or (_00412_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00413_, \oc8051_gm_cxrom_1.cell8.data [0], _00407_);
  and (_00414_, _00413_, _00412_);
  or (_00415_, _00414_, rst);
  or (_00416_, \oc8051_gm_cxrom_1.cell8.data [0], _43223_);
  and (_05478_, _00416_, _00415_);
  or (_00417_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00418_, \oc8051_gm_cxrom_1.cell8.data [1], _00407_);
  and (_00419_, _00418_, _00417_);
  or (_00420_, _00419_, rst);
  or (_00421_, \oc8051_gm_cxrom_1.cell8.data [1], _43223_);
  and (_05482_, _00421_, _00420_);
  or (_00422_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00423_, \oc8051_gm_cxrom_1.cell8.data [2], _00407_);
  and (_00424_, _00423_, _00422_);
  or (_00425_, _00424_, rst);
  or (_00426_, \oc8051_gm_cxrom_1.cell8.data [2], _43223_);
  and (_05486_, _00426_, _00425_);
  or (_00427_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00428_, \oc8051_gm_cxrom_1.cell8.data [3], _00407_);
  and (_00429_, _00428_, _00427_);
  or (_00430_, _00429_, rst);
  or (_00431_, \oc8051_gm_cxrom_1.cell8.data [3], _43223_);
  and (_05490_, _00431_, _00430_);
  or (_00432_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00433_, \oc8051_gm_cxrom_1.cell8.data [4], _00407_);
  and (_00434_, _00433_, _00432_);
  or (_00435_, _00434_, rst);
  or (_00436_, \oc8051_gm_cxrom_1.cell8.data [4], _43223_);
  and (_05494_, _00436_, _00435_);
  or (_00437_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00438_, \oc8051_gm_cxrom_1.cell8.data [5], _00407_);
  and (_00439_, _00438_, _00437_);
  or (_00440_, _00439_, rst);
  or (_00441_, \oc8051_gm_cxrom_1.cell8.data [5], _43223_);
  and (_05498_, _00441_, _00440_);
  or (_00442_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00443_, \oc8051_gm_cxrom_1.cell8.data [6], _00407_);
  and (_00444_, _00443_, _00442_);
  or (_00445_, _00444_, rst);
  or (_00446_, \oc8051_gm_cxrom_1.cell8.data [6], _43223_);
  and (_05502_, _00446_, _00445_);
  or (_00447_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_00448_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_00449_, _00448_, \oc8051_gm_cxrom_1.cell9.data [7]);
  and (_00450_, _00449_, _00447_);
  or (_00451_, _00450_, rst);
  or (_00452_, \oc8051_gm_cxrom_1.cell9.data [7], _43223_);
  and (_05523_, _00452_, _00451_);
  or (_00453_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00454_, \oc8051_gm_cxrom_1.cell9.data [0], _00448_);
  and (_00455_, _00454_, _00453_);
  or (_00456_, _00455_, rst);
  or (_00457_, \oc8051_gm_cxrom_1.cell9.data [0], _43223_);
  and (_05530_, _00457_, _00456_);
  or (_00458_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00459_, \oc8051_gm_cxrom_1.cell9.data [1], _00448_);
  and (_00460_, _00459_, _00458_);
  or (_00461_, _00460_, rst);
  or (_00462_, \oc8051_gm_cxrom_1.cell9.data [1], _43223_);
  and (_05534_, _00462_, _00461_);
  or (_00463_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00464_, \oc8051_gm_cxrom_1.cell9.data [2], _00448_);
  and (_00465_, _00464_, _00463_);
  or (_00466_, _00465_, rst);
  or (_00467_, \oc8051_gm_cxrom_1.cell9.data [2], _43223_);
  and (_05538_, _00467_, _00466_);
  or (_00468_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00469_, \oc8051_gm_cxrom_1.cell9.data [3], _00448_);
  and (_00470_, _00469_, _00468_);
  or (_00471_, _00470_, rst);
  or (_00472_, \oc8051_gm_cxrom_1.cell9.data [3], _43223_);
  and (_05542_, _00472_, _00471_);
  or (_00473_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00474_, \oc8051_gm_cxrom_1.cell9.data [4], _00448_);
  and (_00475_, _00474_, _00473_);
  or (_00476_, _00475_, rst);
  or (_00477_, \oc8051_gm_cxrom_1.cell9.data [4], _43223_);
  and (_05546_, _00477_, _00476_);
  or (_00478_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00479_, \oc8051_gm_cxrom_1.cell9.data [5], _00448_);
  and (_00480_, _00479_, _00478_);
  or (_00481_, _00480_, rst);
  or (_00482_, \oc8051_gm_cxrom_1.cell9.data [5], _43223_);
  and (_05549_, _00482_, _00481_);
  or (_00483_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00484_, \oc8051_gm_cxrom_1.cell9.data [6], _00448_);
  and (_00485_, _00484_, _00483_);
  or (_00486_, _00485_, rst);
  or (_00487_, \oc8051_gm_cxrom_1.cell9.data [6], _43223_);
  and (_05553_, _00487_, _00486_);
  or (_00488_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_00489_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_00490_, _00489_, \oc8051_gm_cxrom_1.cell10.data [7]);
  and (_00491_, _00490_, _00488_);
  or (_00492_, _00491_, rst);
  or (_00493_, \oc8051_gm_cxrom_1.cell10.data [7], _43223_);
  and (_05575_, _00493_, _00492_);
  or (_00494_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00495_, \oc8051_gm_cxrom_1.cell10.data [0], _00489_);
  and (_00496_, _00495_, _00494_);
  or (_00497_, _00496_, rst);
  or (_00498_, \oc8051_gm_cxrom_1.cell10.data [0], _43223_);
  and (_05582_, _00498_, _00497_);
  or (_00499_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00500_, \oc8051_gm_cxrom_1.cell10.data [1], _00489_);
  and (_00501_, _00500_, _00499_);
  or (_00502_, _00501_, rst);
  or (_00503_, \oc8051_gm_cxrom_1.cell10.data [1], _43223_);
  and (_05586_, _00503_, _00502_);
  or (_00504_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00505_, \oc8051_gm_cxrom_1.cell10.data [2], _00489_);
  and (_00506_, _00505_, _00504_);
  or (_00507_, _00506_, rst);
  or (_00508_, \oc8051_gm_cxrom_1.cell10.data [2], _43223_);
  and (_05590_, _00508_, _00507_);
  or (_00509_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00510_, \oc8051_gm_cxrom_1.cell10.data [3], _00489_);
  and (_00511_, _00510_, _00509_);
  or (_00512_, _00511_, rst);
  or (_00513_, \oc8051_gm_cxrom_1.cell10.data [3], _43223_);
  and (_05594_, _00513_, _00512_);
  or (_00514_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00515_, \oc8051_gm_cxrom_1.cell10.data [4], _00489_);
  and (_00516_, _00515_, _00514_);
  or (_00517_, _00516_, rst);
  or (_00518_, \oc8051_gm_cxrom_1.cell10.data [4], _43223_);
  and (_05598_, _00518_, _00517_);
  or (_00519_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00520_, \oc8051_gm_cxrom_1.cell10.data [5], _00489_);
  and (_00521_, _00520_, _00519_);
  or (_00522_, _00521_, rst);
  or (_00523_, \oc8051_gm_cxrom_1.cell10.data [5], _43223_);
  and (_05602_, _00523_, _00522_);
  or (_00524_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00525_, \oc8051_gm_cxrom_1.cell10.data [6], _00489_);
  and (_00526_, _00525_, _00524_);
  or (_00527_, _00526_, rst);
  or (_00528_, \oc8051_gm_cxrom_1.cell10.data [6], _43223_);
  and (_05606_, _00528_, _00527_);
  or (_00529_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_00530_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_00531_, _00530_, \oc8051_gm_cxrom_1.cell11.data [7]);
  and (_00532_, _00531_, _00529_);
  or (_00533_, _00532_, rst);
  or (_00534_, \oc8051_gm_cxrom_1.cell11.data [7], _43223_);
  and (_05628_, _00534_, _00533_);
  or (_00535_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00536_, \oc8051_gm_cxrom_1.cell11.data [0], _00530_);
  and (_00537_, _00536_, _00535_);
  or (_00538_, _00537_, rst);
  or (_00539_, \oc8051_gm_cxrom_1.cell11.data [0], _43223_);
  and (_05635_, _00539_, _00538_);
  or (_00540_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00541_, \oc8051_gm_cxrom_1.cell11.data [1], _00530_);
  and (_00542_, _00541_, _00540_);
  or (_00543_, _00542_, rst);
  or (_00544_, \oc8051_gm_cxrom_1.cell11.data [1], _43223_);
  and (_05639_, _00544_, _00543_);
  or (_00545_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00546_, \oc8051_gm_cxrom_1.cell11.data [2], _00530_);
  and (_00547_, _00546_, _00545_);
  or (_00548_, _00547_, rst);
  or (_00549_, \oc8051_gm_cxrom_1.cell11.data [2], _43223_);
  and (_05643_, _00549_, _00548_);
  or (_00551_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00553_, \oc8051_gm_cxrom_1.cell11.data [3], _00530_);
  and (_00554_, _00553_, _00551_);
  or (_00556_, _00554_, rst);
  or (_00557_, \oc8051_gm_cxrom_1.cell11.data [3], _43223_);
  and (_05647_, _00557_, _00556_);
  or (_00559_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00561_, \oc8051_gm_cxrom_1.cell11.data [4], _00530_);
  and (_00562_, _00561_, _00559_);
  or (_00564_, _00562_, rst);
  or (_00565_, \oc8051_gm_cxrom_1.cell11.data [4], _43223_);
  and (_05651_, _00565_, _00564_);
  or (_00567_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00569_, \oc8051_gm_cxrom_1.cell11.data [5], _00530_);
  and (_00570_, _00569_, _00567_);
  or (_00572_, _00570_, rst);
  or (_00573_, \oc8051_gm_cxrom_1.cell11.data [5], _43223_);
  and (_05655_, _00573_, _00572_);
  or (_00575_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00577_, \oc8051_gm_cxrom_1.cell11.data [6], _00530_);
  and (_00578_, _00577_, _00575_);
  or (_00580_, _00578_, rst);
  or (_00581_, \oc8051_gm_cxrom_1.cell11.data [6], _43223_);
  and (_05659_, _00581_, _00580_);
  or (_00583_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_00585_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_00586_, _00585_, \oc8051_gm_cxrom_1.cell12.data [7]);
  and (_00588_, _00586_, _00583_);
  or (_00589_, _00588_, rst);
  or (_00591_, \oc8051_gm_cxrom_1.cell12.data [7], _43223_);
  and (_05681_, _00591_, _00589_);
  or (_00593_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00594_, \oc8051_gm_cxrom_1.cell12.data [0], _00585_);
  and (_00596_, _00594_, _00593_);
  or (_00597_, _00596_, rst);
  or (_00599_, \oc8051_gm_cxrom_1.cell12.data [0], _43223_);
  and (_05688_, _00599_, _00597_);
  or (_00600_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00601_, \oc8051_gm_cxrom_1.cell12.data [1], _00585_);
  and (_00602_, _00601_, _00600_);
  or (_00603_, _00602_, rst);
  or (_00604_, \oc8051_gm_cxrom_1.cell12.data [1], _43223_);
  and (_05692_, _00604_, _00603_);
  or (_00605_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00606_, \oc8051_gm_cxrom_1.cell12.data [2], _00585_);
  and (_00607_, _00606_, _00605_);
  or (_00608_, _00607_, rst);
  or (_00609_, \oc8051_gm_cxrom_1.cell12.data [2], _43223_);
  and (_05696_, _00609_, _00608_);
  or (_00610_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00611_, \oc8051_gm_cxrom_1.cell12.data [3], _00585_);
  and (_00612_, _00611_, _00610_);
  or (_00613_, _00612_, rst);
  or (_00614_, \oc8051_gm_cxrom_1.cell12.data [3], _43223_);
  and (_05700_, _00614_, _00613_);
  or (_00615_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00616_, \oc8051_gm_cxrom_1.cell12.data [4], _00585_);
  and (_00617_, _00616_, _00615_);
  or (_00618_, _00617_, rst);
  or (_00619_, \oc8051_gm_cxrom_1.cell12.data [4], _43223_);
  and (_05704_, _00619_, _00618_);
  or (_00620_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00621_, \oc8051_gm_cxrom_1.cell12.data [5], _00585_);
  and (_00622_, _00621_, _00620_);
  or (_00623_, _00622_, rst);
  or (_00624_, \oc8051_gm_cxrom_1.cell12.data [5], _43223_);
  and (_05708_, _00624_, _00623_);
  or (_00625_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00626_, \oc8051_gm_cxrom_1.cell12.data [6], _00585_);
  and (_00627_, _00626_, _00625_);
  or (_00628_, _00627_, rst);
  or (_00629_, \oc8051_gm_cxrom_1.cell12.data [6], _43223_);
  and (_05712_, _00629_, _00628_);
  or (_00630_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_00631_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_00632_, _00631_, \oc8051_gm_cxrom_1.cell13.data [7]);
  and (_00633_, _00632_, _00630_);
  or (_00634_, _00633_, rst);
  or (_00635_, \oc8051_gm_cxrom_1.cell13.data [7], _43223_);
  and (_05734_, _00635_, _00634_);
  or (_00636_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00637_, \oc8051_gm_cxrom_1.cell13.data [0], _00631_);
  and (_00638_, _00637_, _00636_);
  or (_00639_, _00638_, rst);
  or (_00640_, \oc8051_gm_cxrom_1.cell13.data [0], _43223_);
  and (_05741_, _00640_, _00639_);
  or (_00641_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00642_, \oc8051_gm_cxrom_1.cell13.data [1], _00631_);
  and (_00643_, _00642_, _00641_);
  or (_00644_, _00643_, rst);
  or (_00645_, \oc8051_gm_cxrom_1.cell13.data [1], _43223_);
  and (_05745_, _00645_, _00644_);
  or (_00646_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00647_, \oc8051_gm_cxrom_1.cell13.data [2], _00631_);
  and (_00648_, _00647_, _00646_);
  or (_00649_, _00648_, rst);
  or (_00650_, \oc8051_gm_cxrom_1.cell13.data [2], _43223_);
  and (_05749_, _00650_, _00649_);
  or (_00651_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00652_, \oc8051_gm_cxrom_1.cell13.data [3], _00631_);
  and (_00653_, _00652_, _00651_);
  or (_00654_, _00653_, rst);
  or (_00655_, \oc8051_gm_cxrom_1.cell13.data [3], _43223_);
  and (_05753_, _00655_, _00654_);
  or (_00656_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00657_, \oc8051_gm_cxrom_1.cell13.data [4], _00631_);
  and (_00658_, _00657_, _00656_);
  or (_00659_, _00658_, rst);
  or (_00660_, \oc8051_gm_cxrom_1.cell13.data [4], _43223_);
  and (_05757_, _00660_, _00659_);
  or (_00661_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00662_, \oc8051_gm_cxrom_1.cell13.data [5], _00631_);
  and (_00663_, _00662_, _00661_);
  or (_00664_, _00663_, rst);
  or (_00665_, \oc8051_gm_cxrom_1.cell13.data [5], _43223_);
  and (_05761_, _00665_, _00664_);
  or (_00666_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00667_, \oc8051_gm_cxrom_1.cell13.data [6], _00631_);
  and (_00668_, _00667_, _00666_);
  or (_00669_, _00668_, rst);
  or (_00670_, \oc8051_gm_cxrom_1.cell13.data [6], _43223_);
  and (_05765_, _00670_, _00669_);
  or (_00671_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_00672_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_00673_, _00672_, \oc8051_gm_cxrom_1.cell14.data [7]);
  and (_00674_, _00673_, _00671_);
  or (_00675_, _00674_, rst);
  or (_00676_, \oc8051_gm_cxrom_1.cell14.data [7], _43223_);
  and (_05787_, _00676_, _00675_);
  or (_00677_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00678_, \oc8051_gm_cxrom_1.cell14.data [0], _00672_);
  and (_00679_, _00678_, _00677_);
  or (_00680_, _00679_, rst);
  or (_00681_, \oc8051_gm_cxrom_1.cell14.data [0], _43223_);
  and (_05794_, _00681_, _00680_);
  or (_00682_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00683_, \oc8051_gm_cxrom_1.cell14.data [1], _00672_);
  and (_00684_, _00683_, _00682_);
  or (_00685_, _00684_, rst);
  or (_00686_, \oc8051_gm_cxrom_1.cell14.data [1], _43223_);
  and (_05798_, _00686_, _00685_);
  or (_00687_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00688_, \oc8051_gm_cxrom_1.cell14.data [2], _00672_);
  and (_00689_, _00688_, _00687_);
  or (_00690_, _00689_, rst);
  or (_00691_, \oc8051_gm_cxrom_1.cell14.data [2], _43223_);
  and (_05802_, _00691_, _00690_);
  or (_00692_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00693_, \oc8051_gm_cxrom_1.cell14.data [3], _00672_);
  and (_00694_, _00693_, _00692_);
  or (_00695_, _00694_, rst);
  or (_00696_, \oc8051_gm_cxrom_1.cell14.data [3], _43223_);
  and (_05806_, _00696_, _00695_);
  or (_00697_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00698_, \oc8051_gm_cxrom_1.cell14.data [4], _00672_);
  and (_00699_, _00698_, _00697_);
  or (_00700_, _00699_, rst);
  or (_00701_, \oc8051_gm_cxrom_1.cell14.data [4], _43223_);
  and (_05810_, _00701_, _00700_);
  or (_00702_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00703_, \oc8051_gm_cxrom_1.cell14.data [5], _00672_);
  and (_00704_, _00703_, _00702_);
  or (_00705_, _00704_, rst);
  or (_00706_, \oc8051_gm_cxrom_1.cell14.data [5], _43223_);
  and (_05814_, _00706_, _00705_);
  or (_00707_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00708_, \oc8051_gm_cxrom_1.cell14.data [6], _00672_);
  and (_00709_, _00708_, _00707_);
  or (_00710_, _00709_, rst);
  or (_00711_, \oc8051_gm_cxrom_1.cell14.data [6], _43223_);
  and (_05818_, _00711_, _00710_);
  or (_00712_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_00713_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_00714_, _00713_, \oc8051_gm_cxrom_1.cell15.data [7]);
  and (_00715_, _00714_, _00712_);
  or (_00716_, _00715_, rst);
  or (_00717_, \oc8051_gm_cxrom_1.cell15.data [7], _43223_);
  and (_05840_, _00717_, _00716_);
  or (_00718_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00719_, \oc8051_gm_cxrom_1.cell15.data [0], _00713_);
  and (_00720_, _00719_, _00718_);
  or (_00721_, _00720_, rst);
  or (_00722_, \oc8051_gm_cxrom_1.cell15.data [0], _43223_);
  and (_05847_, _00722_, _00721_);
  or (_00723_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00724_, \oc8051_gm_cxrom_1.cell15.data [1], _00713_);
  and (_00725_, _00724_, _00723_);
  or (_00726_, _00725_, rst);
  or (_00727_, \oc8051_gm_cxrom_1.cell15.data [1], _43223_);
  and (_05851_, _00727_, _00726_);
  or (_00728_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00729_, \oc8051_gm_cxrom_1.cell15.data [2], _00713_);
  and (_00730_, _00729_, _00728_);
  or (_00731_, _00730_, rst);
  or (_00732_, \oc8051_gm_cxrom_1.cell15.data [2], _43223_);
  and (_05855_, _00732_, _00731_);
  or (_00733_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00734_, \oc8051_gm_cxrom_1.cell15.data [3], _00713_);
  and (_00735_, _00734_, _00733_);
  or (_00736_, _00735_, rst);
  or (_00737_, \oc8051_gm_cxrom_1.cell15.data [3], _43223_);
  and (_05859_, _00737_, _00736_);
  or (_00738_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00739_, \oc8051_gm_cxrom_1.cell15.data [4], _00713_);
  and (_00740_, _00739_, _00738_);
  or (_00741_, _00740_, rst);
  or (_00742_, \oc8051_gm_cxrom_1.cell15.data [4], _43223_);
  and (_05863_, _00742_, _00741_);
  or (_00743_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00744_, \oc8051_gm_cxrom_1.cell15.data [5], _00713_);
  and (_00745_, _00744_, _00743_);
  or (_00746_, _00745_, rst);
  or (_00747_, \oc8051_gm_cxrom_1.cell15.data [5], _43223_);
  and (_05867_, _00747_, _00746_);
  or (_00748_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00749_, \oc8051_gm_cxrom_1.cell15.data [6], _00713_);
  and (_00750_, _00749_, _00748_);
  or (_00751_, _00750_, rst);
  or (_00752_, \oc8051_gm_cxrom_1.cell15.data [6], _43223_);
  and (_05871_, _00752_, _00751_);
  nor (_09646_, _38610_, rst);
  and (_00753_, _37083_, _43223_);
  nand (_00754_, _00753_, _38618_);
  nor (_00755_, _38602_, _38573_);
  or (_09649_, _00755_, _00754_);
  and (_00756_, _38566_, _38544_);
  and (_00757_, _00756_, _38522_);
  and (_00758_, _00757_, _38499_);
  and (_00759_, _38243_, _38001_);
  and (_00760_, _37748_, _37476_);
  and (_00761_, _00760_, _00759_);
  and (_00762_, _00761_, _00758_);
  not (_00763_, _38001_);
  and (_00764_, _38243_, _00763_);
  not (_00765_, _37476_);
  not (_00766_, _38566_);
  nor (_00767_, _00766_, _38544_);
  not (_00768_, _38522_);
  and (_00769_, _38499_, _00768_);
  and (_00770_, _00769_, _00767_);
  and (_00771_, _00770_, _00765_);
  and (_00772_, _00771_, _00764_);
  not (_00773_, _38243_);
  and (_00774_, _00773_, _38001_);
  and (_00775_, _00769_, _00756_);
  and (_00776_, _00775_, _37476_);
  and (_00777_, _00776_, _00774_);
  or (_00778_, _00777_, _00772_);
  nor (_00779_, _00778_, _00762_);
  nand (_00780_, _00758_, _00759_);
  or (_00781_, _00760_, _00780_);
  and (_00782_, _37748_, _00765_);
  and (_00783_, _00782_, _00764_);
  and (_00784_, _00775_, _00783_);
  not (_00785_, _37748_);
  nor (_00786_, _38243_, _38001_);
  and (_00787_, _00786_, _00785_);
  and (_00788_, _00787_, _00775_);
  nor (_00789_, _00788_, _00784_);
  and (_00790_, _00789_, _00781_);
  and (_00791_, _00764_, _37748_);
  not (_00792_, _38499_);
  and (_00793_, _00757_, _00792_);
  and (_00794_, _00793_, _00791_);
  and (_00795_, _00786_, _00760_);
  and (_00796_, _00795_, _00766_);
  nor (_00797_, _00796_, _00794_);
  and (_00798_, _00787_, _00757_);
  and (_00799_, _00798_, _00765_);
  and (_00800_, _00767_, _00768_);
  nor (_00801_, _37748_, _00765_);
  and (_00802_, _00801_, _00764_);
  and (_00803_, _00802_, _00800_);
  nor (_00804_, _00803_, _00799_);
  and (_00805_, _00804_, _00797_);
  nor (_00806_, _37748_, _37476_);
  and (_00807_, _00806_, _00759_);
  or (_00808_, _00807_, _00761_);
  and (_00809_, _00808_, _00775_);
  and (_00810_, _00800_, _00792_);
  and (_00811_, _00810_, _00795_);
  nor (_00812_, _00811_, _00809_);
  and (_00813_, _00812_, _00805_);
  and (_00814_, _00756_, _00768_);
  not (_00815_, _00814_);
  and (_00816_, _00774_, _00806_);
  nor (_00817_, _00816_, _00792_);
  nor (_00818_, _00817_, _00815_);
  and (_00819_, _00801_, _00759_);
  and (_00820_, _00819_, _00775_);
  and (_00821_, _00774_, _00782_);
  and (_00822_, _00821_, _00775_);
  nor (_00823_, _00822_, _00820_);
  not (_00824_, _00823_);
  or (_00825_, _00824_, _00818_);
  nor (_00826_, _00768_, _38544_);
  nor (_00827_, _00826_, _00766_);
  not (_00828_, _00827_);
  and (_00829_, _00828_, _00802_);
  and (_00830_, _00801_, _00774_);
  and (_00831_, _00793_, _00830_);
  and (_00832_, _00798_, _37476_);
  or (_00833_, _00832_, _00831_);
  or (_00834_, _00833_, _00829_);
  nor (_00835_, _00834_, _00825_);
  and (_00836_, _00835_, _00813_);
  and (_00837_, _00836_, _00790_);
  nand (_00838_, _00837_, _00779_);
  and (_00839_, _00838_, _37094_);
  not (_00840_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00841_, _37072_, _18789_);
  and (_00842_, _00841_, _38598_);
  nor (_00843_, _00842_, _00840_);
  or (_00844_, _00843_, rst);
  or (_09652_, _00844_, _00839_);
  nand (_00845_, _38001_, _37017_);
  or (_00846_, _37017_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_00847_, _00846_, _43223_);
  and (_09655_, _00847_, _00845_);
  and (_00848_, \oc8051_top_1.oc8051_sfr1.wait_data , _43223_);
  and (_00849_, _00848_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00850_, _38591_, _38619_);
  and (_00851_, _38574_, _38582_);
  and (_00852_, _00851_, _37553_);
  or (_00853_, _00852_, _00850_);
  and (_00854_, _38587_, _38602_);
  or (_00855_, _00854_, _38603_);
  or (_00856_, _00855_, _38681_);
  and (_00857_, _38657_, _38573_);
  and (_00858_, _38574_, _38654_);
  or (_00859_, _00858_, _00857_);
  nor (_00860_, _00859_, _00856_);
  nand (_00861_, _00860_, _38699_);
  or (_00862_, _00861_, _00853_);
  and (_00863_, _00862_, _00753_);
  or (_09658_, _00863_, _00849_);
  and (_00864_, _37553_, _38571_);
  and (_00865_, _00864_, _38653_);
  or (_00866_, _00865_, _38733_);
  and (_00867_, _38615_, _38589_);
  and (_00868_, _00867_, _38654_);
  or (_00869_, _00868_, _00866_);
  nor (_00870_, _38615_, _38548_);
  and (_00871_, _38504_, _38588_);
  and (_00872_, _00871_, _00870_);
  and (_00873_, _00872_, _38342_);
  and (_00874_, _38602_, _38583_);
  or (_00875_, _00874_, _00873_);
  or (_00876_, _00875_, _00869_);
  and (_00877_, _00876_, _37083_);
  and (_00878_, _38708_, _00840_);
  not (_00879_, _38594_);
  and (_00880_, _00879_, _00878_);
  and (_00881_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00882_, _00881_, _00880_);
  or (_00883_, _00882_, _00877_);
  and (_09661_, _00883_, _43223_);
  and (_00884_, _00848_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_00885_, _38591_, _38644_);
  nor (_00886_, _38657_, _38644_);
  nor (_00887_, _00886_, _38630_);
  or (_00888_, _00887_, _00885_);
  and (_00889_, _00867_, _38667_);
  or (_00890_, _00889_, _00888_);
  nor (_00891_, _00886_, _38588_);
  and (_00892_, _37542_, _38571_);
  and (_00893_, _00892_, _38643_);
  or (_00894_, _00893_, _00891_);
  nand (_00895_, _38669_, _38571_);
  nand (_00896_, _00895_, _38725_);
  or (_00897_, _00896_, _00894_);
  and (_00898_, _38591_, _38626_);
  or (_00899_, _00898_, _00875_);
  or (_00900_, _00899_, _00897_);
  or (_00901_, _00900_, _00890_);
  and (_00902_, _00901_, _00753_);
  or (_09664_, _00902_, _00884_);
  and (_00903_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00904_, _38689_, _37083_);
  or (_00905_, _00904_, _00903_);
  or (_00906_, _00905_, _00880_);
  and (_09667_, _00906_, _43223_);
  and (_00907_, _00872_, _38582_);
  and (_00908_, _38602_, _38619_);
  and (_00909_, _38573_, _38619_);
  or (_00910_, _00909_, _00908_);
  or (_00911_, _00910_, _00907_);
  and (_00912_, _00911_, _00878_);
  or (_00913_, _00912_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00914_, _38667_, _38640_);
  and (_00915_, _38572_, _38616_);
  and (_00916_, _00915_, _37542_);
  or (_00917_, _00916_, _00914_);
  and (_00918_, _00917_, _38600_);
  or (_00919_, _00917_, _00852_);
  and (_00920_, _00919_, _37028_);
  or (_00921_, _00920_, _00918_);
  or (_00922_, _00921_, _00913_);
  or (_00923_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18789_);
  and (_00925_, _00923_, _43223_);
  and (_09670_, _00925_, _00922_);
  and (_00926_, _00848_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_00927_, _00892_, _38653_);
  or (_00928_, _00893_, _00927_);
  or (_00929_, _38667_, _38654_);
  and (_00930_, _00929_, _38623_);
  or (_00931_, _00930_, _00928_);
  and (_00932_, _38640_, _38331_);
  or (_00933_, _00889_, _00857_);
  or (_00934_, _00933_, _00932_);
  or (_00935_, _00865_, _38655_);
  or (_00936_, _38575_, _38674_);
  or (_00937_, _00936_, _00935_);
  or (_00938_, _00937_, _00934_);
  or (_00939_, _00938_, _00931_);
  and (_00940_, _00939_, _00753_);
  or (_09673_, _00940_, _00926_);
  and (_00941_, _00848_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_00942_, _00868_, _38670_);
  and (_00943_, _00867_, _38650_);
  and (_00944_, _38574_, _38631_);
  or (_00945_, _00944_, _00943_);
  or (_00946_, _00945_, _00942_);
  or (_00947_, _00946_, _00894_);
  and (_00948_, _38591_, _38664_);
  or (_00949_, _38673_, _38665_);
  or (_00950_, _00949_, _00948_);
  and (_00951_, _38652_, _38624_);
  or (_00952_, _00951_, _38737_);
  and (_00954_, _38657_, _38623_);
  or (_00955_, _00954_, _00952_);
  or (_00956_, _00955_, _00950_);
  or (_00957_, _00956_, _00947_);
  and (_00958_, _00864_, _38652_);
  and (_00959_, _00864_, _38578_);
  or (_00960_, _00959_, _00958_);
  nor (_00961_, _38724_, _38701_);
  nand (_00962_, _00961_, _38679_);
  or (_00963_, _00962_, _00960_);
  or (_00964_, _00963_, _00890_);
  or (_00965_, _00964_, _00957_);
  and (_00966_, _00965_, _00753_);
  or (_09676_, _00966_, _00941_);
  and (_00967_, _00867_, _38632_);
  and (_00968_, _00892_, _38582_);
  or (_00969_, _00968_, _00967_);
  or (_00970_, _00969_, _38719_);
  and (_00971_, _38632_, _38571_);
  or (_00972_, _00971_, _38734_);
  or (_00974_, _00972_, _00970_);
  and (_00975_, _00867_, _38583_);
  or (_00976_, _00975_, _00974_);
  and (_00977_, _00976_, _37083_);
  nand (_00978_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_00979_, _00978_, _38607_);
  or (_00980_, _00979_, _00977_);
  and (_09679_, _00980_, _43223_);
  or (_00981_, _38658_, _38655_);
  not (_00982_, _38702_);
  or (_00983_, _00887_, _00982_);
  or (_00984_, _00983_, _00981_);
  and (_00985_, _38577_, _37542_);
  and (_00986_, _00985_, _38617_);
  or (_00987_, _00986_, _38668_);
  or (_00988_, _00987_, _38665_);
  or (_00989_, _00988_, _00914_);
  nand (_00990_, _38690_, _38682_);
  or (_00991_, _00990_, _00989_);
  or (_00992_, _00991_, _00984_);
  and (_00993_, _00864_, _38582_);
  or (_00994_, _00993_, _00916_);
  and (_00995_, _00892_, _38577_);
  or (_00996_, _00995_, _38646_);
  or (_00997_, _00996_, _00866_);
  or (_00998_, _00997_, _00994_);
  and (_00999_, _00985_, _38623_);
  or (_01000_, _00999_, _38724_);
  or (_01001_, _01000_, _38625_);
  or (_01002_, _38721_, _38686_);
  or (_01003_, _01002_, _01001_);
  or (_01004_, _01003_, _00998_);
  or (_01005_, _01004_, _00894_);
  or (_01006_, _01005_, _00992_);
  and (_01007_, _01006_, _37083_);
  and (_01008_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01009_, _00918_, _00880_);
  and (_01010_, _38600_, _38697_);
  or (_01011_, _01010_, _01009_);
  or (_01012_, _01011_, _01008_);
  or (_01013_, _01012_, _01007_);
  and (_09682_, _01013_, _43223_);
  nor (_09741_, _38746_, rst);
  nor (_09743_, _38712_, rst);
  nand (_09746_, _00911_, _00753_);
  and (_01014_, _38602_, _38618_);
  or (_01015_, _01014_, _00907_);
  nand (_09749_, _01015_, _00753_);
  and (_01016_, _00759_, _00785_);
  and (_01017_, _01016_, _00758_);
  or (_01018_, _00794_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_01019_, _01018_, _01017_);
  or (_01020_, _01019_, _00772_);
  and (_01021_, _01020_, _00842_);
  nor (_01022_, _00841_, _38598_);
  or (_01023_, _01022_, rst);
  or (_09752_, _01023_, _01021_);
  nand (_01024_, _38499_, _37017_);
  or (_01025_, _37017_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_01026_, _01025_, _43223_);
  and (_09755_, _01026_, _01024_);
  not (_01027_, _37017_);
  or (_01028_, _38522_, _01027_);
  or (_01029_, _37017_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_01030_, _01029_, _43223_);
  and (_09758_, _01030_, _01028_);
  nand (_01031_, _38544_, _37017_);
  or (_01032_, _37017_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_01033_, _01032_, _43223_);
  and (_09761_, _01033_, _01031_);
  nand (_01034_, _38566_, _37017_);
  or (_01035_, _37017_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_01036_, _01035_, _43223_);
  and (_09764_, _01036_, _01034_);
  or (_01037_, _37476_, _01027_);
  or (_01038_, _37017_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_01039_, _01038_, _43223_);
  and (_09767_, _01039_, _01037_);
  nand (_01040_, _37748_, _37017_);
  or (_01041_, _37017_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_01042_, _01041_, _43223_);
  and (_09770_, _01042_, _01040_);
  nand (_01043_, _38243_, _37017_);
  or (_01044_, _37017_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_01045_, _01044_, _43223_);
  and (_09773_, _01045_, _01043_);
  or (_01046_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _18789_);
  and (_01047_, _01046_, _43223_);
  and (_01048_, _01047_, _00913_);
  nor (_01049_, _38636_, _38588_);
  or (_01050_, _01049_, _00970_);
  and (_01051_, _00867_, _38664_);
  or (_01052_, _01051_, _00874_);
  or (_01053_, _38657_, _38643_);
  and (_01054_, _01053_, _38591_);
  or (_01055_, _01054_, _01052_);
  or (_01056_, _01055_, _01050_);
  and (_01057_, _00864_, _38618_);
  and (_01058_, _38635_, _38623_);
  or (_01059_, _01058_, _01057_);
  and (_01060_, _00867_, _38635_);
  and (_01061_, _00867_, _38619_);
  or (_01062_, _01061_, _01060_);
  or (_01063_, _01062_, _01059_);
  or (_01064_, _00943_, _38737_);
  or (_01065_, _00959_, _00944_);
  or (_01066_, _01065_, _01064_);
  or (_01067_, _00975_, _38734_);
  and (_01068_, _00864_, _38634_);
  and (_01069_, _00985_, _38591_);
  or (_01070_, _01069_, _01068_);
  or (_01071_, _01070_, _01067_);
  or (_01072_, _38575_, _38728_);
  or (_01073_, _01072_, _01071_);
  or (_01074_, _01073_, _01066_);
  or (_01075_, _01074_, _01063_);
  or (_01076_, _01075_, _01056_);
  and (_01077_, _01076_, _00753_);
  or (_09776_, _01077_, _01048_);
  and (_01078_, _00848_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_01079_, _38664_, _38650_);
  and (_01080_, _01079_, _38640_);
  or (_01081_, _01052_, _00960_);
  or (_01082_, _01081_, _01080_);
  and (_01083_, _37803_, _38309_);
  and (_01084_, _00892_, _01083_);
  and (_01085_, _01084_, _38056_);
  nor (_01086_, _01085_, _38723_);
  not (_01087_, _01086_);
  nor (_01088_, _01087_, _00898_);
  nand (_01089_, _01088_, _38656_);
  or (_01090_, _01089_, _00853_);
  not (_01091_, _38650_);
  nand (_01092_, _01091_, _38636_);
  and (_01093_, _01092_, _38591_);
  or (_01094_, _01093_, _00955_);
  or (_01095_, _01094_, _01090_);
  or (_01096_, _01095_, _01082_);
  and (_01097_, _01096_, _00753_);
  or (_34165_, _01097_, _01078_);
  or (_01098_, _01002_, _00994_);
  or (_01099_, _01098_, _00992_);
  and (_01100_, _01099_, _37083_);
  and (_01101_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01102_, _01101_, _01011_);
  or (_01103_, _01102_, _01100_);
  and (_34167_, _01103_, _43223_);
  and (_01104_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01105_, _01104_, _01009_);
  and (_01106_, _01105_, _43223_);
  and (_01107_, _38700_, _37553_);
  or (_01108_, _01107_, _38733_);
  or (_01109_, _01108_, _01001_);
  or (_01110_, _01109_, _00917_);
  and (_01111_, _01110_, _00753_);
  or (_34170_, _01111_, _01106_);
  and (_01112_, _00892_, _38581_);
  and (_01113_, _01112_, _38056_);
  or (_01114_, _01113_, _38720_);
  or (_01115_, _01114_, _00917_);
  or (_01116_, _00851_, _38593_);
  and (_01117_, _00967_, _37542_);
  or (_01118_, _01117_, _01060_);
  or (_01119_, _01118_, _01116_);
  or (_01120_, _01079_, _38579_);
  and (_01121_, _01120_, _38591_);
  or (_01122_, _01121_, _01119_);
  or (_01123_, _01122_, _01115_);
  and (_01124_, _38591_, _38654_);
  or (_01125_, _00975_, _00944_);
  or (_01126_, _01125_, _01124_);
  or (_01127_, _01126_, _01049_);
  and (_01128_, _00867_, _38669_);
  or (_01129_, _01128_, _00850_);
  and (_01130_, _38618_, _37542_);
  and (_01131_, _01130_, _38591_);
  or (_01132_, _01131_, _38592_);
  or (_01133_, _01132_, _01054_);
  or (_01134_, _01133_, _01129_);
  and (_01135_, _00967_, _37553_);
  or (_01136_, _01135_, _38580_);
  or (_01137_, _00999_, _38734_);
  or (_01138_, _01137_, _00995_);
  and (_01139_, _01130_, _38617_);
  and (_01140_, _38640_, _38635_);
  or (_01141_, _01140_, _01139_);
  or (_01142_, _01141_, _01138_);
  or (_01143_, _01142_, _01136_);
  or (_01144_, _01143_, _01134_);
  or (_01145_, _01144_, _01127_);
  or (_01146_, _01145_, _01123_);
  and (_01147_, _01146_, _37083_);
  and (_01148_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_01149_, _38594_, _37028_);
  or (_01150_, _00912_, _01149_);
  or (_01151_, _01150_, _01148_);
  or (_01152_, _01151_, _01147_);
  and (_34172_, _01152_, _43223_);
  and (_01153_, _00892_, _38618_);
  or (_01154_, _00986_, _00874_);
  or (_01155_, _01154_, _01153_);
  or (_01156_, _01155_, _38585_);
  and (_01157_, _01079_, _38574_);
  or (_01158_, _01157_, _38637_);
  or (_01159_, _01158_, _01156_);
  and (_01160_, _01130_, _38623_);
  or (_01161_, _38593_, _38734_);
  or (_01162_, _01161_, _38686_);
  or (_01163_, _01162_, _01160_);
  or (_01164_, _01163_, _01114_);
  or (_01165_, _01164_, _01159_);
  or (_01166_, _01134_, _01127_);
  or (_01167_, _01166_, _01165_);
  and (_01168_, _01167_, _37083_);
  and (_01169_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01170_, _01169_, _01150_);
  or (_01171_, _01170_, _01168_);
  and (_34174_, _01171_, _43223_);
  and (_01172_, _00848_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_01173_, _38574_, _38657_);
  and (_01174_, _38574_, _38643_);
  and (_01175_, _01174_, _37542_);
  or (_01176_, _01175_, _01173_);
  not (_01177_, _42725_);
  or (_01178_, _00975_, _01177_);
  or (_01179_, _01178_, _00931_);
  or (_01180_, _01179_, _01176_);
  or (_01181_, _00981_, _00936_);
  or (_01182_, _38622_, _38571_);
  or (_01183_, _01182_, _38574_);
  and (_01184_, _01183_, _38692_);
  and (_01185_, _38591_, _38657_);
  or (_01186_, _01185_, _00889_);
  or (_01187_, _01186_, _01184_);
  or (_01188_, _01187_, _01181_);
  or (_01189_, _01113_, _00865_);
  and (_01190_, _38574_, _38669_);
  or (_01191_, _01190_, _01117_);
  or (_01192_, _01191_, _01189_);
  nor (_01193_, _38734_, _38688_);
  nand (_01194_, _01193_, _42724_);
  or (_01195_, _01194_, _01192_);
  or (_01196_, _01195_, _01188_);
  or (_01197_, _01196_, _01180_);
  and (_01198_, _01197_, _00753_);
  or (_34176_, _01198_, _01172_);
  or (_01199_, _00868_, _38678_);
  or (_01200_, _00954_, _00951_);
  or (_01201_, _01200_, _01199_);
  or (_01202_, _01201_, _00950_);
  or (_01203_, _01202_, _01119_);
  and (_01204_, _38574_, _38692_);
  or (_01205_, _01204_, _01185_);
  or (_01206_, _01175_, _01136_);
  or (_01207_, _01206_, _01205_);
  or (_01208_, _00958_, _38575_);
  or (_01209_, _01208_, _38720_);
  not (_01210_, _38687_);
  or (_01211_, _01049_, _01210_);
  or (_01212_, _01211_, _01209_);
  or (_01213_, _01212_, _01207_);
  or (_01214_, _01213_, _01203_);
  and (_01216_, _01214_, _00753_);
  and (_01218_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01220_, _38593_, _37039_);
  or (_01222_, _01220_, _01218_);
  and (_01224_, _01222_, _43223_);
  or (_34178_, _01224_, _01216_);
  and (_01227_, _38573_, _38669_);
  or (_01229_, _01227_, _01131_);
  nor (_01231_, _00975_, _38677_);
  nand (_01233_, _01231_, _38735_);
  or (_01235_, _01233_, _01129_);
  or (_01237_, _01235_, _01229_);
  or (_01239_, _01060_, _38686_);
  or (_01241_, _01239_, _38685_);
  or (_01243_, _01189_, _00868_);
  and (_01245_, _38574_, _38632_);
  and (_01247_, _01182_, _38635_);
  or (_01249_, _01247_, _01245_);
  or (_01251_, _01249_, _01243_);
  or (_01253_, _01251_, _01241_);
  or (_01255_, _01253_, _01237_);
  or (_01257_, _00897_, _00890_);
  or (_01259_, _01257_, _01255_);
  and (_01261_, _01259_, _37083_);
  and (_01263_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01265_, _01263_, _38605_);
  or (_01267_, _01265_, _01261_);
  and (_34180_, _01267_, _43223_);
  or (_01270_, _01239_, _01186_);
  or (_01272_, _01270_, _01229_);
  or (_01274_, _38733_, _38724_);
  or (_01276_, _01274_, _01174_);
  or (_01278_, _01276_, _01247_);
  or (_01280_, _00935_, _01177_);
  or (_01282_, _01280_, _01278_);
  or (_01284_, _00894_, _00888_);
  or (_01286_, _01284_, _01282_);
  or (_01288_, _01286_, _01272_);
  and (_01290_, _01288_, _37083_);
  and (_01292_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01294_, _01292_, _38606_);
  or (_01296_, _01294_, _01290_);
  and (_34182_, _01296_, _43223_);
  and (_01299_, _00848_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_01301_, _00858_, _38659_);
  nand (_01303_, _01301_, _42724_);
  not (_01305_, _38572_);
  or (_01307_, _38574_, _01305_);
  and (_01309_, _01307_, _38669_);
  or (_01310_, _01309_, _01205_);
  or (_01311_, _01310_, _01303_);
  or (_01312_, _01178_, _00974_);
  or (_01313_, _01312_, _01176_);
  or (_01314_, _01313_, _01311_);
  and (_01315_, _01314_, _00753_);
  or (_34184_, _01315_, _01299_);
  nor (_39248_, _38001_, rst);
  nor (_39249_, _42658_, rst);
  and (_01316_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_01317_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_01318_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_01319_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_01320_, _01319_, _01318_);
  and (_01321_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01322_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_01323_, _01322_, _01321_);
  and (_01324_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_01325_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_01326_, _01325_, _01324_);
  and (_01327_, _01326_, _01323_);
  and (_01328_, _01327_, _01320_);
  nor (_01329_, _01328_, _37269_);
  nor (_01330_, _01329_, _01317_);
  nor (_01331_, _01330_, _42642_);
  nor (_01332_, _01331_, _01316_);
  nor (_39251_, _01332_, rst);
  nor (_39261_, _38499_, rst);
  and (_39263_, _38522_, _43223_);
  nor (_39264_, _38544_, rst);
  nor (_39265_, _38566_, rst);
  and (_39266_, _37476_, _43223_);
  nor (_39267_, _37748_, rst);
  nor (_39268_, _38243_, rst);
  nor (_39269_, _42932_, rst);
  nor (_39270_, _42807_, rst);
  nor (_39272_, _43055_, rst);
  nor (_39273_, _42888_, rst);
  nor (_39274_, _42753_, rst);
  nor (_39275_, _43009_, rst);
  nor (_39276_, _42985_, rst);
  and (_01333_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_01334_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_01335_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_01336_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01337_, _01336_, _01335_);
  and (_01338_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_01339_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01340_, _01339_, _01338_);
  and (_01341_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01342_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_01343_, _01342_, _01341_);
  and (_01344_, _01343_, _01340_);
  and (_01345_, _01344_, _01337_);
  nor (_01346_, _01345_, _37269_);
  nor (_01347_, _01346_, _01334_);
  nor (_01348_, _01347_, _42642_);
  nor (_01349_, _01348_, _01333_);
  nor (_39278_, _01349_, rst);
  and (_01350_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_01351_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_01352_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01353_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01354_, _01353_, _01352_);
  and (_01355_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_01356_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_01357_, _01356_, _01355_);
  and (_01358_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_01359_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_01360_, _01359_, _01358_);
  and (_01361_, _01360_, _01357_);
  and (_01362_, _01361_, _01354_);
  nor (_01363_, _01362_, _37269_);
  nor (_01364_, _01363_, _01351_);
  nor (_01365_, _01364_, _42642_);
  nor (_01366_, _01365_, _01350_);
  nor (_39279_, _01366_, rst);
  and (_01367_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_01368_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_01369_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_01370_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01371_, _01370_, _01369_);
  and (_01372_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_01373_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_01374_, _01373_, _01372_);
  and (_01375_, _01374_, _01371_);
  and (_01376_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_01377_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01378_, _01377_, _01376_);
  and (_01379_, _01378_, _01375_);
  nor (_01380_, _01379_, _37269_);
  nor (_01381_, _01380_, _01368_);
  nor (_01382_, _01381_, _42642_);
  nor (_01383_, _01382_, _01367_);
  nor (_39280_, _01383_, rst);
  and (_01384_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_01385_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_01386_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_01387_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01388_, _01387_, _01386_);
  and (_01389_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_01390_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01391_, _01390_, _01389_);
  and (_01392_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_01393_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_01394_, _01393_, _01392_);
  and (_01395_, _01394_, _01391_);
  and (_01396_, _01395_, _01388_);
  nor (_01397_, _01396_, _37269_);
  nor (_01398_, _01397_, _01385_);
  nor (_01399_, _01398_, _42642_);
  nor (_01400_, _01399_, _01384_);
  nor (_39281_, _01400_, rst);
  and (_01401_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_01402_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_01403_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_01404_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01405_, _01404_, _01403_);
  and (_01406_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_01407_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_01408_, _01407_, _01406_);
  and (_01409_, _01408_, _01405_);
  and (_01410_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_01411_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01412_, _01411_, _01410_);
  and (_01413_, _01412_, _01409_);
  nor (_01414_, _01413_, _37269_);
  nor (_01415_, _01414_, _01402_);
  nor (_01416_, _01415_, _42642_);
  nor (_01417_, _01416_, _01401_);
  nor (_39282_, _01417_, rst);
  and (_01418_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_01419_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_01420_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_01421_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01422_, _01421_, _01420_);
  and (_01423_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_01424_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_01425_, _01424_, _01423_);
  and (_01426_, _01425_, _01422_);
  and (_01427_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_01428_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01429_, _01428_, _01427_);
  and (_01430_, _01429_, _01426_);
  nor (_01431_, _01430_, _37269_);
  nor (_01432_, _01431_, _01419_);
  nor (_01433_, _01432_, _42642_);
  nor (_01434_, _01433_, _01418_);
  nor (_39284_, _01434_, rst);
  and (_01435_, _42642_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_01436_, _37269_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_01437_, _37182_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_01438_, _37302_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01439_, _01438_, _01437_);
  and (_01440_, _37356_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_01441_, _37226_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_01442_, _01441_, _01440_);
  and (_01443_, _01442_, _01439_);
  and (_01444_, _37335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_01445_, _37149_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01446_, _01445_, _01444_);
  and (_01447_, _01446_, _01443_);
  nor (_01448_, _01447_, _37269_);
  nor (_01449_, _01448_, _01436_);
  nor (_01450_, _01449_, _42642_);
  nor (_01451_, _01450_, _01435_);
  nor (_39285_, _01451_, rst);
  and (_01452_, _37094_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_01453_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_01454_, _01452_, _38888_);
  and (_01455_, _01454_, _43223_);
  and (_39310_, _01455_, _01453_);
  not (_01456_, _01452_);
  or (_01457_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _01452_, _43223_);
  and (_01458_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _43223_);
  or (_01459_, _01458_, _00000_);
  and (_39311_, _01459_, _01457_);
  nor (_39346_, _42721_, rst);
  nor (_39349_, _42716_, rst);
  not (_01460_, _38710_);
  not (_01461_, _38600_);
  nor (_01462_, _01461_, _38699_);
  not (_01463_, _01462_);
  and (_01464_, _38604_, _38633_);
  nor (_01465_, _01464_, _42734_);
  and (_01466_, _01465_, _01463_);
  and (_01467_, _01466_, _38614_);
  not (_01468_, _34896_);
  nand (_01469_, _34124_, _29609_);
  nor (_01470_, _01469_, _32034_);
  and (_01471_, _01470_, _01468_);
  and (_01472_, _01471_, _35625_);
  and (_01473_, _01472_, _36365_);
  and (_01474_, _01473_, _01467_);
  and (_01475_, _01474_, _29773_);
  and (_01476_, _01464_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_01477_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_01478_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01479_, _01478_, _01477_);
  nor (_01480_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_01481_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01482_, _01481_, _01480_);
  and (_01483_, _01482_, _01479_);
  and (_01484_, _01483_, _38744_);
  nor (_01485_, _01484_, _01476_);
  not (_01486_, _01485_);
  nor (_01487_, _01486_, _01475_);
  nor (_01488_, _01466_, _01464_);
  and (_01489_, _01488_, _29477_);
  not (_01490_, _01489_);
  and (_01491_, _01490_, _01487_);
  nor (_01492_, _01128_, _38674_);
  and (_01493_, _01492_, _01086_);
  or (_01494_, _38692_, _38579_);
  or (_01495_, _01494_, _38635_);
  and (_01496_, _01495_, _38602_);
  nor (_01497_, _01496_, _00927_);
  and (_01498_, _01497_, _01493_);
  and (_01499_, _01498_, _01491_);
  and (_01500_, _38603_, _37553_);
  not (_01501_, _01500_);
  and (_01502_, _01501_, _38698_);
  not (_01503_, _01502_);
  nor (_01504_, _01503_, _01491_);
  nor (_01505_, _01504_, _01499_);
  nor (_01506_, _00854_, _38580_);
  and (_01507_, _01506_, _38642_);
  not (_01508_, _01507_);
  nor (_01509_, _01508_, _01505_);
  nor (_01510_, _01509_, _01461_);
  and (_01511_, _38643_, _38640_);
  nor (_01512_, _01511_, _00915_);
  nor (_01513_, _01512_, _37039_);
  nor (_01514_, _01513_, _38710_);
  not (_01515_, _01514_);
  nor (_01516_, _01515_, _01510_);
  not (_01517_, _39231_);
  or (_01518_, _39243_, _01517_);
  and (_01519_, _01518_, _01464_);
  not (_01520_, _39511_);
  and (_01521_, _01520_, _38744_);
  or (_01522_, _01521_, _01519_);
  nor (_01523_, _01522_, _01516_);
  not (_01524_, _01523_);
  nor (_01525_, _42892_, _28282_);
  and (_01526_, _42892_, _28282_);
  nor (_01527_, _01526_, _01525_);
  not (_01528_, _01527_);
  nor (_01529_, _42989_, _27821_);
  and (_01530_, _42989_, _27821_);
  nor (_01531_, _01530_, _01529_);
  nor (_01532_, _01531_, _43117_);
  nor (_01533_, _43039_, _27953_);
  and (_01534_, _43039_, _27953_);
  nor (_01535_, _01534_, _01533_);
  nor (_01536_, _42788_, _28424_);
  and (_01537_, _42788_, _28424_);
  nor (_01538_, _01537_, _01536_);
  nor (_01539_, _01538_, _01535_);
  and (_01540_, _01539_, _01532_);
  and (_01541_, _01540_, _01528_);
  nor (_01542_, _31882_, _40230_);
  and (_01543_, _01542_, _01541_);
  and (_01544_, _01543_, _01488_);
  nor (_01545_, _01544_, _01524_);
  and (_01546_, _42835_, _33928_);
  nor (_01547_, _42835_, _33928_);
  or (_01548_, _01547_, _01546_);
  nor (_01549_, _42936_, _33177_);
  and (_01550_, _42936_, _33177_);
  nor (_01551_, _01550_, _01549_);
  not (_01552_, _01551_);
  nor (_01553_, _01552_, _01548_);
  nor (_01554_, _43084_, _31860_);
  and (_01555_, _43084_, _31860_);
  nor (_01556_, _01555_, _01554_);
  and (_01557_, _01556_, _01528_);
  and (_01558_, _01557_, _01553_);
  and (_01559_, _01558_, _01540_);
  and (_01560_, _01559_, _31260_);
  nor (_01561_, _28128_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_01562_, _01561_, _01560_);
  not (_01563_, _01562_);
  and (_01564_, _01563_, _01545_);
  and (_01565_, _01564_, _01460_);
  and (_39353_, _01565_, _43223_);
  and (_39354_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _43223_);
  and (_39355_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _43223_);
  nor (_01566_, _01460_, _31194_);
  not (_01567_, _38973_);
  and (_01568_, _38580_, _38600_);
  and (_01569_, _01568_, _01567_);
  nor (_01570_, _01493_, _01461_);
  not (_01571_, _01570_);
  and (_01572_, _01511_, _37028_);
  not (_01573_, _01572_);
  and (_01574_, _38602_, _38632_);
  and (_01575_, _01574_, _37028_);
  nor (_01576_, _01575_, _38710_);
  and (_01577_, _01576_, _01573_);
  and (_01578_, _01577_, _01463_);
  and (_01579_, _01578_, _01571_);
  and (_01580_, _01579_, _01513_);
  and (_01581_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01582_, _01581_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01583_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01584_, _01583_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01585_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01586_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01587_, _01586_, _01585_);
  and (_01588_, _01587_, _01584_);
  and (_01589_, _01588_, _01582_);
  and (_01590_, _01589_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01591_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01592_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_01593_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01594_, _01593_, _38888_);
  or (_01595_, _01593_, _38888_);
  and (_01596_, _01595_, _01594_);
  and (_01597_, _01596_, _01580_);
  nor (_01598_, _00927_, _38603_);
  and (_01599_, _01598_, _01506_);
  nand (_01600_, _01599_, _01493_);
  and (_01601_, _01600_, _38600_);
  or (_01602_, _01575_, _01462_);
  or (_01603_, _01602_, _01601_);
  nor (_01604_, _01568_, _01513_);
  nand (_01605_, _01604_, _01579_);
  nor (_01606_, _01605_, _01603_);
  and (_01607_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01608_, _01572_, _42659_);
  or (_01609_, _01608_, _01607_);
  or (_01610_, _01609_, _01597_);
  or (_01611_, _01610_, _01569_);
  or (_01613_, _01611_, _01566_);
  and (_01614_, _01579_, _42659_);
  nor (_01616_, _01579_, _01332_);
  nor (_01617_, _01616_, _01614_);
  not (_01619_, _01617_);
  not (_01620_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_01622_, _01617_, _01620_);
  and (_01623_, _01617_, _01620_);
  not (_01625_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01626_, _01579_, _42986_);
  nor (_01628_, _01579_, _01451_);
  nor (_01629_, _01628_, _01626_);
  nor (_01631_, _01629_, _01625_);
  and (_01632_, _01629_, _01625_);
  nor (_01634_, _01632_, _01631_);
  not (_01635_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01637_, _01579_, _43010_);
  nor (_01638_, _01579_, _01434_);
  nor (_01640_, _01638_, _01637_);
  nor (_01641_, _01640_, _01635_);
  and (_01643_, _01640_, _01635_);
  not (_01644_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01645_, _01579_, _42754_);
  nor (_01646_, _01579_, _01417_);
  nor (_01647_, _01646_, _01645_);
  or (_01648_, _01647_, _01644_);
  not (_01649_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01650_, _01579_, _42889_);
  nor (_01651_, _01579_, _01400_);
  nor (_01652_, _01651_, _01650_);
  nor (_01653_, _01652_, _01649_);
  and (_01654_, _01652_, _01649_);
  not (_01655_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01656_, _01579_, _43056_);
  nor (_01657_, _01579_, _01383_);
  nor (_01658_, _01657_, _01656_);
  nor (_01659_, _01658_, _01655_);
  not (_01660_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01661_, _01579_, _42808_);
  nor (_01662_, _01579_, _01366_);
  nor (_01663_, _01662_, _01661_);
  nor (_01664_, _01663_, _01660_);
  and (_01665_, _01579_, _42932_);
  not (_01666_, _01579_);
  and (_01667_, _01666_, _01349_);
  nor (_01668_, _01667_, _01665_);
  and (_01669_, _01668_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_01670_, _01663_, _01660_);
  nor (_01671_, _01670_, _01664_);
  and (_01672_, _01671_, _01669_);
  nor (_01673_, _01672_, _01664_);
  not (_01674_, _01673_);
  and (_01675_, _01658_, _01655_);
  nor (_01676_, _01675_, _01659_);
  and (_01677_, _01676_, _01674_);
  nor (_01678_, _01677_, _01659_);
  nor (_01679_, _01678_, _01654_);
  or (_01680_, _01679_, _01653_);
  nand (_01681_, _01647_, _01644_);
  and (_01682_, _01681_, _01648_);
  nand (_01683_, _01682_, _01680_);
  and (_01684_, _01683_, _01648_);
  nor (_01685_, _01684_, _01643_);
  or (_01686_, _01685_, _01641_);
  and (_01687_, _01686_, _01634_);
  nor (_01688_, _01687_, _01631_);
  nor (_01689_, _01688_, _01623_);
  or (_01690_, _01689_, _01622_);
  and (_01691_, _01690_, _01582_);
  and (_01692_, _01691_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01693_, _01692_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01694_, _01693_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_01695_, _01694_, _01619_);
  nor (_01696_, _01690_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01697_, _01696_, _38910_);
  and (_01698_, _01697_, _38915_);
  and (_01699_, _01698_, _38900_);
  and (_01700_, _01699_, _38921_);
  and (_01701_, _01700_, _38896_);
  nor (_01702_, _01701_, _01617_);
  nor (_01703_, _01702_, _01695_);
  or (_01704_, _01617_, _38892_);
  nand (_01705_, _01617_, _38892_);
  and (_01706_, _01705_, _01704_);
  and (_01707_, _01706_, _01703_);
  or (_01708_, _01707_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_01709_, _01707_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_01710_, _01709_, _01708_);
  or (_01711_, _01604_, _01666_);
  and (_01712_, _38602_, _37028_);
  and (_01713_, _01712_, _38632_);
  or (_01714_, _01713_, _01462_);
  or (_01715_, _01714_, _01601_);
  and (_01716_, _01715_, _01711_);
  and (_01717_, _01716_, _01710_);
  or (_01718_, _01717_, _01613_);
  and (_01719_, _01718_, _01564_);
  nor (_01720_, _37171_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01721_, _01720_, _42642_);
  nor (_01722_, _01721_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_01723_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01725_, _01724_, _01723_);
  not (_01726_, _01725_);
  nor (_01727_, _01726_, _01722_);
  and (_01728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_01729_, _01728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01730_, _01729_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01731_, _01730_, _01727_);
  and (_01732_, _01731_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01733_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01734_, _01733_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01735_, _01734_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_01736_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01737_, _01736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_01738_, _01736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_01739_, _01738_, _01737_);
  nor (_01740_, _01739_, _01564_);
  or (_01741_, _01740_, _01719_);
  and (_39356_, _01741_, _43223_);
  and (_01742_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _43223_);
  and (_01743_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01744_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_01745_, _37083_, _01744_);
  not (_01746_, _01745_);
  not (_01747_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_01748_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01750_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01751_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_01752_, _01751_, _01749_);
  and (_01753_, _01752_, _01750_);
  nor (_01754_, _01753_, _01749_);
  nor (_01755_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01756_, _01755_, _01748_);
  not (_01757_, _01756_);
  nor (_01758_, _01757_, _01754_);
  nor (_01759_, _01758_, _01748_);
  not (_01760_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01761_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_01762_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01763_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_01764_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_01765_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_01766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01767_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_01768_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_01769_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01770_, _01769_, _01768_);
  and (_01771_, _01770_, _01767_);
  and (_01772_, _01771_, _01766_);
  and (_01773_, _01772_, _01765_);
  and (_01774_, _01773_, _01764_);
  and (_01775_, _01774_, _01763_);
  and (_01776_, _01775_, _01762_);
  and (_01777_, _01776_, _01761_);
  and (_01778_, _01777_, _01760_);
  and (_01779_, _01778_, _01759_);
  and (_01780_, _01779_, _01747_);
  nor (_01781_, _01780_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01782_, _01780_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_01783_, _01782_, _01781_);
  nor (_01784_, _01779_, _01747_);
  nor (_01785_, _01784_, _01780_);
  not (_01786_, _01785_);
  and (_01787_, _01777_, _01759_);
  nor (_01788_, _01787_, _01760_);
  or (_01789_, _01788_, _01779_);
  and (_01790_, _01776_, _01759_);
  nor (_01791_, _01790_, _01761_);
  nor (_01792_, _01791_, _01787_);
  not (_01793_, _01792_);
  and (_01794_, _01774_, _01759_);
  and (_01795_, _01794_, _01763_);
  nor (_01796_, _01795_, _01762_);
  nor (_01797_, _01796_, _01790_);
  not (_01798_, _01797_);
  nor (_01799_, _01794_, _01763_);
  nor (_01800_, _01799_, _01795_);
  not (_01801_, _01800_);
  and (_01802_, _01773_, _01759_);
  nor (_01803_, _01802_, _01764_);
  nor (_01804_, _01803_, _01794_);
  not (_01805_, _01804_);
  and (_01806_, _01771_, _01759_);
  nor (_01807_, _01806_, _01766_);
  and (_01808_, _01772_, _01759_);
  or (_01809_, _01808_, _01807_);
  and (_01810_, _01770_, _01759_);
  nor (_01811_, _01810_, _01767_);
  nor (_01812_, _01811_, _01806_);
  not (_01813_, _01812_);
  and (_01814_, _01769_, _01759_);
  nor (_01815_, _01814_, _01768_);
  nor (_01816_, _01815_, _01810_);
  not (_01817_, _01816_);
  not (_01818_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01819_, _01759_, _01818_);
  nor (_01820_, _01759_, _01818_);
  nor (_01821_, _01820_, _01819_);
  not (_01822_, _01821_);
  and (_01823_, _00764_, _00760_);
  and (_01824_, _01823_, _00800_);
  or (_01825_, _00770_, _00758_);
  not (_01826_, _00758_);
  nor (_01827_, _00795_, _00830_);
  nor (_01828_, _01827_, _01826_);
  or (_01829_, _01828_, _00821_);
  and (_01830_, _01829_, _01825_);
  nor (_01831_, _01830_, _01824_);
  not (_01832_, _00816_);
  nor (_01833_, _00800_, _00757_);
  or (_01834_, _01833_, _01832_);
  or (_01835_, _00796_, _00784_);
  or (_01836_, _01835_, _00777_);
  nor (_01837_, _01836_, _00825_);
  and (_01838_, _01837_, _01834_);
  and (_01839_, _01838_, _01831_);
  and (_01840_, _00810_, _00802_);
  and (_01841_, _00774_, _00760_);
  and (_01842_, _00793_, _01841_);
  or (_01843_, _01842_, _01840_);
  and (_01844_, _00759_, _37748_);
  and (_01845_, _00810_, _01844_);
  nor (_01846_, _01845_, _01843_);
  or (_01847_, _00830_, _00783_);
  and (_01848_, _01847_, _00810_);
  and (_01849_, _00806_, _00764_);
  or (_01850_, _01823_, _01849_);
  and (_01851_, _01850_, _00758_);
  nor (_01852_, _01851_, _01848_);
  and (_01853_, _00786_, _00782_);
  nor (_01854_, _01853_, _00802_);
  or (_01855_, _01854_, _01826_);
  nand (_01856_, _01016_, _00810_);
  and (_01857_, _01856_, _01855_);
  and (_01858_, _01844_, _00758_);
  not (_01859_, _01858_);
  and (_01860_, _00786_, _00801_);
  or (_01861_, _00821_, _01860_);
  nand (_01862_, _01861_, _00810_);
  and (_01863_, _01862_, _01859_);
  and (_01864_, _01863_, _01857_);
  and (_01865_, _01864_, _01852_);
  and (_01866_, _01865_, _01846_);
  and (_01867_, _01866_, _01839_);
  and (_01868_, _00802_, _00775_);
  and (_01869_, _00830_, _00770_);
  nor (_01870_, _01869_, _01868_);
  and (_01871_, _01823_, _00775_);
  and (_01872_, _00786_, _00806_);
  and (_01873_, _00810_, _01872_);
  nor (_01874_, _01873_, _01871_);
  and (_01875_, _01874_, _01870_);
  and (_01876_, _01853_, _00810_);
  and (_01877_, _00821_, _00793_);
  or (_01878_, _01877_, _01876_);
  nor (_01879_, _01878_, _00829_);
  and (_01880_, _01879_, _01875_);
  and (_01881_, _00826_, _38566_);
  and (_01882_, _01881_, _00830_);
  and (_01883_, _00783_, _00758_);
  and (_01884_, _00819_, _00770_);
  or (_01885_, _01884_, _01883_);
  nor (_01886_, _01885_, _01882_);
  and (_01887_, _01016_, _00771_);
  and (_01888_, _00764_, _00765_);
  and (_01889_, _01888_, _01881_);
  nor (_01890_, _01889_, _01887_);
  and (_01891_, _01890_, _01886_);
  and (_01892_, _00802_, _00770_);
  not (_01893_, _01892_);
  and (_01894_, _01893_, _00812_);
  not (_01895_, _00775_);
  and (_01896_, _00786_, _37748_);
  nor (_01897_, _01896_, _01849_);
  nor (_01898_, _01897_, _01895_);
  or (_01899_, _01825_, _00810_);
  and (_01900_, _01899_, _01841_);
  nor (_01901_, _01900_, _01898_);
  and (_01902_, _01901_, _01894_);
  nor (_01903_, _00830_, _01849_);
  nor (_01904_, _01903_, _38566_);
  and (_01905_, _00783_, _00766_);
  nor (_01906_, _01905_, _01904_);
  and (_01907_, _01906_, _01902_);
  and (_01908_, _01907_, _01891_);
  and (_01909_, _01908_, _01880_);
  and (_01910_, _01909_, _01867_);
  nor (_01911_, _01752_, _01750_);
  nor (_01912_, _01911_, _01753_);
  not (_01913_, _01912_);
  nor (_01914_, _01913_, _01910_);
  not (_01915_, _01914_);
  or (_01916_, _00829_, _01858_);
  or (_01917_, _01916_, _01848_);
  or (_01918_, _01917_, _01843_);
  and (_01919_, _00816_, _00793_);
  or (_01920_, _01877_, _00820_);
  or (_01921_, _01920_, _01871_);
  nor (_01922_, _01921_, _01919_);
  nand (_01923_, _01922_, _01894_);
  or (_01924_, _01923_, _01918_);
  nor (_01925_, _01924_, _01910_);
  not (_01926_, _01925_);
  nor (_01927_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01928_, _01927_, _01750_);
  and (_01929_, _01928_, _01926_);
  and (_01930_, _01913_, _01910_);
  nor (_01931_, _01930_, _01914_);
  nand (_01932_, _01931_, _01929_);
  and (_01933_, _01932_, _01915_);
  not (_01934_, _01933_);
  and (_01935_, _01757_, _01754_);
  nor (_01936_, _01935_, _01758_);
  and (_01937_, _01936_, _01934_);
  and (_01938_, _01937_, _01822_);
  not (_01939_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_01940_, _01819_, _01939_);
  or (_01941_, _01940_, _01814_);
  and (_01942_, _01941_, _01938_);
  and (_01943_, _01942_, _01817_);
  and (_01944_, _01943_, _01813_);
  and (_01945_, _01944_, _01809_);
  nor (_01946_, _01808_, _01765_);
  or (_01947_, _01946_, _01802_);
  and (_01948_, _01947_, _01945_);
  and (_01949_, _01948_, _01805_);
  and (_01950_, _01949_, _01801_);
  and (_01951_, _01950_, _01798_);
  and (_01952_, _01951_, _01793_);
  and (_01953_, _01952_, _01789_);
  and (_01954_, _01953_, _01786_);
  or (_01955_, _01954_, _01783_);
  nand (_01956_, _01954_, _01783_);
  and (_01957_, _01956_, _01955_);
  or (_01958_, _01957_, _01746_);
  or (_01959_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_01960_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01961_, _01960_, _01959_);
  and (_01962_, _01961_, _01958_);
  or (_39358_, _01962_, _01743_);
  nor (_01963_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_39359_, _01963_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_39360_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _43223_);
  nor (_01964_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01966_, _01965_, _01964_);
  nor (_01967_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_01968_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_01969_, _01968_, _01967_);
  and (_01970_, _01969_, _01966_);
  nor (_01971_, _01970_, rst);
  and (_01972_, \oc8051_top_1.oc8051_rom1.ea_int , _37050_);
  nand (_01973_, _01972_, _37083_);
  and (_01974_, _01973_, _39360_);
  or (_39361_, _01974_, _01971_);
  and (_01975_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_01976_, _01975_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_39363_, _01976_, _43223_);
  nor (_01977_, _01722_, _42642_);
  nor (_01978_, _01910_, _37280_);
  not (_01979_, _01978_);
  nor (_01980_, _01925_, _37204_);
  and (_01981_, _01910_, _37280_);
  nor (_01982_, _01981_, _01978_);
  nand (_01983_, _01982_, _01980_);
  and (_01984_, _01983_, _01979_);
  nor (_01985_, _01984_, _42642_);
  and (_01986_, _01985_, _37127_);
  nor (_01987_, _01985_, _37127_);
  nor (_01988_, _01987_, _01986_);
  nor (_01989_, _01988_, _01977_);
  and (_01990_, _37291_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01991_, _01990_, _01977_);
  and (_01992_, _01991_, _01924_);
  or (_01993_, _01992_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01994_, _01993_, _01989_);
  and (_39364_, _01994_, _43223_);
  nor (_01995_, _37400_, _38516_);
  and (_01996_, _38199_, _37957_);
  and (_01997_, _01996_, _01995_);
  and (_01998_, _37094_, _43223_);
  nand (_01999_, _01998_, _38540_);
  nor (_02000_, _01999_, _38494_);
  not (_02001_, _38562_);
  and (_02002_, _37706_, _02001_);
  and (_02003_, _02002_, _02000_);
  and (_39367_, _02003_, _01997_);
  nor (_02004_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_02005_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_02006_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_39370_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _43223_);
  and (_02007_, _39370_, _02006_);
  or (_39368_, _02007_, _02005_);
  not (_02008_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_02009_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_02010_, _02009_, _02008_);
  and (_02011_, _02009_, _02008_);
  nor (_02012_, _02011_, _02010_);
  not (_02013_, _02012_);
  and (_02014_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_02015_, _02014_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_02016_, _02014_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_02017_, _02016_, _02015_);
  or (_02018_, _02017_, _02009_);
  and (_02019_, _02018_, _02013_);
  nor (_02020_, _02010_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_02021_, _02010_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_02022_, _02021_, _02020_);
  or (_02023_, _02015_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_39372_, _02023_, _43223_);
  and (_02024_, _39372_, _02022_);
  and (_39371_, _02024_, _02019_);
  not (_02025_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_02026_, _01722_, _02025_);
  and (_02027_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_02028_, _02026_);
  and (_02029_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_02030_, _02029_, _02027_);
  and (_39373_, _02030_, _43223_);
  and (_02031_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_02032_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_02033_, _02032_, _02031_);
  and (_39374_, _02033_, _43223_);
  and (_02034_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_02035_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02036_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _02035_);
  and (_02037_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_02038_, _02037_, _02034_);
  and (_39375_, _02038_, _43223_);
  and (_02039_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02040_, _02039_, _02036_);
  and (_39376_, _02040_, _43223_);
  or (_02041_, _02035_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_39378_, _02041_, _43223_);
  not (_02042_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_02043_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_02044_, _02043_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02045_, _02035_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_02046_, _02045_, _43223_);
  and (_39379_, _02046_, _02044_);
  or (_02047_, _02035_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_39380_, _02047_, _43223_);
  nor (_02048_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_02049_, _02048_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02050_, _02049_, _43223_);
  and (_02051_, _39370_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_39381_, _02051_, _02050_);
  and (_02052_, _02025_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_02053_, _02052_, _02049_);
  and (_39382_, _02053_, _43223_);
  nand (_02054_, _02049_, _38973_);
  or (_02055_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_02056_, _02055_, _43223_);
  and (_39383_, _02056_, _02054_);
  nand (_02057_, _38612_, _43223_);
  nor (_39384_, _02057_, _38748_);
  or (_02058_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_02059_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_02060_, _01452_, _02059_);
  and (_02061_, _02060_, _43223_);
  and (_39421_, _02061_, _02058_);
  or (_02062_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_02063_, _01452_, _01660_);
  and (_02064_, _02063_, _43223_);
  and (_39422_, _02064_, _02062_);
  or (_02065_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_02066_, _01452_, _01655_);
  and (_02067_, _02066_, _43223_);
  and (_39423_, _02067_, _02065_);
  or (_02068_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_02069_, _01452_, _01649_);
  and (_02070_, _02069_, _43223_);
  and (_39424_, _02070_, _02068_);
  or (_02071_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_02072_, _01452_, _01644_);
  and (_02073_, _02072_, _43223_);
  and (_39425_, _02073_, _02071_);
  or (_02074_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_02075_, _01452_, _01635_);
  and (_02076_, _02075_, _43223_);
  and (_39427_, _02076_, _02074_);
  or (_02077_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_02078_, _01452_, _01625_);
  and (_02079_, _02078_, _43223_);
  and (_39428_, _02079_, _02077_);
  or (_02080_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_02081_, _01452_, _01620_);
  and (_02082_, _02081_, _43223_);
  and (_39429_, _02082_, _02080_);
  or (_02083_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_02084_, _01452_, _38904_);
  and (_02085_, _02084_, _43223_);
  and (_39430_, _02085_, _02083_);
  or (_02086_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_02087_, _01452_, _38910_);
  and (_02088_, _02087_, _43223_);
  and (_39431_, _02088_, _02086_);
  or (_02089_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_02090_, _01452_, _38915_);
  and (_02091_, _02090_, _43223_);
  and (_39432_, _02091_, _02089_);
  or (_02092_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_02093_, _01452_, _38900_);
  and (_02094_, _02093_, _43223_);
  and (_39433_, _02094_, _02092_);
  or (_02095_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_02096_, _01452_, _38921_);
  and (_02097_, _02096_, _43223_);
  and (_39434_, _02097_, _02095_);
  or (_02098_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_02099_, _01452_, _38896_);
  and (_02100_, _02099_, _43223_);
  and (_39435_, _02100_, _02098_);
  or (_02101_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_02102_, _01452_, _38892_);
  and (_02103_, _02102_, _43223_);
  and (_39436_, _02103_, _02101_);
  and (_02104_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_02105_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_02106_, _02105_, _02104_);
  and (_39441_, _02106_, _43223_);
  and (_02107_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_02108_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_02109_, _02108_, _02107_);
  and (_39442_, _02109_, _43223_);
  and (_02110_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_02111_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_02112_, _02111_, _02110_);
  and (_39443_, _02112_, _43223_);
  and (_02113_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_02114_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_02115_, _02114_, _02113_);
  and (_39444_, _02115_, _43223_);
  and (_02116_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_02117_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_02118_, _02117_, _02116_);
  and (_39445_, _02118_, _43223_);
  and (_02119_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_02120_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or (_02121_, _02120_, _02119_);
  and (_39446_, _02121_, _43223_);
  and (_02122_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_02123_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or (_02124_, _02123_, _02122_);
  and (_39447_, _02124_, _43223_);
  and (_02125_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_02126_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or (_02127_, _02126_, _02125_);
  and (_39448_, _02127_, _43223_);
  and (_02130_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_02132_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02134_, _02132_, _02130_);
  and (_39449_, _02134_, _43223_);
  and (_02137_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02139_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02141_, _02139_, _02137_);
  and (_39450_, _02141_, _43223_);
  and (_02144_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_02146_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02148_, _02146_, _02144_);
  and (_39452_, _02148_, _43223_);
  and (_02151_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_02153_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or (_02155_, _02153_, _02151_);
  and (_39453_, _02155_, _43223_);
  and (_02158_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_02160_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or (_02162_, _02160_, _02158_);
  and (_39454_, _02162_, _43223_);
  and (_02165_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_02167_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or (_02169_, _02167_, _02165_);
  and (_39455_, _02169_, _43223_);
  and (_02172_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_02174_, _01456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_02176_, _02174_, _02172_);
  and (_39456_, _02176_, _43223_);
  and (_39633_, _38504_, _43223_);
  and (_39634_, _38527_, _43223_);
  and (_39635_, _38548_, _43223_);
  nor (_39636_, _42664_, rst);
  and (_02183_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02185_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_02186_, _02185_, _02183_);
  and (_39637_, _02186_, _43223_);
  and (_02187_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02188_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02189_, _02188_, _02026_);
  or (_02190_, _02189_, _02187_);
  and (_39638_, _02190_, _43223_);
  and (_02191_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02192_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_02193_, _02192_, _02191_);
  and (_39639_, _02193_, _43223_);
  and (_02194_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02195_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_02196_, _02195_, _02194_);
  and (_39640_, _02196_, _43223_);
  and (_02197_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02198_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_02199_, _02198_, _02197_);
  and (_39642_, _02199_, _43223_);
  and (_02200_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02201_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_02202_, _02201_, _02026_);
  or (_02203_, _02202_, _02200_);
  and (_39643_, _02203_, _43223_);
  and (_02204_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02205_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_02206_, _02205_, _02026_);
  or (_02207_, _02206_, _02204_);
  and (_39644_, _02207_, _43223_);
  and (_02208_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02209_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_02210_, _02209_, _02208_);
  and (_39645_, _02210_, _43223_);
  and (_02211_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_02212_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_02213_, _02212_, _02211_);
  and (_39646_, _02213_, _43223_);
  and (_02214_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_02215_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_02216_, _02215_, _02214_);
  and (_39647_, _02216_, _43223_);
  and (_02217_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_02218_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_02219_, _02218_, _02217_);
  and (_39648_, _02219_, _43223_);
  and (_02220_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_02221_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_02222_, _02221_, _02220_);
  and (_39649_, _02222_, _43223_);
  and (_02223_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_02224_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_02225_, _02224_, _02223_);
  and (_39650_, _02225_, _43223_);
  and (_02226_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_02227_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_02228_, _02227_, _02226_);
  and (_39651_, _02228_, _43223_);
  and (_02229_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_02230_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_02231_, _02230_, _02229_);
  and (_39653_, _02231_, _43223_);
  and (_02232_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_02233_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_02234_, _02233_, _02232_);
  and (_39654_, _02234_, _43223_);
  and (_02235_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_02236_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_02237_, _02236_, _02235_);
  and (_39655_, _02237_, _43223_);
  and (_02238_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_02239_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_02240_, _02239_, _02238_);
  and (_39656_, _02240_, _43223_);
  and (_02241_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_02242_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_02243_, _02242_, _02241_);
  and (_39657_, _02243_, _43223_);
  and (_02244_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_02245_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_02246_, _02245_, _02244_);
  and (_39658_, _02246_, _43223_);
  and (_02247_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_02248_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_02249_, _02248_, _02247_);
  and (_39659_, _02249_, _43223_);
  and (_02250_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_02251_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_02252_, _02251_, _02250_);
  and (_39660_, _02252_, _43223_);
  and (_02253_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_02254_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_02255_, _02254_, _02253_);
  and (_39661_, _02255_, _43223_);
  and (_02256_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_02257_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_02258_, _02257_, _02256_);
  and (_39662_, _02258_, _43223_);
  and (_02259_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_02260_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_02261_, _02260_, _02259_);
  and (_39664_, _02261_, _43223_);
  and (_02262_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_02263_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_02264_, _02263_, _02262_);
  and (_39665_, _02264_, _43223_);
  and (_02265_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_02266_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_02267_, _02266_, _02265_);
  and (_39666_, _02267_, _43223_);
  and (_02268_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_02269_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_02270_, _02269_, _02268_);
  and (_39667_, _02270_, _43223_);
  and (_02271_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_02272_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_02273_, _02272_, _02271_);
  and (_39668_, _02273_, _43223_);
  and (_02274_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_02275_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_02276_, _02275_, _02274_);
  and (_39669_, _02276_, _43223_);
  and (_02277_, _02026_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_02278_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_02279_, _02278_, _02277_);
  and (_39670_, _02279_, _43223_);
  nor (_39671_, _42914_, rst);
  nor (_39673_, _42830_, rst);
  nor (_39674_, _43076_, rst);
  nor (_39675_, _42869_, rst);
  nor (_39676_, _42779_, rst);
  nor (_39677_, _43030_, rst);
  nor (_39679_, _42966_, rst);
  and (_39694_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _43223_);
  and (_39695_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _43223_);
  and (_39696_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _43223_);
  and (_39697_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _43223_);
  and (_39698_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _43223_);
  and (_39700_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _43223_);
  and (_39701_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _43223_);
  not (_02280_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_02281_, _01565_, _02280_);
  and (_02282_, _01668_, _01513_);
  or (_02283_, _01668_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02284_, _01669_);
  and (_02285_, _01716_, _02284_);
  and (_02286_, _02285_, _02283_);
  or (_02287_, _02286_, _02282_);
  or (_02288_, _01606_, _01568_);
  and (_02289_, _02288_, _32404_);
  or (_02290_, _02289_, _02287_);
  and (_02291_, _02290_, _01564_);
  or (_02292_, _02291_, _02281_);
  and (_39702_, _02292_, _43223_);
  and (_02293_, _02288_, _33101_);
  and (_02294_, _38710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_02295_, _01573_, _01366_);
  and (_02296_, _01661_, _01513_);
  or (_02297_, _02296_, _02295_);
  or (_02298_, _02297_, _02294_);
  or (_02299_, _01671_, _01669_);
  not (_02300_, _01672_);
  and (_02301_, _01716_, _02300_);
  and (_02302_, _02301_, _02299_);
  nor (_02303_, _02302_, _02298_);
  nand (_02304_, _02303_, _01564_);
  or (_02305_, _02304_, _02293_);
  or (_02306_, _01564_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_02307_, _02306_, _43223_);
  and (_39703_, _02307_, _02305_);
  and (_02308_, _02288_, _33819_);
  and (_02309_, _38710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02310_, _01573_, _01383_);
  and (_02311_, _01580_, _43056_);
  or (_02312_, _02311_, _02310_);
  or (_02313_, _02312_, _02309_);
  or (_02314_, _01676_, _01674_);
  not (_02315_, _01677_);
  and (_02316_, _01716_, _02315_);
  and (_02317_, _02316_, _02314_);
  nor (_02318_, _02317_, _02313_);
  nand (_02319_, _02318_, _01564_);
  or (_02320_, _02319_, _02308_);
  not (_02321_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02322_, _01722_, _02321_);
  and (_02323_, _01722_, _02321_);
  nor (_02324_, _02323_, _02322_);
  or (_02325_, _02324_, _01564_);
  and (_02326_, _02325_, _43223_);
  and (_39704_, _02326_, _02320_);
  and (_02327_, _02288_, _34602_);
  and (_02328_, _38710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02329_, _01573_, _01400_);
  and (_02330_, _01650_, _01513_);
  or (_02331_, _02330_, _02329_);
  or (_02332_, _02331_, _02328_);
  or (_02333_, _01654_, _01653_);
  or (_02334_, _02333_, _01678_);
  nand (_02335_, _02333_, _01678_);
  and (_02336_, _02335_, _01716_);
  and (_02337_, _02336_, _02334_);
  nor (_02338_, _02337_, _02332_);
  nand (_02339_, _02338_, _01564_);
  or (_02340_, _02339_, _02327_);
  and (_02341_, _02322_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02342_, _02322_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02343_, _02342_, _02341_);
  or (_02344_, _02343_, _01564_);
  and (_02345_, _02344_, _43223_);
  and (_39705_, _02345_, _02340_);
  and (_02347_, _02288_, _35288_);
  and (_02348_, _38710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02349_, _01573_, _01417_);
  and (_02350_, _01580_, _42754_);
  or (_02351_, _02350_, _02349_);
  or (_02352_, _02351_, _02348_);
  or (_02353_, _01682_, _01680_);
  and (_02354_, _01716_, _01683_);
  and (_02355_, _02354_, _02353_);
  nor (_02356_, _02355_, _02352_);
  nand (_02357_, _02356_, _01564_);
  or (_02358_, _02357_, _02347_);
  and (_02359_, _02341_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02360_, _02341_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02361_, _02360_, _02359_);
  or (_02362_, _02361_, _01564_);
  and (_02363_, _02362_, _43223_);
  and (_39706_, _02363_, _02358_);
  and (_02364_, _02288_, _36094_);
  and (_02365_, _38710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02366_, _01573_, _01434_);
  and (_02367_, _01637_, _01513_);
  or (_02368_, _02367_, _02366_);
  or (_02369_, _02368_, _02365_);
  or (_02370_, _01643_, _01641_);
  or (_02371_, _02370_, _01684_);
  nand (_02372_, _02370_, _01684_);
  and (_02373_, _02372_, _01716_);
  and (_02374_, _02373_, _02371_);
  nor (_02375_, _02374_, _02369_);
  nand (_02376_, _02375_, _01564_);
  or (_02377_, _02376_, _02364_);
  nor (_02378_, _02359_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02379_, _02378_, _01727_);
  or (_02380_, _02379_, _01564_);
  and (_02381_, _02380_, _43223_);
  and (_39707_, _02381_, _02377_);
  nor (_02382_, _01727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02383_, _01727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02384_, _02383_, _02382_);
  or (_02385_, _02384_, _01564_);
  and (_02386_, _02385_, _43223_);
  and (_02387_, _02288_, _36822_);
  and (_02388_, _38710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02389_, _01573_, _01451_);
  and (_02390_, _01626_, _01513_);
  or (_02391_, _02390_, _02389_);
  or (_02392_, _02391_, _02388_);
  or (_02393_, _01686_, _01634_);
  not (_02394_, _01687_);
  and (_02395_, _01716_, _02394_);
  and (_02396_, _02395_, _02393_);
  nor (_02397_, _02396_, _02392_);
  nand (_02398_, _02397_, _01564_);
  or (_02399_, _02398_, _02387_);
  and (_39708_, _02399_, _02386_);
  and (_02400_, _02288_, _31195_);
  or (_02401_, _01622_, _01623_);
  nand (_02402_, _02401_, _01688_);
  and (_02403_, _01603_, _01711_);
  or (_02404_, _02401_, _01688_);
  and (_02405_, _02404_, _02403_);
  and (_02406_, _02405_, _02402_);
  nor (_02407_, _01573_, _01332_);
  and (_02408_, _01580_, _42659_);
  and (_02409_, _38710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_02410_, _02409_, _02408_);
  nor (_02411_, _02410_, _02407_);
  nand (_02412_, _02411_, _01564_);
  or (_02413_, _02412_, _02406_);
  or (_02414_, _02413_, _02400_);
  nor (_02415_, _02383_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02416_, _02383_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_02417_, _02416_, _02415_);
  or (_02418_, _02417_, _01564_);
  and (_02419_, _02418_, _43223_);
  and (_39709_, _02419_, _02414_);
  not (_02420_, _01564_);
  nor (_02421_, _01460_, _32393_);
  not (_02422_, _39012_);
  and (_02423_, _01568_, _02422_);
  and (_02424_, _01572_, _42933_);
  and (_02425_, _01580_, _00785_);
  and (_02426_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_02427_, _02426_, _02425_);
  or (_02428_, _02427_, _02424_);
  and (_02429_, _01690_, _38904_);
  nor (_02430_, _01690_, _38904_);
  nor (_02431_, _02430_, _02429_);
  nor (_02432_, _02431_, _01619_);
  and (_02433_, _02431_, _01619_);
  or (_02434_, _02433_, _02432_);
  and (_02435_, _02434_, _02403_);
  or (_02436_, _02435_, _02428_);
  or (_02437_, _02436_, _02423_);
  or (_02438_, _02437_, _02421_);
  or (_02439_, _02438_, _02420_);
  or (_02440_, _02416_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_02441_, _01729_, _01727_);
  and (_02442_, _02441_, _02440_);
  or (_02443_, _02442_, _01564_);
  and (_02444_, _02443_, _43223_);
  and (_39711_, _02444_, _02439_);
  nor (_02445_, _01460_, _33090_);
  and (_02446_, _01690_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02447_, _02446_, _01617_);
  and (_02448_, _01696_, _01619_);
  nor (_02449_, _02448_, _02447_);
  nor (_02450_, _02449_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_02451_, _02449_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_02452_, _02451_, _02450_);
  and (_02453_, _02452_, _02403_);
  not (_02454_, _39045_);
  and (_02455_, _01568_, _02454_);
  and (_02456_, _01580_, _00773_);
  and (_02457_, _01572_, _42808_);
  or (_02458_, _02457_, _02456_);
  and (_02459_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_02460_, _02459_, _02458_);
  nor (_02461_, _02460_, _02455_);
  nand (_02462_, _02461_, _01564_);
  or (_02463_, _02462_, _02453_);
  or (_02464_, _02463_, _02445_);
  nand (_02465_, _02441_, _01764_);
  or (_02466_, _02441_, _01764_);
  and (_02467_, _02466_, _02465_);
  or (_02468_, _02467_, _01564_);
  and (_02469_, _02468_, _43223_);
  and (_39712_, _02469_, _02464_);
  nor (_02470_, _01460_, _33809_);
  not (_02471_, _39076_);
  and (_02472_, _01568_, _02471_);
  and (_02473_, _01572_, _43056_);
  and (_02474_, _01580_, _00763_);
  and (_02475_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_02476_, _02475_, _02474_);
  or (_02477_, _02476_, _02473_);
  or (_02478_, _02477_, _02472_);
  and (_02479_, _01697_, _01619_);
  and (_02480_, _02447_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02481_, _02480_, _02479_);
  nor (_02482_, _02481_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_02483_, _02481_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_02484_, _02483_, _02482_);
  and (_02485_, _02484_, _02403_);
  or (_02486_, _02485_, _02478_);
  or (_02487_, _02486_, _02470_);
  or (_02488_, _02487_, _02420_);
  nor (_02489_, _01731_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_02490_, _02489_, _01732_);
  or (_02491_, _02490_, _01564_);
  and (_02492_, _02491_, _43223_);
  and (_39713_, _02492_, _02488_);
  nor (_02493_, _01460_, _34591_);
  and (_02494_, _01691_, _01617_);
  and (_02495_, _01698_, _01619_);
  nor (_02496_, _02495_, _02494_);
  nor (_02497_, _02496_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02498_, _02496_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_02499_, _02498_, _02497_);
  and (_02500_, _02499_, _02403_);
  not (_02501_, _39108_);
  and (_02502_, _01568_, _02501_);
  and (_02503_, _01572_, _42889_);
  nor (_02504_, _01589_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02505_, _02504_, _01590_);
  and (_02506_, _02505_, _01580_);
  and (_02507_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_02508_, _02507_, _02506_);
  or (_02509_, _02508_, _02503_);
  nor (_02510_, _02509_, _02502_);
  nand (_02511_, _02510_, _01564_);
  or (_02512_, _02511_, _02500_);
  or (_02513_, _02512_, _02493_);
  nor (_02514_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02515_, _02514_, _01733_);
  or (_02516_, _02515_, _01564_);
  and (_02517_, _02516_, _43223_);
  and (_39714_, _02517_, _02513_);
  nor (_02518_, _01460_, _35277_);
  and (_02519_, _01692_, _01617_);
  and (_02520_, _01699_, _01619_);
  nor (_02521_, _02520_, _02519_);
  nor (_02522_, _02521_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02523_, _02521_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_02524_, _02523_, _02522_);
  and (_02525_, _02524_, _02403_);
  not (_02526_, _39139_);
  and (_02527_, _01568_, _02526_);
  and (_02528_, _01572_, _42754_);
  nor (_02529_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02530_, _02529_, _01591_);
  and (_02531_, _02530_, _01580_);
  and (_02532_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_02533_, _02532_, _02531_);
  or (_02534_, _02533_, _02528_);
  nor (_02535_, _02534_, _02527_);
  nand (_02536_, _02535_, _01564_);
  or (_02537_, _02536_, _02525_);
  or (_02539_, _02537_, _02518_);
  nor (_02540_, _01733_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02541_, _02540_, _01734_);
  or (_02542_, _02541_, _01564_);
  and (_02543_, _02542_, _43223_);
  and (_39715_, _02543_, _02539_);
  and (_02544_, _01693_, _01617_);
  and (_02545_, _01700_, _01619_);
  nor (_02546_, _02545_, _02544_);
  nand (_02547_, _02546_, _38896_);
  or (_02548_, _02546_, _38896_);
  and (_02549_, _02548_, _02403_);
  and (_02550_, _02549_, _02547_);
  not (_02551_, _39173_);
  and (_02552_, _01568_, _02551_);
  and (_02553_, _01572_, _43010_);
  and (_02554_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_02555_, _02554_, _02553_);
  nor (_02556_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_02557_, _02556_, _01592_);
  and (_02558_, _02557_, _01580_);
  or (_02559_, _02558_, _02555_);
  or (_02561_, _02559_, _02552_);
  or (_02562_, _02561_, _02550_);
  nor (_02563_, _01460_, _36083_);
  or (_02564_, _02563_, _02420_);
  or (_02565_, _02564_, _02562_);
  nor (_02566_, _01734_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_02567_, _02566_, _01735_);
  or (_02568_, _02567_, _01564_);
  and (_02569_, _02568_, _43223_);
  and (_39716_, _02569_, _02565_);
  nor (_02570_, _01460_, _36811_);
  nor (_02572_, _01703_, _38892_);
  and (_02573_, _01703_, _38892_);
  or (_02574_, _02573_, _02572_);
  and (_02575_, _02574_, _02403_);
  not (_02576_, _39203_);
  and (_02577_, _01568_, _02576_);
  or (_02578_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02579_, _02578_, _01593_);
  and (_02580_, _02579_, _01580_);
  and (_02581_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_02582_, _01572_, _42986_);
  or (_02583_, _02582_, _02581_);
  or (_02584_, _02583_, _02580_);
  or (_02585_, _02584_, _02577_);
  or (_02586_, _02585_, _02575_);
  or (_02587_, _02586_, _02570_);
  or (_02588_, _02587_, _02420_);
  nor (_02589_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02590_, _02589_, _01736_);
  or (_02591_, _02590_, _01564_);
  and (_02592_, _02591_, _43223_);
  and (_39717_, _02592_, _02588_);
  and (_02593_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_02594_, _01928_, _01926_);
  nor (_02595_, _02594_, _01929_);
  or (_02596_, _02595_, _01746_);
  or (_02597_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02598_, _02597_, _01960_);
  and (_02599_, _02598_, _02596_);
  or (_39718_, _02599_, _02593_);
  or (_02600_, _01931_, _01929_);
  and (_02601_, _02600_, _01932_);
  or (_02602_, _02601_, _01746_);
  or (_02603_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02604_, _02603_, _01960_);
  and (_02605_, _02604_, _02602_);
  and (_02606_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39719_, _02606_, _02605_);
  and (_02607_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02608_, _01936_, _01934_);
  nor (_02609_, _02608_, _01937_);
  or (_02610_, _02609_, _01746_);
  or (_02611_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_02612_, _02611_, _01960_);
  and (_02613_, _02612_, _02610_);
  or (_39720_, _02613_, _02607_);
  nor (_02614_, _01937_, _01822_);
  nor (_02615_, _02614_, _01938_);
  or (_02616_, _02615_, _01746_);
  or (_02617_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_02618_, _02617_, _01960_);
  and (_02619_, _02618_, _02616_);
  and (_02620_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_39722_, _02620_, _02619_);
  and (_02621_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02622_, _01941_, _01938_);
  nor (_02623_, _02622_, _01942_);
  or (_02624_, _02623_, _01746_);
  or (_02625_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_02626_, _02625_, _01960_);
  and (_02627_, _02626_, _02624_);
  or (_39723_, _02627_, _02621_);
  and (_02628_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02629_, _01942_, _01817_);
  nor (_02630_, _02629_, _01943_);
  or (_02631_, _02630_, _01746_);
  or (_02632_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_02633_, _02632_, _01960_);
  and (_02634_, _02633_, _02631_);
  or (_39724_, _02634_, _02628_);
  nor (_02635_, _01943_, _01813_);
  nor (_02636_, _02635_, _01944_);
  or (_02637_, _02636_, _01746_);
  or (_02638_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02639_, _02638_, _01960_);
  and (_02640_, _02639_, _02637_);
  and (_02641_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39725_, _02641_, _02640_);
  or (_02642_, _01944_, _01809_);
  nor (_02643_, _01945_, _01746_);
  and (_02644_, _02643_, _02642_);
  nor (_02645_, _01745_, _01620_);
  or (_02646_, _02645_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02647_, _02646_, _02644_);
  or (_02648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _37050_);
  and (_02649_, _02648_, _43223_);
  and (_39726_, _02649_, _02647_);
  or (_02650_, _01947_, _01945_);
  nor (_02651_, _01948_, _01746_);
  and (_02652_, _02651_, _02650_);
  nor (_02653_, _01745_, _38904_);
  or (_02654_, _02653_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02655_, _02654_, _02652_);
  or (_02656_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _37050_);
  and (_02657_, _02656_, _43223_);
  and (_39727_, _02657_, _02655_);
  nor (_02658_, _01948_, _01805_);
  nor (_02659_, _02658_, _01949_);
  or (_02660_, _02659_, _01746_);
  or (_02661_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_02662_, _02661_, _01960_);
  and (_02663_, _02662_, _02660_);
  and (_02664_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39728_, _02664_, _02663_);
  nor (_02665_, _01949_, _01801_);
  nor (_02666_, _02665_, _01950_);
  or (_02667_, _02666_, _01746_);
  or (_02668_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_02669_, _02668_, _01960_);
  and (_02670_, _02669_, _02667_);
  and (_02671_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_39729_, _02671_, _02670_);
  nor (_02672_, _01950_, _01798_);
  nor (_02673_, _02672_, _01951_);
  or (_02674_, _02673_, _01746_);
  or (_02675_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02676_, _02675_, _01960_);
  and (_02677_, _02676_, _02674_);
  and (_02678_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39730_, _02678_, _02677_);
  nor (_02679_, _01951_, _01793_);
  nor (_02680_, _02679_, _01952_);
  or (_02681_, _02680_, _01746_);
  or (_02682_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02683_, _02682_, _01960_);
  and (_02684_, _02683_, _02681_);
  and (_02685_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39731_, _02685_, _02684_);
  nor (_02686_, _01952_, _01789_);
  nor (_02687_, _02686_, _01953_);
  or (_02688_, _02687_, _01746_);
  or (_02689_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_02690_, _02689_, _01960_);
  and (_02691_, _02690_, _02688_);
  and (_02692_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39733_, _02692_, _02691_);
  nor (_02693_, _01953_, _01786_);
  nor (_02694_, _02693_, _01954_);
  or (_02695_, _02694_, _01746_);
  or (_02696_, _01745_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02697_, _02696_, _01960_);
  and (_02698_, _02697_, _02695_);
  and (_02699_, _01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_39734_, _02699_, _02698_);
  and (_02700_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_02701_, _02700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39735_, _02701_, _43223_);
  and (_02702_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_02703_, _02702_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39736_, _02703_, _43223_);
  and (_02704_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_02705_, _02704_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39737_, _02705_, _43223_);
  and (_02706_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_02707_, _02706_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39738_, _02707_, _43223_);
  and (_02708_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_02709_, _02708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39739_, _02709_, _43223_);
  and (_02710_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_02711_, _02710_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39740_, _02711_, _43223_);
  and (_02712_, _01970_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_02713_, _02712_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39741_, _02713_, _43223_);
  nor (_02714_, _01925_, _42642_);
  nand (_02715_, _02714_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_02717_, _02714_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_02718_, _02717_, _01960_);
  and (_39742_, _02718_, _02715_);
  or (_02719_, _01982_, _01980_);
  and (_02720_, _02719_, _01983_);
  or (_02721_, _02720_, _42642_);
  or (_02722_, _37083_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_02723_, _02722_, _01960_);
  and (_39744_, _02723_, _02721_);
  and (_02724_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_02725_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_02726_, _02725_, _39370_);
  or (_39760_, _02726_, _02724_);
  and (_02727_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_02728_, _02188_, _39370_);
  or (_39761_, _02728_, _02727_);
  and (_02729_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_02730_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_02731_, _02730_, _39370_);
  or (_39762_, _02731_, _02729_);
  and (_02732_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_02733_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_02734_, _02733_, _39370_);
  or (_39763_, _02734_, _02732_);
  and (_02735_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_02736_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_02737_, _02736_, _39370_);
  or (_39764_, _02737_, _02735_);
  and (_02738_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_02739_, _02201_, _39370_);
  or (_39766_, _02739_, _02738_);
  and (_02740_, _02004_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_02741_, _02205_, _39370_);
  or (_39767_, _02741_, _02740_);
  and (_39768_, _02012_, _43223_);
  nor (_39769_, _02022_, rst);
  and (_39770_, _02018_, _43223_);
  and (_02742_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02743_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_02744_, _02743_, _02742_);
  and (_39771_, _02744_, _43223_);
  and (_02745_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02746_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_02747_, _02746_, _02745_);
  and (_39772_, _02747_, _43223_);
  and (_02748_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02749_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_02750_, _02749_, _02748_);
  and (_39773_, _02750_, _43223_);
  and (_02751_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02752_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_02753_, _02752_, _02751_);
  and (_39774_, _02753_, _43223_);
  and (_02754_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02755_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_02756_, _02755_, _02754_);
  and (_39775_, _02756_, _43223_);
  and (_02757_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02758_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_02759_, _02758_, _02757_);
  and (_39777_, _02759_, _43223_);
  and (_02760_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02761_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_02762_, _02761_, _02760_);
  and (_39778_, _02762_, _43223_);
  and (_02763_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02764_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_02765_, _02764_, _02763_);
  and (_39779_, _02765_, _43223_);
  and (_02766_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_02767_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_02768_, _02767_, _02766_);
  and (_39780_, _02768_, _43223_);
  and (_02769_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_02770_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_02771_, _02770_, _02769_);
  and (_39781_, _02771_, _43223_);
  and (_02772_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_02773_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_02774_, _02773_, _02772_);
  and (_39782_, _02774_, _43223_);
  and (_02775_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_02776_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_02777_, _02776_, _02775_);
  and (_39783_, _02777_, _43223_);
  and (_02778_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_02779_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_02780_, _02779_, _02778_);
  and (_39784_, _02780_, _43223_);
  and (_02781_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_02782_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_02783_, _02782_, _02781_);
  and (_39785_, _02783_, _43223_);
  and (_02784_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_02785_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_02786_, _02785_, _02784_);
  and (_39786_, _02786_, _43223_);
  and (_02787_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_02788_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_02789_, _02788_, _02787_);
  and (_39788_, _02789_, _43223_);
  and (_02790_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_02791_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_02792_, _02791_, _02790_);
  and (_39789_, _02792_, _43223_);
  and (_02793_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_02794_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_02795_, _02794_, _02793_);
  and (_39790_, _02795_, _43223_);
  and (_02796_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_02797_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_02798_, _02797_, _02796_);
  and (_39791_, _02798_, _43223_);
  and (_02799_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_02800_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_02801_, _02800_, _02799_);
  and (_39792_, _02801_, _43223_);
  and (_02802_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02803_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_02804_, _02803_, _02802_);
  and (_39793_, _02804_, _43223_);
  and (_02805_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02807_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_02808_, _02807_, _02805_);
  and (_39794_, _02808_, _43223_);
  and (_02809_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_02810_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_02812_, _02810_, _02809_);
  and (_39795_, _02812_, _43223_);
  and (_02813_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_02814_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_02815_, _02814_, _02813_);
  and (_39796_, _02815_, _43223_);
  and (_02817_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_02818_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_02819_, _02818_, _02817_);
  and (_39797_, _02819_, _43223_);
  and (_02821_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_02822_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_02823_, _02822_, _02821_);
  and (_39799_, _02823_, _43223_);
  and (_02824_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_02826_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_02827_, _02826_, _02824_);
  and (_39800_, _02827_, _43223_);
  and (_02828_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_02829_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_02831_, _02829_, _02828_);
  and (_39801_, _02831_, _43223_);
  and (_02832_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_02833_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_02834_, _02833_, _02832_);
  and (_39802_, _02834_, _43223_);
  and (_02836_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_02838_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_02839_, _02838_, _02836_);
  and (_39803_, _02839_, _43223_);
  and (_02840_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_02841_, _02028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_02842_, _02841_, _02840_);
  and (_39804_, _02842_, _43223_);
  and (_02845_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02846_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_02847_, _02846_, _02845_);
  and (_39805_, _02847_, _43223_);
  and (_02849_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02850_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_02852_, _02850_, _02849_);
  and (_39806_, _02852_, _43223_);
  and (_02853_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02856_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_02857_, _02856_, _02853_);
  and (_39807_, _02857_, _43223_);
  and (_02859_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02860_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_02861_, _02860_, _02859_);
  and (_39808_, _02861_, _43223_);
  and (_02863_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02864_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_02866_, _02864_, _02863_);
  and (_39810_, _02866_, _43223_);
  and (_02868_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02869_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_02870_, _02869_, _02868_);
  and (_39811_, _02870_, _43223_);
  and (_02871_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02872_, _02036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_02873_, _02872_, _02871_);
  and (_39812_, _02873_, _43223_);
  and (_02875_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02877_, _42914_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02879_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_02880_, _02879_, _02035_);
  and (_02881_, _02880_, _02877_);
  or (_02883_, _02881_, _02875_);
  and (_39813_, _02883_, _43223_);
  and (_02884_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02886_, _42830_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02887_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_02888_, _02887_, _02035_);
  and (_02891_, _02888_, _02886_);
  or (_02892_, _02891_, _02884_);
  and (_39814_, _02892_, _43223_);
  and (_02894_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02895_, _43076_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02896_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_02898_, _02896_, _02035_);
  and (_02899_, _02898_, _02895_);
  or (_02901_, _02899_, _02894_);
  and (_39815_, _02901_, _43223_);
  and (_02903_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02904_, _42869_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02905_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_02907_, _02905_, _02035_);
  and (_02908_, _02907_, _02904_);
  or (_02909_, _02908_, _02903_);
  and (_39816_, _02909_, _43223_);
  and (_02911_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02912_, _42779_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02914_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_02915_, _02914_, _02035_);
  and (_02916_, _02915_, _02912_);
  or (_02918_, _02916_, _02911_);
  and (_39817_, _02918_, _43223_);
  and (_02919_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02921_, _43030_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02922_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_02923_, _02922_, _02035_);
  and (_02925_, _02923_, _02921_);
  or (_02926_, _02925_, _02919_);
  and (_39818_, _02926_, _43223_);
  and (_02929_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02930_, _42966_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02932_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02933_, _02932_, _02035_);
  and (_02934_, _02933_, _02930_);
  or (_02935_, _02934_, _02929_);
  and (_39819_, _02935_, _43223_);
  and (_02936_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02937_, _42716_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02940_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_02941_, _02940_, _02035_);
  and (_02942_, _02941_, _02937_);
  or (_02944_, _02942_, _02936_);
  and (_39821_, _02944_, _43223_);
  and (_02945_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_02947_, _02945_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02948_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _02035_);
  and (_02949_, _02948_, _43223_);
  and (_39822_, _02949_, _02947_);
  and (_02952_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_02953_, _02952_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02955_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _02035_);
  and (_02956_, _02955_, _43223_);
  and (_39823_, _02956_, _02953_);
  and (_02958_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_02959_, _02958_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02960_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _02035_);
  and (_02962_, _02960_, _43223_);
  and (_39824_, _02962_, _02959_);
  and (_02965_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_02966_, _02965_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02967_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _02035_);
  and (_02968_, _02967_, _43223_);
  and (_39825_, _02968_, _02966_);
  and (_02970_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_02971_, _02970_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02973_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _02035_);
  and (_02974_, _02973_, _43223_);
  and (_39826_, _02974_, _02971_);
  and (_02977_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_02978_, _02977_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02979_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _02035_);
  and (_02981_, _02979_, _43223_);
  and (_39827_, _02981_, _02978_);
  and (_02982_, _02042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_02984_, _02982_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02985_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _02035_);
  and (_02986_, _02985_, _43223_);
  and (_39828_, _02986_, _02984_);
  nand (_02989_, _02049_, _32393_);
  or (_02990_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02992_, _02990_, _43223_);
  and (_39829_, _02992_, _02989_);
  nand (_02994_, _02049_, _33090_);
  or (_02995_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02996_, _02995_, _43223_);
  and (_39830_, _02996_, _02994_);
  nand (_02998_, _02049_, _33809_);
  or (_02999_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_03001_, _02999_, _43223_);
  and (_39832_, _03001_, _02998_);
  nand (_03003_, _02049_, _34591_);
  or (_03004_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_03006_, _03004_, _43223_);
  and (_39833_, _03006_, _03003_);
  nand (_03007_, _02049_, _35277_);
  or (_03009_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_03010_, _03009_, _43223_);
  and (_39834_, _03010_, _03007_);
  nand (_03013_, _02049_, _36083_);
  or (_03014_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_03015_, _03014_, _43223_);
  and (_39835_, _03015_, _03013_);
  nand (_03017_, _02049_, _36811_);
  or (_03018_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_03020_, _03018_, _43223_);
  and (_39836_, _03020_, _03017_);
  nand (_03022_, _02049_, _31194_);
  or (_03023_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_03025_, _03023_, _43223_);
  and (_39837_, _03025_, _03022_);
  nand (_03027_, _02049_, _39012_);
  or (_03028_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_03029_, _03028_, _43223_);
  and (_39838_, _03029_, _03027_);
  nand (_03031_, _02049_, _39045_);
  or (_03032_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_03034_, _03032_, _43223_);
  and (_39839_, _03034_, _03031_);
  nand (_03035_, _02049_, _39076_);
  or (_03037_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_03038_, _03037_, _43223_);
  and (_39840_, _03038_, _03035_);
  nand (_03040_, _02049_, _39108_);
  or (_03041_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_03042_, _03041_, _43223_);
  and (_39841_, _03042_, _03040_);
  nand (_03044_, _02049_, _39139_);
  or (_03045_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_03047_, _03045_, _43223_);
  and (_39843_, _03047_, _03044_);
  nand (_03049_, _02049_, _39173_);
  or (_03050_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_03051_, _03050_, _43223_);
  and (_39844_, _03051_, _03049_);
  nand (_03052_, _02049_, _39203_);
  or (_03053_, _02049_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_03054_, _03053_, _43223_);
  and (_39845_, _03054_, _03052_);
  nor (_40063_, _42736_, rst);
  and (_03056_, _42672_, _38753_);
  and (_03058_, _03056_, _39409_);
  and (_03059_, _03058_, _42674_);
  nand (_03060_, _03059_, _38837_);
  or (_03062_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_03063_, _03062_, _43223_);
  and (_40064_, _03063_, _03060_);
  and (_03065_, _03056_, _39699_);
  not (_03066_, _03065_);
  nor (_03067_, _03066_, _38837_);
  not (_03069_, _42674_);
  and (_03070_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03071_, _03070_, _03069_);
  or (_03073_, _03071_, _03067_);
  or (_03074_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03075_, _03074_, _43223_);
  and (_40065_, _03075_, _03073_);
  and (_03077_, _27624_, _28293_);
  and (_03079_, _03056_, _03077_);
  and (_03080_, _03079_, _42674_);
  nand (_03081_, _03080_, _38837_);
  or (_03082_, _03080_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_03084_, _03082_, _43223_);
  and (_40066_, _03084_, _03081_);
  and (_03085_, _03056_, _41781_);
  and (_03087_, _03085_, _42674_);
  not (_03088_, _03087_);
  nor (_03089_, _03088_, _38837_);
  and (_03091_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_03092_, _03091_, _03089_);
  and (_40068_, _03092_, _43223_);
  and (_03094_, _42672_, _39235_);
  and (_03095_, _03094_, _39409_);
  and (_03096_, _03095_, _42674_);
  not (_03098_, _03096_);
  and (_03099_, _03098_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_03100_, _03098_, _38837_);
  or (_03102_, _03100_, _03099_);
  and (_40069_, _03102_, _43223_);
  or (_03103_, _03085_, _03079_);
  or (_03105_, _03095_, _03103_);
  and (_03106_, _03105_, _42674_);
  not (_03108_, _03079_);
  nor (_03109_, _03095_, _03085_);
  and (_03110_, _03094_, _39699_);
  not (_03111_, _03110_);
  and (_03113_, _03111_, _03109_);
  and (_03114_, _03113_, _03108_);
  nor (_03115_, _03065_, _03058_);
  nand (_03117_, _03115_, _42674_);
  or (_03118_, _03117_, _03114_);
  or (_03119_, _03118_, _03106_);
  and (_03121_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_03122_, _03110_, _42674_);
  and (_03123_, _03122_, _42714_);
  or (_03125_, _03123_, _03121_);
  and (_40070_, _03125_, _43223_);
  and (_03126_, _03094_, _03077_);
  and (_03128_, _03126_, _42714_);
  not (_03130_, _03113_);
  nor (_03131_, _03126_, _03110_);
  and (_03133_, _03131_, _03109_);
  and (_03134_, _03108_, _03115_);
  nand (_03135_, _03134_, _42674_);
  or (_03137_, _03135_, _03133_);
  or (_03138_, _03137_, _03130_);
  and (_03140_, _03138_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_03141_, _03140_, _03128_);
  or (_03142_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_03143_, _03142_, _43223_);
  and (_40071_, _03143_, _03141_);
  and (_03145_, _03094_, _41781_);
  and (_03146_, _03145_, _42674_);
  not (_03148_, _03146_);
  nor (_03149_, _03148_, _38837_);
  not (_03150_, _03095_);
  and (_03152_, _03131_, _03150_);
  not (_03153_, _03152_);
  nor (_03154_, _03153_, _03145_);
  not (_03156_, _03085_);
  and (_03157_, _03156_, _03134_);
  nand (_03158_, _03157_, _42674_);
  or (_03160_, _03158_, _03154_);
  or (_03161_, _03160_, _03153_);
  and (_03162_, _03161_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_03164_, _03162_, _03149_);
  and (_40072_, _03164_, _43223_);
  nand (_03165_, _03059_, _38816_);
  or (_03167_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03168_, _03167_, _43223_);
  and (_40162_, _03168_, _03165_);
  nand (_03170_, _03059_, _38808_);
  or (_03171_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03172_, _03171_, _43223_);
  and (_40163_, _03172_, _03170_);
  nand (_03174_, _03059_, _38801_);
  or (_03175_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_03176_, _03175_, _43223_);
  and (_40164_, _03176_, _03174_);
  nand (_03178_, _03059_, _38793_);
  or (_03179_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_03181_, _03179_, _43223_);
  and (_40165_, _03181_, _03178_);
  nand (_03182_, _03059_, _38786_);
  or (_03184_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_03185_, _03184_, _43223_);
  and (_40166_, _03185_, _03182_);
  nand (_03187_, _03059_, _38778_);
  or (_03188_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03189_, _03188_, _43223_);
  and (_40167_, _03189_, _03187_);
  nand (_03191_, _03059_, _38770_);
  or (_03192_, _03059_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03194_, _03192_, _43223_);
  and (_40168_, _03194_, _03191_);
  and (_03196_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_03197_, _03065_, _38817_);
  or (_03198_, _03197_, _03069_);
  or (_03199_, _03198_, _03196_);
  or (_03201_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_03202_, _03201_, _43223_);
  and (_40169_, _03202_, _03199_);
  nor (_03204_, _03066_, _38808_);
  and (_03205_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_03206_, _03205_, _03069_);
  or (_03208_, _03206_, _03204_);
  or (_03209_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03210_, _03209_, _43223_);
  and (_40170_, _03210_, _03208_);
  nor (_03212_, _03066_, _38801_);
  and (_03213_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03215_, _03213_, _03069_);
  or (_03216_, _03215_, _03212_);
  or (_03217_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03219_, _03217_, _43223_);
  and (_40171_, _03219_, _03216_);
  nor (_03220_, _03066_, _38793_);
  and (_03222_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03223_, _03222_, _03069_);
  or (_03225_, _03223_, _03220_);
  or (_03226_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03227_, _03226_, _43223_);
  and (_40173_, _03227_, _03225_);
  nor (_03229_, _03066_, _38786_);
  and (_03230_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_03231_, _03230_, _03069_);
  or (_03233_, _03231_, _03229_);
  or (_03234_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_03235_, _03234_, _43223_);
  and (_40174_, _03235_, _03233_);
  nor (_03237_, _03066_, _38778_);
  and (_03238_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_03240_, _03238_, _03069_);
  or (_03241_, _03240_, _03237_);
  or (_03242_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_03244_, _03242_, _43223_);
  and (_40175_, _03244_, _03241_);
  nor (_03245_, _03066_, _38770_);
  and (_03247_, _03066_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03248_, _03247_, _03069_);
  or (_03249_, _03248_, _03245_);
  or (_03251_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03252_, _03251_, _43223_);
  and (_40176_, _03252_, _03249_);
  nand (_03254_, _03080_, _38816_);
  or (_03255_, _03080_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_03256_, _03255_, _03254_);
  and (_40177_, _03256_, _43223_);
  not (_03258_, _03080_);
  nor (_03259_, _03258_, _38808_);
  and (_03261_, _03258_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_03262_, _03261_, _03259_);
  and (_40178_, _03262_, _43223_);
  nor (_03264_, _03258_, _38801_);
  and (_03265_, _03258_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_03266_, _03265_, _03264_);
  and (_40179_, _03266_, _43223_);
  nor (_03268_, _03258_, _38793_);
  and (_03269_, _03258_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_03271_, _03269_, _03268_);
  and (_40180_, _03271_, _43223_);
  nand (_03272_, _03080_, _38786_);
  or (_03274_, _03080_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_03275_, _03274_, _43223_);
  and (_40181_, _03275_, _03272_);
  nor (_03277_, _03258_, _38778_);
  and (_03278_, _03258_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_03279_, _03278_, _03277_);
  and (_40182_, _03279_, _43223_);
  nor (_03280_, _03258_, _38770_);
  and (_03281_, _03258_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_03282_, _03281_, _03280_);
  and (_40184_, _03282_, _43223_);
  and (_03283_, _03087_, _38817_);
  and (_03284_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_03285_, _03284_, _03283_);
  and (_40185_, _03285_, _43223_);
  and (_03286_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_03287_, _03088_, _38808_);
  or (_03288_, _03287_, _03286_);
  and (_40186_, _03288_, _43223_);
  nor (_03289_, _03088_, _38801_);
  and (_03290_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_03291_, _03290_, _03289_);
  and (_40187_, _03291_, _43223_);
  nor (_03292_, _03088_, _38793_);
  and (_03293_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_03294_, _03293_, _03292_);
  and (_40188_, _03294_, _43223_);
  and (_03295_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_03296_, _03088_, _38786_);
  or (_03297_, _03296_, _03295_);
  and (_40189_, _03297_, _43223_);
  nor (_03298_, _03088_, _38778_);
  and (_03299_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_03300_, _03299_, _03298_);
  and (_40190_, _03300_, _43223_);
  nor (_03301_, _03088_, _38770_);
  and (_03302_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03303_, _03302_, _03301_);
  and (_40191_, _03303_, _43223_);
  and (_03304_, _03098_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_03305_, _03096_, _38817_);
  or (_03306_, _03305_, _03304_);
  and (_40192_, _03306_, _43223_);
  and (_03307_, _03098_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_03308_, _03098_, _38808_);
  or (_03309_, _03308_, _03307_);
  and (_40193_, _03309_, _43223_);
  nor (_03310_, _03098_, _38801_);
  and (_03311_, _03109_, _03134_);
  or (_03312_, _03311_, _03069_);
  or (_03313_, _03103_, _03065_);
  and (_03314_, _03313_, _42674_);
  or (_03315_, _03314_, _03058_);
  or (_03316_, _03315_, _03312_);
  and (_03317_, _03316_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_03318_, _03317_, _03310_);
  and (_40195_, _03318_, _43223_);
  nor (_03319_, _03098_, _38793_);
  and (_03320_, _03316_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_03321_, _03320_, _03319_);
  and (_40196_, _03321_, _43223_);
  nor (_03322_, _03098_, _38786_);
  not (_03323_, _03157_);
  or (_03324_, _03312_, _03323_);
  and (_03325_, _03324_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or (_03326_, _03325_, _03322_);
  and (_40197_, _03326_, _43223_);
  nor (_03327_, _03098_, _38778_);
  and (_03328_, _03324_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_03329_, _03328_, _03327_);
  and (_40198_, _03329_, _43223_);
  nor (_03330_, _03098_, _38770_);
  and (_03331_, _03316_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_03332_, _03331_, _03330_);
  and (_40199_, _03332_, _43223_);
  and (_03333_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_03334_, _03069_, _38816_);
  and (_03336_, _03334_, _03110_);
  or (_03337_, _03336_, _03333_);
  and (_40200_, _03337_, _43223_);
  and (_03338_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_03339_, _03122_, _42828_);
  or (_03340_, _03339_, _03338_);
  and (_40201_, _03340_, _43223_);
  and (_03341_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_03342_, _03122_, _43074_);
  or (_03343_, _03342_, _03341_);
  and (_40202_, _03343_, _43223_);
  and (_03344_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_03345_, _03122_, _42867_);
  or (_03346_, _03345_, _03344_);
  and (_40203_, _03346_, _43223_);
  and (_03347_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_03348_, _03122_, _42777_);
  or (_03349_, _03348_, _03347_);
  and (_40204_, _03349_, _43223_);
  and (_03350_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03351_, _03122_, _43028_);
  or (_03352_, _03351_, _03350_);
  and (_40206_, _03352_, _43223_);
  and (_03353_, _03119_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_03354_, _03122_, _42964_);
  or (_03355_, _03354_, _03353_);
  and (_40207_, _03355_, _43223_);
  and (_03356_, _03126_, _42674_);
  and (_03357_, _03356_, _38817_);
  not (_03358_, _03356_);
  and (_03359_, _03358_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or (_03360_, _03359_, _03357_);
  and (_40208_, _03360_, _43223_);
  and (_03361_, _03137_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03362_, _03358_, _38808_);
  nand (_03363_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03364_, _03363_, _03113_);
  or (_03365_, _03364_, _03362_);
  or (_03366_, _03365_, _03361_);
  and (_40209_, _03366_, _43223_);
  and (_03367_, _03358_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_03368_, _03358_, _38801_);
  or (_03369_, _03368_, _03367_);
  and (_40210_, _03369_, _43223_);
  nor (_03370_, _03358_, _38793_);
  and (_03371_, _03138_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or (_03372_, _03371_, _03370_);
  and (_40211_, _03372_, _43223_);
  nor (_03373_, _03358_, _38786_);
  and (_03374_, _03138_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or (_03375_, _03374_, _03373_);
  and (_40212_, _03375_, _43223_);
  nor (_03376_, _03358_, _38778_);
  and (_03377_, _03138_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_03378_, _03377_, _03376_);
  and (_40213_, _03378_, _43223_);
  nor (_03379_, _03358_, _38770_);
  and (_03380_, _03138_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_03381_, _03380_, _03379_);
  and (_40214_, _03381_, _43223_);
  and (_03382_, _03160_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03383_, _03146_, _38817_);
  nand (_03384_, _42674_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_03385_, _03384_, _03152_);
  or (_03386_, _03385_, _03383_);
  or (_03387_, _03386_, _03382_);
  and (_40215_, _03387_, _43223_);
  and (_03388_, _03161_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_03389_, _03148_, _38808_);
  or (_03390_, _03389_, _03388_);
  and (_40217_, _03390_, _43223_);
  nor (_03391_, _03148_, _38801_);
  and (_03392_, _03161_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_03393_, _03392_, _03391_);
  and (_40218_, _03393_, _43223_);
  nor (_03394_, _03148_, _38793_);
  and (_03395_, _03161_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or (_03396_, _03395_, _03394_);
  and (_40219_, _03396_, _43223_);
  nor (_03397_, _03148_, _38786_);
  and (_03398_, _03148_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_03399_, _03398_, _03397_);
  and (_40220_, _03399_, _43223_);
  and (_03400_, _03148_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_03401_, _03148_, _38778_);
  or (_03402_, _03401_, _03400_);
  and (_40221_, _03402_, _43223_);
  nor (_03403_, _03148_, _38770_);
  and (_03404_, _03161_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_03405_, _03404_, _03403_);
  and (_40222_, _03405_, _43223_);
  not (_03406_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03407_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_03408_, _03407_, _03406_);
  and (_03409_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _43223_);
  and (_40283_, _03409_, _03408_);
  nor (_03410_, _03408_, rst);
  nand (_03411_, _03407_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03412_, _03407_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03413_, _03412_, _03411_);
  and (_40285_, _03413_, _03410_);
  not (_03414_, _42989_);
  and (_03415_, _03414_, _43039_);
  not (_03416_, _42721_);
  and (_03417_, _42892_, _03416_);
  and (_03418_, _03417_, _42789_);
  and (_03419_, _03418_, _03415_);
  not (_03420_, _43084_);
  and (_03421_, _39496_, _39483_);
  nor (_03422_, _39496_, _39483_);
  or (_03423_, _03422_, _03421_);
  nor (_03424_, _39522_, _39508_);
  and (_03425_, _39522_, _39508_);
  nor (_03426_, _03425_, _03424_);
  nor (_03427_, _03426_, _03423_);
  and (_03428_, _03426_, _03423_);
  nor (_03429_, _03428_, _03427_);
  and (_03430_, _39546_, _39534_);
  nor (_03431_, _39546_, _39534_);
  nor (_03432_, _03431_, _03430_);
  nor (_03433_, _39557_, _39462_);
  and (_03434_, _39557_, _39462_);
  nor (_03435_, _03434_, _03433_);
  or (_03436_, _03435_, _03432_);
  nand (_03437_, _03435_, _03432_);
  and (_03438_, _03437_, _03436_);
  nor (_03439_, _03438_, _03429_);
  and (_03440_, _03438_, _03429_);
  nor (_03441_, _03440_, _03439_);
  or (_03442_, _03441_, _03420_);
  and (_03443_, _42936_, _42835_);
  or (_03444_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03445_, _03444_, _03443_);
  and (_03446_, _03445_, _03442_);
  nor (_03447_, _42936_, _42835_);
  and (_03448_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not (_03449_, _42936_);
  and (_03450_, _03449_, _42835_);
  and (_03451_, _03450_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_03452_, _03451_, _03448_);
  and (_03453_, _03452_, _03420_);
  nor (_03454_, _03449_, _42835_);
  nor (_03455_, _43084_, _34319_);
  and (_03456_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03457_, _03456_, _03455_);
  and (_03458_, _03457_, _03454_);
  and (_03459_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_03460_, _03450_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_03461_, _03460_, _03459_);
  and (_03462_, _03461_, _43084_);
  or (_03463_, _03462_, _03458_);
  or (_03464_, _03463_, _03453_);
  or (_03465_, _03464_, _03446_);
  and (_03466_, _03465_, _03419_);
  nor (_03467_, _43039_, _42788_);
  and (_03468_, _03417_, _03414_);
  and (_03469_, _03468_, _03467_);
  and (_03470_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_03471_, _43084_, _31281_);
  or (_03472_, _03471_, _03470_);
  and (_03473_, _03472_, _03447_);
  or (_03474_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_03475_, _43084_, _32426_);
  and (_03476_, _03475_, _03443_);
  and (_03477_, _03476_, _03474_);
  or (_03478_, _03477_, _03473_);
  and (_03479_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_03480_, _43084_, _36116_);
  or (_03481_, _03480_, _03479_);
  and (_03482_, _03481_, _03450_);
  nand (_03483_, _43084_, _33841_);
  or (_03484_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03485_, _03484_, _03454_);
  and (_03486_, _03485_, _03483_);
  or (_03487_, _03486_, _03482_);
  or (_03488_, _03487_, _03478_);
  and (_03489_, _03488_, _03469_);
  and (_03490_, _42788_, _03416_);
  and (_03491_, _42989_, _43039_);
  and (_03492_, _03491_, _03490_);
  and (_03493_, _03492_, _42892_);
  nor (_03494_, _01060_, _01210_);
  and (_03495_, _38601_, _38624_);
  or (_03496_, _03495_, _38651_);
  or (_03497_, _03496_, _38718_);
  nor (_03498_, _03497_, _00891_);
  and (_03499_, _38634_, _38571_);
  or (_03500_, _03499_, _00893_);
  nor (_03501_, _03500_, _00959_);
  nor (_03502_, _38658_, _38645_);
  and (_03503_, _03502_, _03501_);
  and (_03504_, _03503_, _00961_);
  and (_03505_, _03504_, _03498_);
  and (_03506_, _03505_, _38684_);
  and (_03507_, _03506_, _03494_);
  nor (_03508_, _03507_, _37039_);
  nor (_03509_, _03508_, p0_in[7]);
  and (_03510_, _03508_, _39570_);
  nor (_03511_, _03510_, _03509_);
  and (_03512_, _03511_, _03420_);
  or (_03514_, _03508_, p0_in[3]);
  not (_03515_, _03508_);
  or (_03516_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03517_, _03516_, _03514_);
  and (_03518_, _03517_, _43084_);
  or (_03519_, _03518_, _03512_);
  and (_03520_, _03519_, _03447_);
  nor (_03521_, _03508_, p0_in[0]);
  and (_03522_, _03508_, _39652_);
  nor (_03523_, _03522_, _03521_);
  or (_03524_, _03523_, _03420_);
  or (_03525_, _03508_, p0_in[4]);
  or (_03526_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03527_, _03526_, _03525_);
  or (_03528_, _03527_, _43084_);
  and (_03529_, _03528_, _03443_);
  and (_03530_, _03529_, _03524_);
  or (_03531_, _03508_, p0_in[6]);
  or (_03532_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03533_, _03532_, _03531_);
  and (_03534_, _03533_, _03420_);
  or (_03535_, _03508_, p0_in[2]);
  or (_03536_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03537_, _03536_, _03535_);
  and (_03538_, _03537_, _43084_);
  or (_03539_, _03538_, _03534_);
  and (_03540_, _03539_, _03454_);
  or (_03541_, _03508_, p0_in[1]);
  or (_03542_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03543_, _03542_, _03541_);
  or (_03544_, _03543_, _03420_);
  or (_03545_, _03508_, p0_in[5]);
  or (_03546_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03547_, _03546_, _03545_);
  or (_03548_, _03547_, _43084_);
  and (_03549_, _03548_, _03450_);
  and (_03550_, _03549_, _03544_);
  or (_03551_, _03550_, _03540_);
  or (_03552_, _03551_, _03530_);
  or (_03553_, _03552_, _03520_);
  and (_03554_, _03553_, _03493_);
  or (_03555_, _03554_, _03489_);
  or (_03556_, _42892_, _42721_);
  nor (_03557_, _03556_, _42788_);
  and (_03558_, _42989_, _43040_);
  and (_03559_, _03558_, _03557_);
  and (_03560_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03561_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03562_, _03561_, _03560_);
  and (_03563_, _03562_, _03447_);
  or (_03564_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nand (_03565_, _43084_, _41086_);
  and (_03566_, _03565_, _03443_);
  and (_03567_, _03566_, _03564_);
  or (_03568_, _03567_, _03563_);
  and (_03569_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03570_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03571_, _03570_, _03569_);
  and (_03572_, _03571_, _03454_);
  or (_03573_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  nand (_03574_, _43084_, _41089_);
  and (_03575_, _03574_, _03450_);
  and (_03576_, _03575_, _03573_);
  or (_03577_, _03576_, _03572_);
  or (_03578_, _03577_, _03568_);
  and (_03579_, _03578_, _03559_);
  nor (_03580_, _42989_, _42721_);
  and (_03581_, _43040_, _42788_);
  and (_03582_, _03581_, _03580_);
  and (_03583_, _03582_, _42892_);
  and (_03584_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03585_, _03450_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03586_, _03585_, _03584_);
  and (_03587_, _03586_, _43084_);
  and (_03588_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03589_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03590_, _03589_, _03588_);
  and (_03591_, _03590_, _03454_);
  and (_03592_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03593_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03594_, _03593_, _03592_);
  and (_03595_, _03594_, _03443_);
  or (_03596_, _03595_, _03591_);
  and (_03597_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03598_, _03450_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03599_, _03598_, _03597_);
  and (_03600_, _03599_, _03420_);
  or (_03601_, _03600_, _03596_);
  or (_03602_, _03601_, _03587_);
  and (_03603_, _03602_, _03583_);
  or (_03604_, _03603_, _03579_);
  or (_03605_, _03604_, _03555_);
  and (_03606_, _03417_, _42989_);
  and (_03607_, _03606_, _03467_);
  nor (_03608_, _03508_, p3_in[7]);
  and (_03609_, _03508_, _39611_);
  nor (_03610_, _03609_, _03608_);
  and (_03611_, _03610_, _03420_);
  or (_03612_, _03508_, p3_in[3]);
  or (_03613_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03614_, _03613_, _03612_);
  and (_03615_, _03614_, _43084_);
  or (_03616_, _03615_, _03611_);
  and (_03617_, _03616_, _03447_);
  nor (_03618_, _03508_, p3_in[0]);
  and (_03619_, _03508_, _40098_);
  nor (_03620_, _03619_, _03618_);
  or (_03621_, _03620_, _03420_);
  or (_03622_, _03508_, p3_in[4]);
  or (_03623_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03624_, _03623_, _03622_);
  or (_03625_, _03624_, _43084_);
  and (_03626_, _03625_, _03443_);
  and (_03627_, _03626_, _03621_);
  or (_03628_, _03627_, _03617_);
  or (_03629_, _03508_, p3_in[5]);
  or (_03630_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03631_, _03630_, _03629_);
  and (_03632_, _03631_, _03420_);
  or (_03633_, _03508_, p3_in[1]);
  or (_03634_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03635_, _03634_, _03633_);
  and (_03636_, _03635_, _43084_);
  or (_03637_, _03636_, _03632_);
  and (_03638_, _03637_, _03450_);
  or (_03639_, _03508_, p3_in[2]);
  or (_03640_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03641_, _03640_, _03639_);
  or (_03642_, _03641_, _03420_);
  or (_03643_, _03508_, p3_in[6]);
  or (_03644_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03645_, _03644_, _03643_);
  or (_03646_, _03645_, _43084_);
  and (_03647_, _03646_, _03454_);
  and (_03648_, _03647_, _03642_);
  or (_03649_, _03648_, _03638_);
  or (_03650_, _03649_, _03628_);
  and (_03651_, _03650_, _03607_);
  and (_03652_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_03653_, _03652_, _43084_);
  and (_03654_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03655_, _03450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_03656_, _03454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03657_, _03656_, _03655_);
  or (_03658_, _03657_, _03654_);
  or (_03659_, _03658_, _03653_);
  and (_03660_, _03490_, _42893_);
  and (_03661_, _03660_, _03415_);
  and (_03662_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_03663_, _03662_, _03420_);
  and (_03664_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03665_, _03450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_03666_, _03454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03667_, _03666_, _03665_);
  or (_03668_, _03667_, _03664_);
  or (_03669_, _03668_, _03663_);
  and (_03670_, _03669_, _03661_);
  and (_03671_, _03670_, _03659_);
  or (_03672_, _03671_, _03651_);
  and (_03673_, _01560_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_03674_, _03606_, _03581_);
  or (_03675_, _03508_, p2_in[1]);
  or (_03676_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03677_, _03676_, _03675_);
  or (_03678_, _03677_, _03420_);
  or (_03679_, _03508_, p2_in[5]);
  or (_03680_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03681_, _03680_, _03679_);
  or (_03682_, _03681_, _43084_);
  and (_03683_, _03682_, _03450_);
  and (_03684_, _03683_, _03678_);
  or (_03685_, _03508_, p2_in[6]);
  or (_03686_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03687_, _03686_, _03685_);
  and (_03688_, _03687_, _03420_);
  or (_03689_, _03508_, p2_in[2]);
  or (_03690_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03691_, _03690_, _03689_);
  and (_03692_, _03691_, _43084_);
  or (_03693_, _03692_, _03688_);
  and (_03694_, _03693_, _03454_);
  nor (_03695_, _03508_, p2_in[7]);
  and (_03696_, _03508_, _39601_);
  nor (_03697_, _03696_, _03695_);
  and (_03698_, _03697_, _03420_);
  or (_03699_, _03508_, p2_in[3]);
  or (_03700_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03701_, _03700_, _03699_);
  and (_03702_, _03701_, _43084_);
  or (_03703_, _03702_, _03698_);
  and (_03704_, _03703_, _03447_);
  nor (_03705_, _03508_, p2_in[0]);
  and (_03706_, _03508_, _40005_);
  nor (_03707_, _03706_, _03705_);
  or (_03708_, _03707_, _03420_);
  or (_03709_, _03508_, p2_in[4]);
  or (_03710_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03711_, _03710_, _03709_);
  or (_03712_, _03711_, _43084_);
  and (_03713_, _03712_, _03443_);
  and (_03715_, _03713_, _03708_);
  or (_03716_, _03715_, _03704_);
  or (_03717_, _03716_, _03694_);
  or (_03718_, _03717_, _03684_);
  and (_03719_, _03718_, _03674_);
  or (_03720_, _03719_, _03673_);
  or (_03721_, _03720_, _03672_);
  or (_03722_, _03721_, _03605_);
  nor (_03723_, _43084_, _40343_);
  and (_03724_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_03725_, _03724_, _03723_);
  and (_03726_, _03725_, _03443_);
  or (_03727_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03728_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03729_, _03728_, _03447_);
  and (_03730_, _03729_, _03727_);
  or (_03731_, _03730_, _03726_);
  and (_03732_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03733_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03734_, _03733_, _03732_);
  and (_03735_, _03734_, _03454_);
  or (_03736_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03737_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_03738_, _03737_, _03450_);
  and (_03739_, _03738_, _03736_);
  or (_03740_, _03739_, _03735_);
  or (_03741_, _03740_, _03731_);
  and (_03742_, _03741_, _03491_);
  nor (_03743_, _43084_, _41067_);
  and (_03744_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03745_, _03744_, _03743_);
  and (_03746_, _03745_, _03443_);
  or (_03747_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03748_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03749_, _03748_, _03447_);
  and (_03750_, _03749_, _03747_);
  or (_03751_, _03750_, _03746_);
  and (_03752_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03753_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03754_, _03753_, _03752_);
  and (_03755_, _03754_, _03454_);
  or (_03756_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_03757_, _03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03758_, _03757_, _03450_);
  and (_03759_, _03758_, _03756_);
  or (_03760_, _03759_, _03755_);
  or (_03761_, _03760_, _03751_);
  and (_03762_, _03761_, _03558_);
  or (_03763_, _03762_, _03742_);
  and (_03764_, _03763_, _03660_);
  and (_03765_, _03557_, _03491_);
  nor (_03766_, _43084_, _41640_);
  and (_03767_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03768_, _03767_, _03766_);
  and (_03769_, _03768_, _03447_);
  or (_03770_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand (_03771_, _43084_, _41657_);
  and (_03772_, _03771_, _03443_);
  and (_03773_, _03772_, _03770_);
  or (_03774_, _03773_, _03769_);
  nor (_03775_, _43084_, _42065_);
  and (_03776_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03777_, _03776_, _03775_);
  and (_03778_, _03777_, _03450_);
  nand (_03779_, _43084_, _42090_);
  or (_03780_, _43084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03781_, _03780_, _03454_);
  and (_03782_, _03781_, _03779_);
  or (_03783_, _03782_, _03778_);
  or (_03784_, _03783_, _03774_);
  and (_03785_, _03784_, _03765_);
  and (_03786_, _42989_, _03416_);
  nand (_03787_, _03786_, _42893_);
  nand (_03788_, _03787_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_03789_, _03788_, _03418_);
  nor (_03790_, _03583_, _03493_);
  nor (_03791_, _03674_, _03661_);
  and (_03792_, _03791_, _03790_);
  and (_03793_, _03792_, _03789_);
  and (_03794_, _03491_, _03418_);
  nor (_03795_, _03508_, p1_in[7]);
  and (_03796_, _03508_, _39586_);
  nor (_03797_, _03796_, _03795_);
  and (_03798_, _03797_, _03420_);
  or (_03799_, _03508_, p1_in[3]);
  or (_03800_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03801_, _03800_, _03799_);
  and (_03802_, _03801_, _43084_);
  or (_03803_, _03802_, _03798_);
  and (_03804_, _03803_, _03447_);
  nor (_03805_, _03508_, p1_in[0]);
  and (_03806_, _03508_, _39922_);
  nor (_03807_, _03806_, _03805_);
  or (_03808_, _03807_, _03420_);
  or (_03809_, _03508_, p1_in[4]);
  or (_03810_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03811_, _03810_, _03809_);
  or (_03812_, _03811_, _43084_);
  and (_03813_, _03812_, _03443_);
  and (_03814_, _03813_, _03808_);
  or (_03815_, _03814_, _03804_);
  or (_03816_, _03508_, p1_in[5]);
  or (_03817_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03818_, _03817_, _03816_);
  and (_03819_, _03818_, _03420_);
  or (_03820_, _03508_, p1_in[1]);
  or (_03821_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03822_, _03821_, _03820_);
  and (_03823_, _03822_, _43084_);
  or (_03824_, _03823_, _03819_);
  and (_03825_, _03824_, _03450_);
  or (_03826_, _03508_, p1_in[2]);
  or (_03827_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03828_, _03827_, _03826_);
  or (_03829_, _03828_, _03420_);
  or (_03830_, _03508_, p1_in[6]);
  or (_03831_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03832_, _03831_, _03830_);
  or (_03833_, _03832_, _43084_);
  and (_03834_, _03833_, _03454_);
  and (_03835_, _03834_, _03829_);
  or (_03836_, _03835_, _03825_);
  or (_03837_, _03836_, _03815_);
  and (_03838_, _03837_, _03794_);
  or (_03839_, _03838_, _03793_);
  or (_03840_, _03839_, _03785_);
  or (_03841_, _03840_, _03764_);
  or (_03842_, _03841_, _03722_);
  or (_03843_, _03842_, _03466_);
  and (_03844_, _03583_, _39408_);
  nor (_03845_, _03844_, _01543_);
  nand (_03846_, _03673_, _31849_);
  and (_03847_, _03846_, _03845_);
  and (_03848_, _03847_, _03843_);
  and (_03849_, _03447_, _42714_);
  and (_03850_, _03450_, _43028_);
  or (_03851_, _03850_, _03849_);
  and (_03852_, _03851_, _03420_);
  nor (_03853_, _43084_, _38786_);
  and (_03854_, _43084_, _38817_);
  or (_03855_, _03854_, _03853_);
  and (_03856_, _03855_, _03443_);
  nor (_03857_, _43084_, _38770_);
  and (_03858_, _43084_, _43074_);
  or (_03859_, _03858_, _03857_);
  and (_03860_, _03859_, _03454_);
  or (_03861_, _03860_, _03856_);
  and (_03862_, _03447_, _42867_);
  and (_03863_, _03450_, _42828_);
  or (_03864_, _03863_, _03862_);
  and (_03865_, _03864_, _43084_);
  or (_03866_, _03865_, _03861_);
  nor (_03867_, _03866_, _03852_);
  nor (_03868_, _03867_, _03845_);
  or (_03869_, _03868_, _03848_);
  and (_40286_, _03869_, _43223_);
  and (_03870_, _42892_, _43084_);
  and (_03871_, _03870_, _03447_);
  and (_03872_, _03871_, _03492_);
  and (_03873_, _03872_, _38885_);
  nor (_03874_, _43040_, _42788_);
  and (_03875_, _03870_, _03443_);
  and (_03876_, _03875_, _03580_);
  and (_03877_, _03876_, _03874_);
  and (_03878_, _03877_, _01517_);
  and (_03879_, _03875_, _03582_);
  and (_03880_, _03879_, _39405_);
  or (_03881_, _03880_, _03878_);
  nor (_03882_, _03881_, _03873_);
  nor (_03883_, _03882_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_03884_, _03883_);
  and (_03885_, _03879_, _39408_);
  not (_03886_, _39418_);
  and (_03887_, _03447_, _03420_);
  nor (_03888_, _03887_, _03886_);
  and (_03889_, _03888_, _01541_);
  nor (_03890_, _03889_, _03885_);
  and (_03891_, _03890_, _01563_);
  and (_03892_, _03891_, _03884_);
  and (_03893_, _03870_, _03454_);
  and (_03894_, _03893_, _03492_);
  and (_03895_, _03894_, _38885_);
  or (_03896_, _03895_, rst);
  nor (_40287_, _03896_, _03892_);
  nand (_03897_, _03895_, _31194_);
  and (_03898_, _03490_, _03415_);
  and (_03899_, _42893_, _43084_);
  and (_03900_, _03899_, _03443_);
  and (_03901_, _03900_, _03898_);
  nor (_03902_, _42892_, _43084_);
  and (_03903_, _03902_, _03443_);
  and (_03904_, _03903_, _03898_);
  nor (_03905_, _03904_, _03901_);
  and (_03906_, _03902_, _03450_);
  and (_03907_, _03906_, _03898_);
  and (_03908_, _03899_, _03454_);
  and (_03909_, _03908_, _03898_);
  nor (_03910_, _03909_, _03907_);
  and (_03911_, _03910_, _03905_);
  and (_03912_, _03899_, _03447_);
  and (_03914_, _03912_, _03898_);
  and (_03915_, _03900_, _03492_);
  nor (_03916_, _03915_, _03914_);
  and (_03917_, _03581_, _03786_);
  and (_03918_, _03900_, _03917_);
  and (_03919_, _03887_, _42892_);
  and (_03920_, _03786_, _03467_);
  and (_03921_, _03920_, _03919_);
  nor (_03922_, _03921_, _03918_);
  and (_03923_, _03922_, _03916_);
  and (_03924_, _03923_, _03911_);
  and (_03925_, _03912_, _03492_);
  and (_03926_, _03899_, _03450_);
  and (_03927_, _03926_, _03492_);
  nor (_03928_, _03927_, _03925_);
  and (_03929_, _03908_, _03492_);
  and (_03930_, _03906_, _03492_);
  nor (_03931_, _03930_, _03929_);
  and (_03932_, _03931_, _03928_);
  and (_03933_, _03903_, _03492_);
  and (_03934_, _03887_, _03493_);
  nor (_03935_, _03934_, _03933_);
  and (_03936_, _03874_, _03786_);
  and (_03937_, _03936_, _03900_);
  and (_03938_, _03926_, _03936_);
  nor (_03939_, _03938_, _03937_);
  and (_03940_, _03939_, _03935_);
  and (_03941_, _03940_, _03932_);
  and (_03942_, _03941_, _03924_);
  nand (_03943_, _03875_, _03786_);
  nor (_03944_, _03894_, _03872_);
  and (_03945_, _03876_, _03467_);
  and (_03946_, _03870_, _03450_);
  and (_03947_, _03946_, _03492_);
  nor (_03948_, _03947_, _03945_);
  and (_03949_, _03948_, _03944_);
  and (_03950_, _03949_, _03943_);
  nor (_03951_, _03879_, _03877_);
  and (_03952_, _03951_, _03950_);
  and (_03953_, _03952_, _03942_);
  nand (_03954_, _01560_, _28139_);
  nor (_03955_, _03954_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not (_03956_, _03887_);
  nand (_03957_, _03956_, _01541_);
  nor (_03958_, _03957_, _03886_);
  or (_03959_, _03958_, _03885_);
  or (_03960_, _03959_, _03955_);
  or (_03961_, _03960_, _03883_);
  nor (_03962_, _03961_, _03953_);
  nor (_03963_, _03962_, _20658_);
  not (_03964_, _03895_);
  nand (_03965_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_03966_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_03967_, _03966_, _03965_);
  nand (_03968_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand (_03969_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_03970_, _03969_, _03968_);
  and (_03971_, _03970_, _03967_);
  nand (_03972_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand (_03973_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_03974_, _03973_, _03972_);
  nand (_03975_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_03976_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03977_, _03976_, _03975_);
  and (_03978_, _03977_, _03974_);
  and (_03979_, _03978_, _03971_);
  nand (_03980_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand (_03981_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_03982_, _03981_, _03980_);
  nand (_03983_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand (_03984_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_03985_, _03984_, _03983_);
  and (_03986_, _03985_, _03982_);
  nand (_03987_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand (_03988_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03989_, _03988_, _03987_);
  nand (_03990_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_03991_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_03992_, _03991_, _03990_);
  and (_03993_, _03992_, _03989_);
  and (_03994_, _03993_, _03986_);
  and (_03995_, _03994_, _03979_);
  nand (_03996_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_03997_, _03947_, _38839_);
  and (_03998_, _03997_, _03996_);
  nand (_03999_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand (_04000_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_04001_, _04000_, _03999_);
  and (_04002_, _04001_, _03998_);
  and (_04003_, _03875_, _03492_);
  nand (_04004_, _04003_, _03511_);
  and (_04005_, _03936_, _03875_);
  nand (_04006_, _04005_, _03797_);
  and (_04007_, _04006_, _04004_);
  and (_04008_, _03875_, _03917_);
  nand (_04009_, _04008_, _03697_);
  and (_04010_, _03920_, _03875_);
  nand (_04011_, _04010_, _03610_);
  and (_04012_, _04011_, _04009_);
  and (_04013_, _04012_, _04007_);
  and (_04015_, _04013_, _04002_);
  nand (_04016_, _03877_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_04017_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_04018_, _04017_, _04016_);
  and (_04019_, _04018_, _04015_);
  nand (_04020_, _04019_, _03995_);
  nand (_04021_, _04020_, _03892_);
  nand (_04022_, _04021_, _03964_);
  or (_04023_, _04022_, _03963_);
  and (_04024_, _04023_, _43223_);
  and (_40288_, _04024_, _03897_);
  nor (_40369_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_04025_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_04026_, _03407_, rst);
  and (_40370_, _04026_, _04025_);
  nor (_04027_, _03407_, _03406_);
  or (_04028_, _04027_, _03408_);
  and (_04029_, _03411_, _43223_);
  and (_40371_, _04029_, _04028_);
  nand (_04030_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_04031_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_04032_, _04031_, _04030_);
  nand (_04033_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_04034_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_04035_, _04034_, _04033_);
  and (_04036_, _04035_, _04032_);
  nand (_04037_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_04038_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_04039_, _04038_, _04037_);
  nand (_04040_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_04041_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_04042_, _04041_, _04040_);
  and (_04043_, _04042_, _04039_);
  and (_04044_, _04043_, _04036_);
  nand (_04045_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_04046_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_04047_, _04046_, _04045_);
  nand (_04048_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_04049_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_04050_, _04049_, _04048_);
  and (_04051_, _04050_, _04047_);
  nand (_04052_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_04053_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_04054_, _04053_, _04052_);
  nand (_04055_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_04056_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_04057_, _04056_, _04055_);
  and (_04058_, _04057_, _04054_);
  and (_04059_, _04058_, _04051_);
  and (_04060_, _04059_, _04044_);
  nand (_04061_, _03947_, _42895_);
  nand (_04062_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_04063_, _04062_, _04061_);
  nand (_04064_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_04065_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_04066_, _04065_, _04064_);
  and (_04067_, _04066_, _04063_);
  nand (_04068_, _04008_, _03707_);
  nand (_04069_, _04010_, _03620_);
  and (_04070_, _04069_, _04068_);
  nand (_04071_, _04005_, _03807_);
  nand (_04072_, _04003_, _03523_);
  and (_04073_, _04072_, _04071_);
  and (_04074_, _04073_, _04070_);
  and (_04075_, _04074_, _04067_);
  nand (_04076_, _03877_, _03441_);
  nand (_04077_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_04078_, _04077_, _04076_);
  and (_04079_, _04078_, _04075_);
  and (_04080_, _04079_, _04060_);
  nor (_04081_, _04080_, _03961_);
  or (_04082_, _03962_, _19489_);
  nand (_04083_, _04082_, _03964_);
  or (_04084_, _04083_, _04081_);
  nand (_04085_, _03895_, _32393_);
  and (_04086_, _04085_, _43223_);
  and (_40373_, _04086_, _04084_);
  and (_04087_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_04088_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_04089_, _04088_, _04087_);
  and (_04090_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_04091_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_04092_, _04091_, _04090_);
  or (_04093_, _04092_, _04089_);
  and (_04094_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_04095_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_04096_, _04095_, _04094_);
  and (_04097_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04098_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_04099_, _04098_, _04097_);
  or (_04100_, _04099_, _04096_);
  or (_04101_, _04100_, _04093_);
  and (_04102_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_04103_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_04104_, _04103_, _04102_);
  and (_04105_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_04106_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_04107_, _04106_, _04105_);
  or (_04108_, _04107_, _04104_);
  and (_04109_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_04111_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_04112_, _04111_, _04109_);
  and (_04113_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_04114_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_04115_, _04114_, _04113_);
  or (_04116_, _04115_, _04112_);
  or (_04117_, _04116_, _04108_);
  or (_04118_, _04117_, _04101_);
  and (_04119_, _03947_, _42810_);
  and (_04120_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_04121_, _04120_, _04119_);
  and (_04122_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_04123_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_04124_, _04123_, _04122_);
  or (_04125_, _04124_, _04121_);
  and (_04126_, _04003_, _03543_);
  and (_04127_, _04005_, _03822_);
  or (_04128_, _04127_, _04126_);
  and (_04129_, _04008_, _03677_);
  and (_04130_, _04010_, _03635_);
  or (_04131_, _04130_, _04129_);
  or (_04132_, _04131_, _04128_);
  or (_04133_, _04132_, _04125_);
  and (_04134_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_04135_, _03877_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_04136_, _04135_, _04134_);
  or (_04137_, _04136_, _04133_);
  or (_04138_, _04137_, _04118_);
  nand (_04139_, _03961_, _20474_);
  and (_04140_, _04139_, _04138_);
  nor (_04141_, _03962_, _20474_);
  or (_04142_, _04141_, _03895_);
  or (_04143_, _04142_, _04140_);
  nand (_04144_, _03895_, _33090_);
  and (_04145_, _04144_, _43223_);
  and (_40374_, _04145_, _04143_);
  and (_04146_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_04147_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_04148_, _04147_, _04146_);
  and (_04149_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04150_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_04151_, _04150_, _04149_);
  or (_04152_, _04151_, _04148_);
  and (_04153_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_04154_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_04155_, _04154_, _04153_);
  and (_04156_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_04157_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_04158_, _04157_, _04156_);
  or (_04159_, _04158_, _04155_);
  or (_04160_, _04159_, _04152_);
  and (_04161_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_04162_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_04163_, _04162_, _04161_);
  and (_04164_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_04165_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_04166_, _04165_, _04164_);
  or (_04167_, _04166_, _04163_);
  and (_04168_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_04169_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_04170_, _04169_, _04168_);
  and (_04171_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_04172_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_04173_, _04172_, _04171_);
  or (_04174_, _04173_, _04170_);
  or (_04175_, _04174_, _04167_);
  or (_04176_, _04175_, _04160_);
  and (_04177_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_04178_, _03947_, _43080_);
  or (_04179_, _04178_, _04177_);
  and (_04180_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_04181_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or (_04182_, _04181_, _04180_);
  or (_04183_, _04182_, _04179_);
  and (_04184_, _04005_, _03828_);
  and (_04185_, _04003_, _03537_);
  or (_04186_, _04185_, _04184_);
  and (_04187_, _04008_, _03691_);
  and (_04188_, _04010_, _03641_);
  or (_04189_, _04188_, _04187_);
  or (_04190_, _04189_, _04186_);
  or (_04191_, _04190_, _04183_);
  and (_04192_, _03877_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_04193_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_04194_, _04193_, _04192_);
  or (_04195_, _04194_, _04191_);
  or (_04196_, _04195_, _04176_);
  nand (_04197_, _03961_, _19128_);
  and (_04198_, _04197_, _04196_);
  nor (_04199_, _03962_, _19128_);
  or (_04200_, _04199_, _03895_);
  or (_04201_, _04200_, _04198_);
  nand (_04202_, _03895_, _33809_);
  and (_04203_, _04202_, _43223_);
  and (_40375_, _04203_, _04201_);
  nand (_04204_, _03895_, _34591_);
  and (_04205_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_04206_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_04207_, _04206_, _04205_);
  and (_04208_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_04210_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_04211_, _04210_, _04208_);
  or (_04212_, _04211_, _04207_);
  and (_04213_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_04214_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_04215_, _04214_, _04213_);
  and (_04216_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_04217_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_04218_, _04217_, _04216_);
  or (_04219_, _04218_, _04215_);
  or (_04220_, _04219_, _04212_);
  and (_04221_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_04222_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_04223_, _04222_, _04221_);
  and (_04224_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_04225_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_04226_, _04225_, _04224_);
  or (_04227_, _04226_, _04223_);
  and (_04228_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_04229_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_04230_, _04229_, _04228_);
  and (_04231_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_04232_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_04233_, _04232_, _04231_);
  or (_04234_, _04233_, _04230_);
  or (_04235_, _04234_, _04227_);
  or (_04236_, _04235_, _04220_);
  and (_04237_, _03947_, _42849_);
  and (_04238_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_04239_, _04238_, _04237_);
  and (_04240_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_04241_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_04242_, _04241_, _04240_);
  or (_04243_, _04242_, _04239_);
  and (_04244_, _04003_, _03517_);
  and (_04245_, _04005_, _03801_);
  or (_04246_, _04245_, _04244_);
  and (_04247_, _04008_, _03701_);
  and (_04248_, _04010_, _03614_);
  or (_04249_, _04248_, _04247_);
  or (_04250_, _04249_, _04246_);
  or (_04251_, _04250_, _04243_);
  and (_04252_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_04253_, _03877_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_04254_, _04253_, _04252_);
  or (_04255_, _04254_, _04251_);
  or (_04256_, _04255_, _04236_);
  nand (_04257_, _03961_, _20159_);
  and (_04258_, _04257_, _04256_);
  nor (_04259_, _03962_, _20159_);
  or (_04260_, _04259_, _03895_);
  or (_04261_, _04260_, _04258_);
  and (_04262_, _04261_, _43223_);
  and (_40376_, _04262_, _04204_);
  and (_04263_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_04264_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_04265_, _04264_, _04263_);
  and (_04266_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_04267_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_04268_, _04267_, _04266_);
  or (_04269_, _04268_, _04265_);
  and (_04270_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_04271_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_04272_, _04271_, _04270_);
  and (_04273_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_04274_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_04275_, _04274_, _04273_);
  or (_04276_, _04275_, _04272_);
  or (_04277_, _04276_, _04269_);
  and (_04278_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_04279_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or (_04280_, _04279_, _04278_);
  and (_04281_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_04282_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_04283_, _04282_, _04281_);
  or (_04284_, _04283_, _04280_);
  and (_04285_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_04286_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_04287_, _04286_, _04285_);
  and (_04288_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_04289_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_04290_, _04289_, _04288_);
  or (_04291_, _04290_, _04287_);
  or (_04292_, _04291_, _04284_);
  or (_04293_, _04292_, _04277_);
  and (_04294_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_04295_, _03947_, _42783_);
  or (_04296_, _04295_, _04294_);
  and (_04297_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_04298_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_04299_, _04298_, _04297_);
  or (_04300_, _04299_, _04296_);
  and (_04301_, _04003_, _03527_);
  and (_04302_, _04005_, _03811_);
  or (_04303_, _04302_, _04301_);
  and (_04304_, _04008_, _03711_);
  and (_04305_, _04010_, _03624_);
  or (_04306_, _04305_, _04304_);
  or (_04307_, _04306_, _04303_);
  or (_04308_, _04307_, _04300_);
  and (_04310_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_04311_, _03877_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_04312_, _04311_, _04310_);
  or (_04313_, _04312_, _04308_);
  or (_04314_, _04313_, _04293_);
  nand (_04315_, _03961_, _19326_);
  and (_04316_, _04315_, _04314_);
  nor (_04317_, _03962_, _19326_);
  or (_04318_, _04317_, _03895_);
  or (_04319_, _04318_, _04316_);
  nand (_04320_, _03895_, _35277_);
  and (_04321_, _04320_, _43223_);
  and (_40377_, _04321_, _04319_);
  and (_04322_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04323_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_04324_, _04323_, _04322_);
  and (_04325_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_04326_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04327_, _04326_, _04325_);
  or (_04328_, _04327_, _04324_);
  and (_04329_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04330_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_04331_, _04330_, _04329_);
  and (_04332_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_04333_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_04334_, _04333_, _04332_);
  or (_04335_, _04334_, _04331_);
  or (_04336_, _04335_, _04328_);
  and (_04337_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_04338_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_04339_, _04338_, _04337_);
  and (_04340_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_04341_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_04342_, _04341_, _04340_);
  or (_04343_, _04342_, _04339_);
  and (_04344_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_04345_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_04346_, _04345_, _04344_);
  and (_04347_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_04348_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_04349_, _04348_, _04347_);
  or (_04350_, _04349_, _04346_);
  or (_04351_, _04350_, _04343_);
  or (_04352_, _04351_, _04336_);
  and (_04353_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_04354_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_04355_, _04354_, _04353_);
  not (_04356_, _38877_);
  and (_04357_, _03947_, _04356_);
  and (_04358_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_04359_, _04358_, _04357_);
  or (_04360_, _04359_, _04355_);
  and (_04361_, _04003_, _03547_);
  and (_04362_, _04005_, _03818_);
  or (_04363_, _04362_, _04361_);
  and (_04364_, _04008_, _03681_);
  and (_04365_, _04010_, _03631_);
  or (_04366_, _04365_, _04364_);
  or (_04367_, _04366_, _04363_);
  or (_04368_, _04367_, _04360_);
  and (_04369_, _03877_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_04370_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_04371_, _04370_, _04369_);
  or (_04372_, _04371_, _04368_);
  or (_04373_, _04372_, _04352_);
  nand (_04374_, _03961_, _20311_);
  and (_04375_, _04374_, _04373_);
  nor (_04376_, _03962_, _20311_);
  or (_04377_, _04376_, _03895_);
  or (_04378_, _04377_, _04375_);
  nand (_04379_, _03895_, _36083_);
  and (_04380_, _04379_, _43223_);
  and (_40378_, _04380_, _04378_);
  and (_04381_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_04382_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_04383_, _04382_, _04381_);
  and (_04384_, _03907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_04385_, _03909_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_04386_, _04385_, _04384_);
  or (_04387_, _04386_, _04383_);
  and (_04388_, _03914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_04389_, _03915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_04390_, _04389_, _04388_);
  and (_04391_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04392_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_04393_, _04392_, _04391_);
  or (_04394_, _04393_, _04390_);
  or (_04395_, _04394_, _04387_);
  and (_04396_, _03925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_04397_, _03927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or (_04398_, _04397_, _04396_);
  and (_04399_, _03930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_04400_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_04401_, _04400_, _04399_);
  or (_04402_, _04401_, _04398_);
  and (_04403_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_04404_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04405_, _04404_, _04403_);
  and (_04406_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_04407_, _03934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_04409_, _04407_, _04406_);
  or (_04410_, _04409_, _04405_);
  or (_04411_, _04410_, _04402_);
  or (_04412_, _04411_, _04395_);
  and (_04413_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_04414_, _03947_, _42970_);
  or (_04415_, _04414_, _04413_);
  and (_04416_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_04417_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_04418_, _04417_, _04416_);
  or (_04419_, _04418_, _04415_);
  and (_04420_, _04003_, _03533_);
  and (_04421_, _04005_, _03832_);
  or (_04422_, _04421_, _04420_);
  and (_04423_, _04008_, _03687_);
  and (_04424_, _04010_, _03645_);
  or (_04425_, _04424_, _04423_);
  or (_04426_, _04425_, _04422_);
  or (_04427_, _04426_, _04419_);
  and (_04428_, _03877_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_04429_, _03879_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_04430_, _04429_, _04428_);
  or (_04431_, _04430_, _04427_);
  or (_04432_, _04431_, _04412_);
  nand (_04433_, _03961_, _19663_);
  and (_04434_, _04433_, _04432_);
  nor (_04435_, _03962_, _19663_);
  or (_04436_, _04435_, _03895_);
  or (_04437_, _04436_, _04434_);
  nand (_04438_, _03895_, _36811_);
  and (_04439_, _04438_, _43223_);
  and (_40379_, _04439_, _04437_);
  and (_40449_, _43121_, _43223_);
  nor (_40452_, _43084_, rst);
  and (_40473_, _43282_, _43223_);
  nor (_40476_, _42936_, rst);
  nor (_40478_, _42835_, rst);
  nor (_04440_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_04441_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04442_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04441_);
  nor (_04443_, _04442_, _04440_);
  nor (_04444_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04441_);
  nor (_04446_, _04445_, _04444_);
  and (_04447_, _04446_, _04443_);
  nor (_04448_, _02324_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04449_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04441_);
  nor (_04450_, _04449_, _04448_);
  nor (_04451_, _04450_, _04447_);
  and (_04452_, _04450_, _04447_);
  nor (_04453_, _04452_, _04451_);
  not (_04454_, _04453_);
  nor (_04455_, _02343_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04456_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04441_);
  or (_04457_, _04456_, _04455_);
  nor (_04458_, _04457_, _04454_);
  not (_04459_, _04443_);
  nor (_04460_, _04446_, _04459_);
  and (_04461_, _04460_, _04458_);
  and (_04462_, _04461_, _00674_);
  and (_04463_, _04458_, _04447_);
  and (_04464_, _04463_, _00588_);
  and (_04465_, _04446_, _04459_);
  and (_04466_, _04457_, _04453_);
  and (_04467_, _04466_, _04465_);
  and (_04468_, _04467_, _00368_);
  or (_04469_, _04468_, _04464_);
  or (_04470_, _04469_, _04462_);
  nor (_04471_, _04446_, _04443_);
  and (_04472_, _04471_, _04466_);
  and (_04473_, _04472_, _00286_);
  and (_04474_, _04466_, _04447_);
  and (_04475_, _04474_, _00245_);
  and (_04476_, _04457_, _04452_);
  and (_04477_, _04476_, _00409_);
  not (_04478_, _04452_);
  nor (_04479_, _04457_, _04478_);
  and (_04480_, _04479_, _00050_);
  or (_04481_, _04480_, _04477_);
  or (_04482_, _04481_, _04475_);
  or (_04483_, _04482_, _04473_);
  and (_04484_, _04471_, _04458_);
  and (_04485_, _04484_, _00633_);
  and (_04486_, _04466_, _04460_);
  and (_04487_, _04486_, _00327_);
  or (_04488_, _04487_, _04485_);
  or (_04489_, _04488_, _04483_);
  nor (_04490_, _04457_, _04452_);
  or (_04491_, _04490_, _04476_);
  and (_04492_, _04491_, _04454_);
  and (_04493_, _04492_, _04465_);
  and (_04494_, _04493_, _00532_);
  nor (_04495_, _04491_, _04453_);
  and (_04496_, _04495_, _04465_);
  and (_04497_, _04496_, _00204_);
  or (_04498_, _04497_, _04494_);
  or (_04499_, _04498_, _04489_);
  or (_04500_, _04499_, _04470_);
  nand (_04501_, _04495_, _04459_);
  and (_04503_, _04495_, _04460_);
  nand (_04504_, _04450_, _04446_);
  nand (_04505_, _04457_, _04451_);
  and (_04506_, _04505_, _04504_);
  or (_04507_, _04506_, _04452_);
  or (_04508_, _04507_, _04467_);
  nor (_04509_, _04508_, _04503_);
  and (_04510_, _04509_, _04501_);
  and (_04511_, _04510_, _00715_);
  and (_04512_, _04492_, _04460_);
  and (_04513_, _04512_, _00491_);
  and (_04514_, _04503_, _00132_);
  or (_04515_, _04514_, _04513_);
  and (_04516_, _04492_, _04471_);
  and (_04517_, _04516_, _00450_);
  and (_04518_, _04495_, _04471_);
  and (_04519_, _04518_, _00091_);
  or (_04520_, _04519_, _04517_);
  or (_04521_, _04520_, _04515_);
  or (_04522_, _04521_, _04511_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04522_, _04500_);
  and (_04523_, _04461_, _00715_);
  and (_04524_, _04463_, _00633_);
  and (_04525_, _04467_, _00409_);
  or (_04526_, _04525_, _04524_);
  or (_04527_, _04526_, _04523_);
  and (_04528_, _04472_, _00327_);
  and (_04529_, _04474_, _00286_);
  and (_04530_, _04476_, _00450_);
  and (_04531_, _04479_, _00091_);
  or (_04532_, _04531_, _04530_);
  or (_04533_, _04532_, _04529_);
  or (_04534_, _04533_, _04528_);
  and (_04535_, _04484_, _00674_);
  and (_04536_, _04486_, _00368_);
  or (_04537_, _04536_, _04535_);
  or (_04538_, _04537_, _04534_);
  and (_04539_, _04493_, _00588_);
  and (_04540_, _04496_, _00245_);
  or (_04541_, _04540_, _04539_);
  or (_04542_, _04541_, _04538_);
  or (_04543_, _04542_, _04527_);
  and (_04544_, _04510_, _00050_);
  and (_04545_, _04512_, _00532_);
  and (_04546_, _04503_, _00204_);
  or (_04547_, _04546_, _04545_);
  and (_04548_, _04516_, _00491_);
  and (_04549_, _04518_, _00132_);
  or (_04550_, _04549_, _04548_);
  or (_04551_, _04550_, _04547_);
  or (_04552_, _04551_, _04544_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04552_, _04543_);
  and (_04553_, _04463_, _00674_);
  and (_04554_, _04484_, _00715_);
  and (_04555_, _04472_, _00368_);
  or (_04556_, _04555_, _04554_);
  or (_04557_, _04556_, _04553_);
  and (_04558_, _04486_, _00409_);
  and (_04559_, _04474_, _00327_);
  and (_04560_, _04476_, _00491_);
  and (_04561_, _04479_, _00132_);
  or (_04562_, _04561_, _04560_);
  or (_04563_, _04562_, _04559_);
  or (_04564_, _04563_, _04558_);
  and (_04565_, _04467_, _00450_);
  and (_04566_, _04461_, _00050_);
  or (_04567_, _04566_, _04565_);
  or (_04568_, _04567_, _04564_);
  and (_04569_, _04493_, _00633_);
  and (_04570_, _04496_, _00286_);
  or (_04571_, _04570_, _04569_);
  or (_04572_, _04571_, _04568_);
  or (_04573_, _04572_, _04557_);
  and (_04574_, _04510_, _00091_);
  and (_04575_, _04512_, _00588_);
  and (_04576_, _04503_, _00245_);
  or (_04577_, _04576_, _04575_);
  and (_04578_, _04516_, _00532_);
  and (_04579_, _04518_, _00204_);
  or (_04580_, _04579_, _04578_);
  or (_04581_, _04580_, _04577_);
  or (_04582_, _04581_, _04574_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04582_, _04573_);
  and (_04583_, _04484_, _00588_);
  and (_04584_, _04461_, _00633_);
  and (_04585_, _04463_, _00532_);
  or (_04586_, _04585_, _04584_);
  or (_04587_, _04586_, _04583_);
  and (_04588_, _04486_, _00286_);
  and (_04589_, _04474_, _00204_);
  and (_04590_, _04479_, _00715_);
  and (_04591_, _04476_, _00368_);
  or (_04592_, _04591_, _04590_);
  or (_04593_, _04592_, _04589_);
  or (_04594_, _04593_, _04588_);
  and (_04595_, _04467_, _00327_);
  and (_04596_, _04472_, _00245_);
  or (_04597_, _04596_, _04595_);
  or (_04598_, _04597_, _04594_);
  and (_04599_, _04512_, _00450_);
  and (_04601_, _04516_, _00409_);
  or (_04602_, _04601_, _04599_);
  or (_04603_, _04602_, _04598_);
  or (_04604_, _04603_, _04587_);
  and (_04605_, _04510_, _00674_);
  and (_04606_, _04493_, _00491_);
  and (_04607_, _04496_, _00132_);
  or (_04608_, _04607_, _04606_);
  and (_04609_, _04518_, _00050_);
  and (_04610_, _04503_, _00091_);
  or (_04611_, _04610_, _04609_);
  or (_04612_, _04611_, _04608_);
  or (_04613_, _04612_, _04605_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04613_, _04604_);
  and (_04614_, _04484_, _00720_);
  and (_04615_, _04463_, _00679_);
  and (_04616_, _04472_, _00373_);
  or (_04617_, _04616_, _04615_);
  or (_04618_, _04617_, _04614_);
  and (_04619_, _04467_, _00455_);
  and (_04620_, _04486_, _00414_);
  or (_04621_, _04620_, _04619_);
  and (_04622_, _04461_, _00055_);
  and (_04623_, _04474_, _00332_);
  and (_04624_, _04476_, _00496_);
  and (_04625_, _04479_, _00138_);
  or (_04626_, _04625_, _04624_);
  or (_04627_, _04626_, _04623_);
  or (_04628_, _04627_, _04622_);
  or (_04629_, _04628_, _04621_);
  and (_04630_, _04512_, _00596_);
  and (_04631_, _04503_, _00250_);
  or (_04632_, _04631_, _04630_);
  or (_04633_, _04632_, _04629_);
  or (_04634_, _04633_, _04618_);
  and (_04635_, _04510_, _00096_);
  and (_04636_, _04516_, _00537_);
  and (_04637_, _04493_, _00638_);
  or (_04638_, _04637_, _04636_);
  and (_04639_, _04496_, _00291_);
  and (_04640_, _04518_, _00209_);
  or (_04641_, _04640_, _04639_);
  or (_04642_, _04641_, _04638_);
  or (_04643_, _04642_, _04635_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04643_, _04634_);
  and (_04644_, _04484_, _00725_);
  and (_04645_, _04463_, _00684_);
  and (_04646_, _04472_, _00378_);
  or (_04647_, _04646_, _04645_);
  or (_04648_, _04647_, _04644_);
  and (_04649_, _04467_, _00460_);
  and (_04650_, _04486_, _00419_);
  or (_04651_, _04650_, _04649_);
  and (_04652_, _04461_, _00060_);
  and (_04653_, _04474_, _00337_);
  and (_04654_, _04476_, _00501_);
  and (_04655_, _04479_, _00149_);
  or (_04656_, _04655_, _04654_);
  or (_04657_, _04656_, _04653_);
  or (_04658_, _04657_, _04652_);
  or (_04659_, _04658_, _04651_);
  and (_04660_, _04512_, _00602_);
  and (_04661_, _04503_, _00255_);
  or (_04662_, _04661_, _04660_);
  or (_04663_, _04662_, _04659_);
  or (_04664_, _04663_, _04648_);
  and (_04665_, _04510_, _00101_);
  and (_04666_, _04516_, _00542_);
  and (_04667_, _04493_, _00643_);
  or (_04668_, _04667_, _04666_);
  and (_04669_, _04496_, _00296_);
  and (_04670_, _04518_, _00214_);
  or (_04671_, _04670_, _04669_);
  or (_04672_, _04671_, _04668_);
  or (_04673_, _04672_, _04665_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04673_, _04664_);
  and (_04674_, _04463_, _00689_);
  and (_04675_, _04484_, _00730_);
  and (_04676_, _04472_, _00383_);
  or (_04677_, _04676_, _04675_);
  or (_04678_, _04677_, _04674_);
  and (_04679_, _04486_, _00424_);
  and (_04680_, _04474_, _00342_);
  and (_04681_, _04476_, _00506_);
  and (_04682_, _04479_, _00160_);
  or (_04683_, _04682_, _04681_);
  or (_04684_, _04683_, _04680_);
  or (_04685_, _04684_, _04679_);
  and (_04686_, _04467_, _00465_);
  and (_04687_, _04461_, _00065_);
  or (_04688_, _04687_, _04686_);
  or (_04689_, _04688_, _04685_);
  and (_04690_, _04493_, _00648_);
  and (_04691_, _04496_, _00301_);
  or (_04692_, _04691_, _04690_);
  or (_04693_, _04692_, _04689_);
  or (_04694_, _04693_, _04678_);
  and (_04695_, _04510_, _00106_);
  and (_04696_, _04512_, _00607_);
  and (_04697_, _04503_, _00260_);
  or (_04698_, _04697_, _04696_);
  and (_04699_, _04516_, _00547_);
  and (_04700_, _04518_, _00219_);
  or (_04701_, _04700_, _04699_);
  or (_04702_, _04701_, _04698_);
  or (_04703_, _04702_, _04695_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04703_, _04694_);
  and (_04704_, _04484_, _00735_);
  and (_04705_, _04463_, _00694_);
  and (_04706_, _04472_, _00388_);
  or (_04707_, _04706_, _04705_);
  or (_04708_, _04707_, _04704_);
  and (_04709_, _04467_, _00470_);
  and (_04710_, _04486_, _00429_);
  or (_04711_, _04710_, _04709_);
  and (_04712_, _04461_, _00070_);
  and (_04713_, _04474_, _00347_);
  and (_04714_, _04476_, _00511_);
  and (_04715_, _04479_, _00171_);
  or (_04716_, _04715_, _04714_);
  or (_04717_, _04716_, _04713_);
  or (_04718_, _04717_, _04712_);
  or (_04719_, _04718_, _04711_);
  and (_04720_, _04512_, _00612_);
  and (_04721_, _04503_, _00265_);
  or (_04722_, _04721_, _04720_);
  or (_04723_, _04722_, _04719_);
  or (_04724_, _04723_, _04708_);
  and (_04725_, _04510_, _00111_);
  and (_04726_, _04516_, _00554_);
  and (_04727_, _04493_, _00653_);
  or (_04728_, _04727_, _04726_);
  and (_04729_, _04496_, _00306_);
  and (_04730_, _04518_, _00224_);
  or (_04731_, _04730_, _04729_);
  or (_04732_, _04731_, _04728_);
  or (_04733_, _04732_, _04725_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04733_, _04724_);
  and (_04734_, _04463_, _00699_);
  and (_04735_, _04484_, _00740_);
  and (_04736_, _04472_, _00393_);
  or (_04737_, _04736_, _04735_);
  or (_04738_, _04737_, _04734_);
  and (_04739_, _04486_, _00434_);
  and (_04740_, _04474_, _00352_);
  and (_04741_, _04476_, _00516_);
  and (_04742_, _04479_, _00182_);
  or (_04743_, _04742_, _04741_);
  or (_04744_, _04743_, _04740_);
  or (_04745_, _04744_, _04739_);
  and (_04746_, _04467_, _00475_);
  and (_04747_, _04461_, _00075_);
  or (_04748_, _04747_, _04746_);
  or (_04749_, _04748_, _04745_);
  and (_04750_, _04493_, _00658_);
  and (_04751_, _04496_, _00311_);
  or (_04752_, _04751_, _04750_);
  or (_04753_, _04752_, _04749_);
  or (_04754_, _04753_, _04738_);
  and (_04755_, _04510_, _00116_);
  and (_04756_, _04512_, _00617_);
  and (_04757_, _04503_, _00270_);
  or (_04758_, _04757_, _04756_);
  and (_04759_, _04516_, _00562_);
  and (_04760_, _04518_, _00229_);
  or (_04761_, _04760_, _04759_);
  or (_04762_, _04761_, _04758_);
  or (_04763_, _04762_, _04755_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _04763_, _04754_);
  and (_04764_, _04484_, _00745_);
  and (_04765_, _04463_, _00704_);
  and (_04766_, _04472_, _00398_);
  or (_04767_, _04766_, _04765_);
  or (_04768_, _04767_, _04764_);
  and (_04769_, _04467_, _00480_);
  and (_04770_, _04486_, _00439_);
  or (_04771_, _04770_, _04769_);
  and (_04772_, _04461_, _00080_);
  and (_04773_, _04474_, _00357_);
  and (_04774_, _04476_, _00521_);
  and (_04775_, _04479_, _00193_);
  or (_04776_, _04775_, _04774_);
  or (_04777_, _04776_, _04773_);
  or (_04778_, _04777_, _04772_);
  or (_04779_, _04778_, _04771_);
  and (_04780_, _04512_, _00622_);
  and (_04781_, _04503_, _00275_);
  or (_04782_, _04781_, _04780_);
  or (_04783_, _04782_, _04779_);
  or (_04784_, _04783_, _04768_);
  and (_04785_, _04510_, _00121_);
  and (_04786_, _04516_, _00570_);
  and (_04787_, _04493_, _00663_);
  or (_04788_, _04787_, _04786_);
  and (_04789_, _04496_, _00316_);
  and (_04790_, _04518_, _00234_);
  or (_04791_, _04790_, _04789_);
  or (_04792_, _04791_, _04788_);
  or (_04793_, _04792_, _04785_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _04793_, _04784_);
  and (_04794_, _04463_, _00709_);
  and (_04795_, _04484_, _00750_);
  and (_04796_, _04472_, _00403_);
  or (_04797_, _04796_, _04795_);
  or (_04798_, _04797_, _04794_);
  and (_04799_, _04486_, _00444_);
  and (_04800_, _04474_, _00362_);
  and (_04801_, _04476_, _00526_);
  and (_04802_, _04479_, _00198_);
  or (_04803_, _04802_, _04801_);
  or (_04804_, _04803_, _04800_);
  or (_04805_, _04804_, _04799_);
  and (_04806_, _04467_, _00485_);
  and (_04807_, _04461_, _00085_);
  or (_04808_, _04807_, _04806_);
  or (_04809_, _04808_, _04805_);
  and (_04810_, _04493_, _00668_);
  and (_04811_, _04496_, _00321_);
  or (_04812_, _04811_, _04810_);
  or (_04813_, _04812_, _04809_);
  or (_04814_, _04813_, _04798_);
  and (_04815_, _04510_, _00126_);
  and (_04816_, _04512_, _00627_);
  and (_04817_, _04503_, _00280_);
  or (_04818_, _04817_, _04816_);
  and (_04819_, _04516_, _00578_);
  and (_04820_, _04518_, _00239_);
  or (_04821_, _04820_, _04819_);
  or (_04822_, _04821_, _04818_);
  or (_04823_, _04822_, _04815_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _04823_, _04814_);
  and (_04824_, _04461_, _00720_);
  and (_04825_, _04463_, _00638_);
  and (_04826_, _04467_, _00414_);
  or (_04827_, _04826_, _04825_);
  or (_04828_, _04827_, _04824_);
  and (_04829_, _04472_, _00332_);
  and (_04830_, _04474_, _00291_);
  and (_04831_, _04476_, _00455_);
  and (_04832_, _04479_, _00096_);
  or (_04833_, _04832_, _04831_);
  or (_04834_, _04833_, _04830_);
  or (_04835_, _04834_, _04829_);
  and (_04836_, _04484_, _00679_);
  and (_04837_, _04486_, _00373_);
  or (_04838_, _04837_, _04836_);
  or (_04839_, _04838_, _04835_);
  and (_04840_, _04493_, _00596_);
  and (_04841_, _04496_, _00250_);
  or (_04842_, _04841_, _04840_);
  or (_04843_, _04842_, _04839_);
  or (_04844_, _04843_, _04828_);
  and (_04845_, _04510_, _00055_);
  and (_04846_, _04512_, _00537_);
  and (_04847_, _04503_, _00209_);
  or (_04848_, _04847_, _04846_);
  and (_04849_, _04516_, _00496_);
  and (_04850_, _04518_, _00138_);
  or (_04851_, _04850_, _04849_);
  or (_04852_, _04851_, _04848_);
  or (_04853_, _04852_, _04845_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _04853_, _04844_);
  and (_04854_, _04484_, _00684_);
  and (_04855_, _04461_, _00725_);
  and (_04856_, _04467_, _00419_);
  or (_04857_, _04856_, _04855_);
  or (_04858_, _04857_, _04854_);
  and (_04859_, _04486_, _00378_);
  and (_04860_, _04472_, _00337_);
  or (_04861_, _04860_, _04859_);
  and (_04862_, _04463_, _00643_);
  and (_04863_, _04474_, _00296_);
  and (_04864_, _04476_, _00460_);
  and (_04865_, _04479_, _00101_);
  or (_04866_, _04865_, _04864_);
  or (_04867_, _04866_, _04863_);
  or (_04868_, _04867_, _04862_);
  or (_04869_, _04868_, _04861_);
  and (_04870_, _04493_, _00602_);
  and (_04871_, _04516_, _00501_);
  or (_04872_, _04871_, _04870_);
  or (_04873_, _04872_, _04869_);
  or (_04874_, _04873_, _04858_);
  and (_04875_, _04510_, _00060_);
  and (_04876_, _04503_, _00214_);
  and (_04877_, _04496_, _00255_);
  or (_04878_, _04877_, _04876_);
  and (_04879_, _04512_, _00542_);
  and (_04880_, _04518_, _00149_);
  or (_04881_, _04880_, _04879_);
  or (_04882_, _04881_, _04878_);
  or (_04883_, _04882_, _04875_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _04883_, _04874_);
  and (_04884_, _04484_, _00689_);
  and (_04885_, _04461_, _00730_);
  and (_04886_, _04463_, _00648_);
  or (_04887_, _04886_, _04885_);
  or (_04888_, _04887_, _04884_);
  and (_04889_, _04486_, _00383_);
  and (_04890_, _04467_, _00424_);
  or (_04891_, _04890_, _04889_);
  and (_04892_, _04472_, _00342_);
  and (_04893_, _04474_, _00301_);
  and (_04894_, _04476_, _00465_);
  and (_04895_, _04479_, _00106_);
  or (_04896_, _04895_, _04894_);
  or (_04897_, _04896_, _04893_);
  or (_04898_, _04897_, _04892_);
  or (_04899_, _04898_, _04891_);
  and (_04900_, _04512_, _00547_);
  and (_04901_, _04496_, _00260_);
  or (_04902_, _04901_, _04900_);
  or (_04903_, _04902_, _04899_);
  or (_04904_, _04903_, _04888_);
  and (_04905_, _04510_, _00065_);
  and (_04906_, _04516_, _00506_);
  and (_04907_, _04503_, _00219_);
  or (_04908_, _04907_, _04906_);
  and (_04909_, _04493_, _00607_);
  and (_04910_, _04518_, _00160_);
  or (_04911_, _04910_, _04909_);
  or (_04912_, _04911_, _04908_);
  or (_04913_, _04912_, _04905_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _04913_, _04904_);
  and (_04914_, _04484_, _00694_);
  and (_04915_, _04461_, _00735_);
  and (_04916_, _04463_, _00653_);
  or (_04917_, _04916_, _04915_);
  or (_04918_, _04917_, _04914_);
  and (_04919_, _04486_, _00388_);
  and (_04920_, _04467_, _00429_);
  or (_04921_, _04920_, _04919_);
  and (_04922_, _04472_, _00347_);
  and (_04923_, _04474_, _00306_);
  and (_04924_, _04476_, _00470_);
  and (_04925_, _04479_, _00111_);
  or (_04926_, _04925_, _04924_);
  or (_04927_, _04926_, _04923_);
  or (_04928_, _04927_, _04922_);
  or (_04929_, _04928_, _04921_);
  and (_04930_, _04512_, _00554_);
  and (_04931_, _04496_, _00265_);
  or (_04932_, _04931_, _04930_);
  or (_04933_, _04932_, _04929_);
  or (_04934_, _04933_, _04918_);
  and (_04935_, _04510_, _00070_);
  and (_04936_, _04516_, _00511_);
  and (_04937_, _04503_, _00224_);
  or (_04938_, _04937_, _04936_);
  and (_04939_, _04493_, _00612_);
  and (_04940_, _04518_, _00171_);
  or (_04941_, _04940_, _04939_);
  or (_04942_, _04941_, _04938_);
  or (_04943_, _04942_, _04935_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _04943_, _04934_);
  and (_04944_, _04484_, _00699_);
  and (_04945_, _04461_, _00740_);
  and (_04946_, _04463_, _00658_);
  or (_04947_, _04946_, _04945_);
  or (_04948_, _04947_, _04944_);
  and (_04949_, _04486_, _00393_);
  and (_04950_, _04467_, _00434_);
  or (_04951_, _04950_, _04949_);
  and (_04952_, _04472_, _00352_);
  and (_04953_, _04474_, _00311_);
  and (_04954_, _04476_, _00475_);
  and (_04955_, _04479_, _00116_);
  or (_04956_, _04955_, _04954_);
  or (_04957_, _04956_, _04953_);
  or (_04958_, _04957_, _04952_);
  or (_04959_, _04958_, _04951_);
  and (_04960_, _04512_, _00562_);
  and (_04961_, _04518_, _00182_);
  or (_04962_, _04961_, _04960_);
  or (_04963_, _04962_, _04959_);
  or (_04964_, _04963_, _04948_);
  and (_04965_, _04510_, _00075_);
  and (_04966_, _04516_, _00516_);
  and (_04967_, _04503_, _00229_);
  or (_04968_, _04967_, _04966_);
  and (_04969_, _04493_, _00617_);
  and (_04970_, _04496_, _00270_);
  or (_04971_, _04970_, _04969_);
  or (_04972_, _04971_, _04968_);
  or (_04973_, _04972_, _04965_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _04973_, _04964_);
  and (_04974_, _04461_, _00745_);
  and (_04975_, _04463_, _00663_);
  and (_04976_, _04467_, _00439_);
  or (_04977_, _04976_, _04975_);
  or (_04978_, _04977_, _04974_);
  and (_04979_, _04472_, _00357_);
  and (_04980_, _04474_, _00316_);
  and (_04981_, _04476_, _00480_);
  and (_04982_, _04479_, _00121_);
  or (_04983_, _04982_, _04981_);
  or (_04984_, _04983_, _04980_);
  or (_04985_, _04984_, _04979_);
  and (_04986_, _04484_, _00704_);
  and (_04987_, _04486_, _00398_);
  or (_04988_, _04987_, _04986_);
  or (_04989_, _04988_, _04985_);
  and (_04990_, _04493_, _00622_);
  and (_04991_, _04496_, _00275_);
  or (_04992_, _04991_, _04990_);
  or (_04993_, _04992_, _04989_);
  or (_04994_, _04993_, _04978_);
  and (_04995_, _04510_, _00080_);
  and (_04996_, _04512_, _00570_);
  and (_04997_, _04503_, _00234_);
  or (_04998_, _04997_, _04996_);
  and (_04999_, _04516_, _00521_);
  and (_05000_, _04518_, _00193_);
  or (_05001_, _05000_, _04999_);
  or (_05002_, _05001_, _04998_);
  or (_05003_, _05002_, _04995_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _05003_, _04994_);
  and (_05004_, _04484_, _00709_);
  and (_05005_, _04461_, _00750_);
  and (_05006_, _04463_, _00668_);
  or (_05007_, _05006_, _05005_);
  or (_05008_, _05007_, _05004_);
  and (_05009_, _04486_, _00403_);
  and (_05010_, _04467_, _00444_);
  or (_05011_, _05010_, _05009_);
  and (_05012_, _04472_, _00362_);
  and (_05013_, _04474_, _00321_);
  and (_05014_, _04476_, _00485_);
  and (_05015_, _04479_, _00126_);
  or (_05016_, _05015_, _05014_);
  or (_05017_, _05016_, _05013_);
  or (_05018_, _05017_, _05012_);
  or (_05019_, _05018_, _05011_);
  and (_05020_, _04512_, _00578_);
  and (_05021_, _04518_, _00198_);
  or (_05022_, _05021_, _05020_);
  or (_05023_, _05022_, _05019_);
  or (_05024_, _05023_, _05008_);
  and (_05025_, _04510_, _00085_);
  and (_05026_, _04516_, _00526_);
  and (_05027_, _04503_, _00239_);
  or (_05028_, _05027_, _05026_);
  and (_05029_, _04493_, _00627_);
  and (_05030_, _04496_, _00280_);
  or (_05031_, _05030_, _05029_);
  or (_05032_, _05031_, _05028_);
  or (_05033_, _05032_, _05025_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _05033_, _05024_);
  and (_05034_, _04486_, _00291_);
  and (_05035_, _04467_, _00332_);
  and (_05036_, _04472_, _00250_);
  or (_05037_, _05036_, _05035_);
  or (_05038_, _05037_, _05034_);
  and (_05040_, _04484_, _00596_);
  and (_05042_, _04463_, _00537_);
  or (_05044_, _05042_, _05040_);
  and (_05046_, _04461_, _00638_);
  and (_05048_, _04474_, _00209_);
  and (_05050_, _04479_, _00720_);
  and (_05052_, _04476_, _00373_);
  or (_05053_, _05052_, _05050_);
  or (_05054_, _05053_, _05048_);
  or (_05055_, _05054_, _05046_);
  or (_05056_, _05055_, _05044_);
  and (_05057_, _04503_, _00096_);
  and (_05058_, _04512_, _00455_);
  or (_05060_, _05058_, _05057_);
  or (_05061_, _05060_, _05056_);
  or (_05063_, _05061_, _05038_);
  and (_05064_, _04510_, _00679_);
  and (_05065_, _04496_, _00138_);
  and (_05067_, _04516_, _00414_);
  or (_05068_, _05067_, _05065_);
  and (_05069_, _04518_, _00055_);
  and (_05071_, _04493_, _00496_);
  or (_05072_, _05071_, _05069_);
  or (_05073_, _05072_, _05068_);
  or (_05075_, _05073_, _05064_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _05075_, _05063_);
  and (_05076_, _04472_, _00255_);
  and (_05078_, _04461_, _00643_);
  and (_05079_, _04467_, _00337_);
  or (_05080_, _05079_, _05078_);
  or (_05082_, _05080_, _05076_);
  and (_05083_, _04484_, _00602_);
  and (_05084_, _04474_, _00214_);
  and (_05086_, _04479_, _00725_);
  and (_05087_, _04476_, _00378_);
  or (_05088_, _05087_, _05086_);
  or (_05090_, _05088_, _05084_);
  or (_05091_, _05090_, _05083_);
  and (_05092_, _04463_, _00542_);
  and (_05093_, _04486_, _00296_);
  or (_05094_, _05093_, _05092_);
  or (_05095_, _05094_, _05091_);
  and (_05096_, _04512_, _00460_);
  and (_05097_, _04516_, _00419_);
  or (_05098_, _05097_, _05096_);
  or (_05099_, _05098_, _05095_);
  or (_05100_, _05099_, _05082_);
  and (_05101_, _04510_, _00684_);
  and (_05102_, _04503_, _00101_);
  and (_05103_, _04496_, _00149_);
  or (_05104_, _05103_, _05102_);
  and (_05105_, _04493_, _00501_);
  and (_05106_, _04518_, _00060_);
  or (_05107_, _05106_, _05105_);
  or (_05108_, _05107_, _05104_);
  or (_05109_, _05108_, _05101_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _05109_, _05100_);
  and (_05111_, _04472_, _00260_);
  and (_05112_, _04461_, _00648_);
  and (_05114_, _04467_, _00342_);
  or (_05115_, _05114_, _05112_);
  or (_05116_, _05115_, _05111_);
  and (_05118_, _04484_, _00607_);
  and (_05119_, _04474_, _00219_);
  and (_05120_, _04479_, _00730_);
  and (_05122_, _04476_, _00383_);
  or (_05123_, _05122_, _05120_);
  or (_05124_, _05123_, _05119_);
  or (_05126_, _05124_, _05118_);
  and (_05127_, _04463_, _00547_);
  and (_05128_, _04486_, _00301_);
  or (_05130_, _05128_, _05127_);
  or (_05131_, _05130_, _05126_);
  and (_05132_, _04512_, _00465_);
  and (_05134_, _04516_, _00424_);
  or (_05135_, _05134_, _05132_);
  or (_05136_, _05135_, _05131_);
  or (_05138_, _05136_, _05116_);
  and (_05139_, _04510_, _00689_);
  and (_05140_, _04503_, _00106_);
  and (_05142_, _04496_, _00160_);
  or (_05143_, _05142_, _05140_);
  and (_05144_, _04493_, _00506_);
  and (_05145_, _04518_, _00065_);
  or (_05146_, _05145_, _05144_);
  or (_05147_, _05146_, _05143_);
  or (_05148_, _05147_, _05139_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _05148_, _05138_);
  and (_05149_, _04484_, _00612_);
  and (_05150_, _04461_, _00653_);
  and (_05151_, _04463_, _00554_);
  or (_05152_, _05151_, _05150_);
  or (_05153_, _05152_, _05149_);
  and (_05154_, _04467_, _00347_);
  and (_05155_, _04486_, _00306_);
  or (_05156_, _05155_, _05154_);
  and (_05157_, _04472_, _00265_);
  and (_05158_, _04474_, _00224_);
  and (_05159_, _04479_, _00735_);
  and (_05160_, _04476_, _00388_);
  or (_05161_, _05160_, _05159_);
  or (_05163_, _05161_, _05158_);
  or (_05164_, _05163_, _05157_);
  or (_05166_, _05164_, _05156_);
  and (_05167_, _04512_, _00470_);
  and (_05168_, _04516_, _00429_);
  or (_05170_, _05168_, _05167_);
  or (_05171_, _05170_, _05166_);
  or (_05172_, _05171_, _05153_);
  and (_05174_, _04510_, _00694_);
  and (_05175_, _04493_, _00511_);
  and (_05176_, _04496_, _00171_);
  or (_05178_, _05176_, _05175_);
  and (_05179_, _04518_, _00070_);
  and (_05180_, _04503_, _00111_);
  or (_05182_, _05180_, _05179_);
  or (_05183_, _05182_, _05178_);
  or (_05184_, _05183_, _05174_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _05184_, _05172_);
  and (_05186_, _04484_, _00617_);
  and (_05187_, _04461_, _00658_);
  and (_05189_, _04463_, _00562_);
  or (_05190_, _05189_, _05187_);
  or (_05191_, _05190_, _05186_);
  and (_05193_, _04467_, _00352_);
  and (_05194_, _04486_, _00311_);
  or (_05195_, _05194_, _05193_);
  and (_05196_, _04472_, _00270_);
  and (_05197_, _04474_, _00229_);
  and (_05198_, _04479_, _00740_);
  and (_05199_, _04476_, _00393_);
  or (_05200_, _05199_, _05198_);
  or (_05201_, _05200_, _05197_);
  or (_05202_, _05201_, _05196_);
  or (_05203_, _05202_, _05195_);
  and (_05204_, _04512_, _00475_);
  and (_05205_, _04503_, _00116_);
  or (_05206_, _05205_, _05204_);
  or (_05207_, _05206_, _05203_);
  or (_05208_, _05207_, _05191_);
  and (_05209_, _04510_, _00699_);
  and (_05210_, _04493_, _00516_);
  and (_05211_, _04496_, _00182_);
  or (_05212_, _05211_, _05210_);
  and (_05213_, _04516_, _00434_);
  and (_05215_, _04518_, _00075_);
  or (_05216_, _05215_, _05213_);
  or (_05218_, _05216_, _05212_);
  or (_05219_, _05218_, _05209_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _05219_, _05208_);
  and (_05221_, _04484_, _00622_);
  and (_05222_, _04461_, _00663_);
  and (_05223_, _04463_, _00570_);
  or (_05225_, _05223_, _05222_);
  or (_05226_, _05225_, _05221_);
  and (_05227_, _04486_, _00316_);
  and (_05229_, _04467_, _00357_);
  or (_05230_, _05229_, _05227_);
  and (_05231_, _04472_, _00275_);
  and (_05233_, _04474_, _00234_);
  and (_05234_, _04479_, _00745_);
  and (_05235_, _04476_, _00398_);
  or (_05237_, _05235_, _05234_);
  or (_05238_, _05237_, _05233_);
  or (_05239_, _05238_, _05231_);
  or (_05241_, _05239_, _05230_);
  and (_05242_, _04512_, _00480_);
  and (_05243_, _04503_, _00121_);
  or (_05245_, _05243_, _05242_);
  or (_05246_, _05245_, _05241_);
  or (_05247_, _05246_, _05226_);
  and (_05248_, _04510_, _00704_);
  and (_05249_, _04493_, _00521_);
  and (_05250_, _04496_, _00193_);
  or (_05251_, _05250_, _05249_);
  and (_05252_, _04516_, _00439_);
  and (_05253_, _04518_, _00080_);
  or (_05254_, _05253_, _05252_);
  or (_05255_, _05254_, _05251_);
  or (_05256_, _05255_, _05248_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _05256_, _05247_);
  and (_05257_, _04484_, _00627_);
  and (_05258_, _04461_, _00668_);
  and (_05259_, _04463_, _00578_);
  or (_05260_, _05259_, _05258_);
  or (_05261_, _05260_, _05257_);
  and (_05262_, _04486_, _00321_);
  and (_05263_, _04467_, _00362_);
  or (_05264_, _05263_, _05262_);
  and (_05266_, _04472_, _00280_);
  and (_05267_, _04474_, _00239_);
  and (_05269_, _04479_, _00750_);
  and (_05270_, _04476_, _00403_);
  or (_05271_, _05270_, _05269_);
  or (_05273_, _05271_, _05267_);
  or (_05274_, _05273_, _05266_);
  or (_05275_, _05274_, _05264_);
  and (_05277_, _04512_, _00485_);
  and (_05278_, _04516_, _00444_);
  or (_05279_, _05278_, _05277_);
  or (_05281_, _05279_, _05275_);
  or (_05282_, _05281_, _05261_);
  and (_05283_, _04510_, _00709_);
  and (_05285_, _04493_, _00526_);
  and (_05286_, _04496_, _00198_);
  or (_05287_, _05286_, _05285_);
  and (_05289_, _04518_, _00085_);
  and (_05290_, _04503_, _00126_);
  or (_05291_, _05290_, _05289_);
  or (_05293_, _05291_, _05287_);
  or (_05294_, _05293_, _05283_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _05294_, _05282_);
  and (_05296_, _04461_, _00679_);
  and (_05297_, _04463_, _00596_);
  and (_05298_, _04467_, _00373_);
  or (_05299_, _05298_, _05297_);
  or (_05300_, _05299_, _05296_);
  and (_05301_, _04512_, _00496_);
  and (_05302_, _04516_, _00455_);
  or (_05303_, _05302_, _05301_);
  and (_05304_, _04472_, _00291_);
  and (_05305_, _04486_, _00332_);
  or (_05306_, _05305_, _05304_);
  and (_05307_, _04484_, _00638_);
  and (_05308_, _04474_, _00250_);
  and (_05309_, _04476_, _00414_);
  and (_05310_, _04479_, _00055_);
  or (_05311_, _05310_, _05309_);
  or (_05312_, _05311_, _05308_);
  or (_05313_, _05312_, _05307_);
  or (_05314_, _05313_, _05306_);
  or (_05315_, _05314_, _05303_);
  or (_05316_, _05315_, _05300_);
  and (_05318_, _04510_, _00720_);
  and (_05319_, _04493_, _00537_);
  and (_05321_, _04518_, _00096_);
  or (_05322_, _05321_, _05319_);
  and (_05323_, _04503_, _00138_);
  and (_05325_, _04496_, _00209_);
  or (_05326_, _05325_, _05323_);
  or (_05327_, _05326_, _05322_);
  or (_05329_, _05327_, _05318_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05329_, _05316_);
  and (_05330_, _04484_, _00643_);
  and (_05332_, _04461_, _00684_);
  and (_05333_, _04463_, _00602_);
  or (_05334_, _05333_, _05332_);
  or (_05336_, _05334_, _05330_);
  and (_05337_, _04472_, _00296_);
  and (_05338_, _04474_, _00255_);
  and (_05340_, _04476_, _00419_);
  and (_05341_, _04479_, _00060_);
  or (_05342_, _05341_, _05340_);
  or (_05344_, _05342_, _05338_);
  or (_05345_, _05344_, _05337_);
  and (_05346_, _04467_, _00378_);
  and (_05348_, _04486_, _00337_);
  or (_05349_, _05348_, _05346_);
  or (_05350_, _05349_, _05345_);
  and (_05351_, _04512_, _00501_);
  and (_05352_, _04496_, _00214_);
  or (_05353_, _05352_, _05351_);
  or (_05354_, _05353_, _05350_);
  or (_05355_, _05354_, _05336_);
  and (_05356_, _04510_, _00725_);
  and (_05357_, _04516_, _00460_);
  and (_05358_, _04503_, _00149_);
  or (_05359_, _05358_, _05357_);
  and (_05360_, _04493_, _00542_);
  and (_05361_, _04518_, _00101_);
  or (_05362_, _05361_, _05360_);
  or (_05363_, _05362_, _05359_);
  or (_05364_, _05363_, _05356_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05364_, _05355_);
  and (_05365_, _04461_, _00689_);
  and (_05366_, _04484_, _00648_);
  or (_05367_, _05366_, _05365_);
  and (_05369_, _04486_, _00342_);
  or (_05370_, _05369_, _05367_);
  and (_05372_, _04472_, _00301_);
  and (_05373_, _04474_, _00260_);
  and (_05374_, _04476_, _00424_);
  and (_05376_, _04479_, _00065_);
  or (_05377_, _05376_, _05374_);
  or (_05378_, _05377_, _05373_);
  or (_05380_, _05378_, _05372_);
  and (_05381_, _04463_, _00607_);
  and (_05382_, _04467_, _00383_);
  or (_05384_, _05382_, _05381_);
  or (_05385_, _05384_, _05380_);
  and (_05386_, _04512_, _00506_);
  and (_05388_, _04518_, _00106_);
  or (_05389_, _05388_, _05386_);
  or (_05390_, _05389_, _05385_);
  or (_05392_, _05390_, _05370_);
  and (_05393_, _04510_, _00730_);
  and (_05394_, _04516_, _00465_);
  and (_05396_, _04503_, _00160_);
  or (_05397_, _05396_, _05394_);
  and (_05398_, _04493_, _00547_);
  and (_05400_, _04496_, _00219_);
  or (_05401_, _05400_, _05398_);
  or (_05402_, _05401_, _05397_);
  or (_05403_, _05402_, _05393_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05403_, _05392_);
  and (_05404_, _04461_, _00694_);
  and (_05405_, _04463_, _00612_);
  and (_05406_, _04467_, _00388_);
  or (_05407_, _05406_, _05405_);
  or (_05408_, _05407_, _05404_);
  and (_05409_, _04472_, _00306_);
  and (_05410_, _04474_, _00265_);
  and (_05411_, _04476_, _00429_);
  and (_05412_, _04479_, _00070_);
  or (_05413_, _05412_, _05411_);
  or (_05414_, _05413_, _05410_);
  or (_05415_, _05414_, _05409_);
  and (_05416_, _04484_, _00653_);
  and (_05417_, _04486_, _00347_);
  or (_05418_, _05417_, _05416_);
  or (_05419_, _05418_, _05415_);
  and (_05421_, _04493_, _00554_);
  and (_05422_, _04496_, _00224_);
  or (_05424_, _05422_, _05421_);
  or (_05425_, _05424_, _05419_);
  or (_05426_, _05425_, _05408_);
  and (_05428_, _04510_, _00735_);
  and (_05429_, _04512_, _00511_);
  and (_05430_, _04503_, _00171_);
  or (_05432_, _05430_, _05429_);
  and (_05433_, _04516_, _00470_);
  and (_05434_, _04518_, _00111_);
  or (_05436_, _05434_, _05433_);
  or (_05437_, _05436_, _05432_);
  or (_05438_, _05437_, _05428_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05438_, _05426_);
  and (_05440_, _04461_, _00699_);
  and (_05441_, _04463_, _00617_);
  and (_05443_, _04467_, _00393_);
  or (_05444_, _05443_, _05441_);
  or (_05445_, _05444_, _05440_);
  and (_05447_, _04472_, _00311_);
  and (_05448_, _04474_, _00270_);
  and (_05449_, _04476_, _00434_);
  and (_05451_, _04479_, _00075_);
  or (_05452_, _05451_, _05449_);
  or (_05453_, _05452_, _05448_);
  or (_05454_, _05453_, _05447_);
  and (_05455_, _04484_, _00658_);
  and (_05456_, _04486_, _00352_);
  or (_05457_, _05456_, _05455_);
  or (_05458_, _05457_, _05454_);
  and (_05459_, _04493_, _00562_);
  and (_05460_, _04496_, _00229_);
  or (_05461_, _05460_, _05459_);
  or (_05462_, _05461_, _05458_);
  or (_05463_, _05462_, _05445_);
  and (_05464_, _04510_, _00740_);
  and (_05465_, _04512_, _00516_);
  and (_05466_, _04503_, _00182_);
  or (_05467_, _05466_, _05465_);
  and (_05468_, _04516_, _00475_);
  and (_05469_, _04518_, _00116_);
  or (_05470_, _05469_, _05468_);
  or (_05471_, _05470_, _05467_);
  or (_05473_, _05471_, _05464_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05473_, _05463_);
  and (_05475_, _04486_, _00357_);
  and (_05476_, _04484_, _00663_);
  and (_05477_, _04467_, _00398_);
  or (_05479_, _05477_, _05476_);
  or (_05480_, _05479_, _05475_);
  and (_05481_, _04472_, _00316_);
  and (_05483_, _04474_, _00275_);
  and (_05484_, _04476_, _00439_);
  and (_05485_, _04479_, _00080_);
  or (_05487_, _05485_, _05484_);
  or (_05488_, _05487_, _05483_);
  or (_05489_, _05488_, _05481_);
  and (_05491_, _04461_, _00704_);
  and (_05492_, _04463_, _00622_);
  or (_05493_, _05492_, _05491_);
  or (_05495_, _05493_, _05489_);
  and (_05496_, _04512_, _00521_);
  and (_05497_, _04503_, _00193_);
  or (_05499_, _05497_, _05496_);
  or (_05500_, _05499_, _05495_);
  or (_05501_, _05500_, _05480_);
  and (_05503_, _04510_, _00745_);
  and (_05504_, _04516_, _00480_);
  and (_05505_, _04518_, _00121_);
  or (_05506_, _05505_, _05504_);
  and (_05507_, _04493_, _00570_);
  and (_05508_, _04496_, _00234_);
  or (_05509_, _05508_, _05507_);
  or (_05510_, _05509_, _05506_);
  or (_05511_, _05510_, _05503_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05511_, _05501_);
  and (_05512_, _04484_, _00668_);
  and (_05513_, _04461_, _00709_);
  and (_05514_, _04463_, _00627_);
  or (_05515_, _05514_, _05513_);
  or (_05516_, _05515_, _05512_);
  and (_05517_, _04472_, _00321_);
  and (_05518_, _04474_, _00280_);
  and (_05519_, _04476_, _00444_);
  and (_05520_, _04479_, _00085_);
  or (_05521_, _05520_, _05519_);
  or (_05522_, _05521_, _05518_);
  or (_05524_, _05522_, _05517_);
  and (_05525_, _04467_, _00403_);
  and (_05527_, _04486_, _00362_);
  or (_05528_, _05527_, _05525_);
  or (_05529_, _05528_, _05524_);
  and (_05531_, _04512_, _00526_);
  and (_05532_, _04518_, _00126_);
  or (_05533_, _05532_, _05531_);
  or (_05535_, _05533_, _05529_);
  or (_05536_, _05535_, _05516_);
  and (_05537_, _04510_, _00750_);
  and (_05539_, _04516_, _00485_);
  and (_05540_, _04503_, _00198_);
  or (_05541_, _05540_, _05539_);
  and (_05543_, _04493_, _00578_);
  and (_05544_, _04496_, _00239_);
  or (_05545_, _05544_, _05543_);
  or (_05547_, _05545_, _05541_);
  or (_05548_, _05547_, _05537_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05548_, _05536_);
  not (_05550_, \oc8051_golden_model_1.PC [1]);
  and (_05551_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_05552_, \oc8051_golden_model_1.PC [2]);
  and (_05554_, _05552_, \oc8051_golden_model_1.PC [3]);
  and (_05555_, _05554_, _05551_);
  nand (_05556_, _05555_, _00547_);
  not (_05557_, \oc8051_golden_model_1.PC [0]);
  and (_05558_, \oc8051_golden_model_1.PC [1], _05557_);
  and (_05559_, _05558_, _05554_);
  nand (_05560_, _05559_, _00506_);
  and (_05561_, _05560_, _05556_);
  not (_05562_, \oc8051_golden_model_1.PC [3]);
  and (_05563_, \oc8051_golden_model_1.PC [2], _05562_);
  and (_05564_, _05563_, _05551_);
  nand (_05565_, _05564_, _00383_);
  and (_05566_, _05563_, _05558_);
  nand (_05567_, _05566_, _00342_);
  and (_05568_, _05567_, _05565_);
  and (_05569_, _05568_, _05561_);
  and (_05570_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_05571_, _05570_, _05551_);
  nand (_05572_, _05571_, _00730_);
  and (_05573_, _05570_, _05558_);
  nand (_05574_, _05573_, _00689_);
  and (_05576_, _05574_, _05572_);
  nor (_05577_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_05579_, _05577_, _05551_);
  nand (_05580_, _05579_, _00219_);
  and (_05581_, _05577_, _05558_);
  nand (_05583_, _05581_, _00160_);
  and (_05584_, _05583_, _05580_);
  and (_05585_, _05584_, _05576_);
  and (_05587_, _05585_, _05569_);
  and (_05588_, _05550_, \oc8051_golden_model_1.PC [0]);
  and (_05589_, _05588_, _05570_);
  nand (_05591_, _05589_, _00648_);
  nor (_05592_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and (_05593_, _05592_, _05570_);
  nand (_05595_, _05593_, _00607_);
  and (_05596_, _05595_, _05591_);
  and (_05597_, _05577_, _05592_);
  nand (_05599_, _05597_, _00065_);
  and (_05600_, _05577_, _05588_);
  nand (_05601_, _05600_, _00106_);
  and (_05603_, _05601_, _05599_);
  and (_05604_, _05603_, _05596_);
  and (_05605_, _05588_, _05554_);
  nand (_05607_, _05605_, _00465_);
  and (_05608_, _05592_, _05554_);
  nand (_05609_, _05608_, _00424_);
  and (_05610_, _05609_, _05607_);
  and (_05611_, _05588_, _05563_);
  nand (_05612_, _05611_, _00301_);
  and (_05613_, _05592_, _05563_);
  nand (_05614_, _05613_, _00260_);
  and (_05615_, _05614_, _05612_);
  and (_05616_, _05615_, _05610_);
  and (_05617_, _05616_, _05604_);
  nand (_05618_, _05617_, _05587_);
  nand (_05619_, _05555_, _00554_);
  nand (_05620_, _05559_, _00511_);
  and (_05621_, _05620_, _05619_);
  nand (_05622_, _05564_, _00388_);
  nand (_05623_, _05566_, _00347_);
  and (_05624_, _05623_, _05622_);
  and (_05625_, _05624_, _05621_);
  nand (_05626_, _05571_, _00735_);
  nand (_05627_, _05573_, _00694_);
  and (_05629_, _05627_, _05626_);
  nand (_05630_, _05579_, _00224_);
  nand (_05632_, _05581_, _00171_);
  and (_05633_, _05632_, _05630_);
  and (_05634_, _05633_, _05629_);
  and (_05636_, _05634_, _05625_);
  nand (_05637_, _05589_, _00653_);
  nand (_05638_, _05593_, _00612_);
  and (_05640_, _05638_, _05637_);
  nand (_05641_, _05597_, _00070_);
  nand (_05642_, _05600_, _00111_);
  and (_05644_, _05642_, _05641_);
  and (_05645_, _05644_, _05640_);
  nand (_05646_, _05605_, _00470_);
  nand (_05648_, _05608_, _00429_);
  and (_05649_, _05648_, _05646_);
  nand (_05650_, _05611_, _00306_);
  nand (_05652_, _05613_, _00265_);
  and (_05653_, _05652_, _05650_);
  and (_05654_, _05653_, _05649_);
  and (_05656_, _05654_, _05645_);
  nand (_05657_, _05656_, _05636_);
  or (_05658_, _05657_, _05618_);
  nand (_05660_, _05555_, _00537_);
  nand (_05661_, _05559_, _00496_);
  and (_05662_, _05661_, _05660_);
  nand (_05663_, _05564_, _00373_);
  nand (_05664_, _05566_, _00332_);
  and (_05665_, _05664_, _05663_);
  and (_05666_, _05665_, _05662_);
  nand (_05667_, _05571_, _00720_);
  nand (_05668_, _05573_, _00679_);
  and (_05669_, _05668_, _05667_);
  nand (_05670_, _05579_, _00209_);
  nand (_05671_, _05581_, _00138_);
  and (_05672_, _05671_, _05670_);
  and (_05673_, _05672_, _05669_);
  and (_05674_, _05673_, _05666_);
  nand (_05675_, _05589_, _00638_);
  nand (_05676_, _05593_, _00596_);
  and (_05677_, _05676_, _05675_);
  nand (_05678_, _05597_, _00055_);
  nand (_05679_, _05600_, _00096_);
  and (_05680_, _05679_, _05678_);
  and (_05682_, _05680_, _05677_);
  nand (_05683_, _05605_, _00455_);
  nand (_05685_, _05608_, _00414_);
  and (_05686_, _05685_, _05683_);
  nand (_05687_, _05611_, _00291_);
  nand (_05689_, _05613_, _00250_);
  and (_05690_, _05689_, _05687_);
  and (_05691_, _05690_, _05686_);
  and (_05693_, _05691_, _05682_);
  and (_05694_, _05693_, _05674_);
  nand (_05695_, _05555_, _00542_);
  nand (_05697_, _05559_, _00501_);
  and (_05698_, _05697_, _05695_);
  nand (_05699_, _05564_, _00378_);
  nand (_05701_, _05566_, _00337_);
  and (_05702_, _05701_, _05699_);
  and (_05703_, _05702_, _05698_);
  nand (_05705_, _05571_, _00725_);
  nand (_05706_, _05573_, _00684_);
  and (_05707_, _05706_, _05705_);
  nand (_05709_, _05579_, _00214_);
  nand (_05710_, _05581_, _00149_);
  and (_05711_, _05710_, _05709_);
  and (_05713_, _05711_, _05707_);
  and (_05714_, _05713_, _05703_);
  nand (_05715_, _05589_, _00643_);
  nand (_05716_, _05593_, _00602_);
  and (_05717_, _05716_, _05715_);
  nand (_05718_, _05597_, _00060_);
  nand (_05719_, _05600_, _00101_);
  and (_05720_, _05719_, _05718_);
  and (_05721_, _05720_, _05717_);
  nand (_05722_, _05605_, _00460_);
  nand (_05723_, _05608_, _00419_);
  and (_05724_, _05723_, _05722_);
  nand (_05725_, _05611_, _00296_);
  nand (_05726_, _05613_, _00255_);
  and (_05727_, _05726_, _05725_);
  and (_05728_, _05727_, _05724_);
  and (_05729_, _05728_, _05721_);
  nand (_05730_, _05729_, _05714_);
  or (_05731_, _05730_, _05694_);
  or (_05732_, _05731_, _05658_);
  not (_05733_, _05732_);
  nand (_05735_, _05555_, _00562_);
  nand (_05736_, _05559_, _00516_);
  and (_05738_, _05736_, _05735_);
  nand (_05739_, _05564_, _00393_);
  nand (_05740_, _05566_, _00352_);
  and (_05742_, _05740_, _05739_);
  and (_05743_, _05742_, _05738_);
  nand (_05744_, _05571_, _00740_);
  nand (_05746_, _05573_, _00699_);
  and (_05747_, _05746_, _05744_);
  nand (_05748_, _05579_, _00229_);
  nand (_05750_, _05581_, _00182_);
  and (_05751_, _05750_, _05748_);
  and (_05752_, _05751_, _05747_);
  and (_05754_, _05752_, _05743_);
  nand (_05755_, _05589_, _00658_);
  nand (_05756_, _05593_, _00617_);
  and (_05758_, _05756_, _05755_);
  nand (_05759_, _05597_, _00075_);
  nand (_05760_, _05600_, _00116_);
  and (_05762_, _05760_, _05759_);
  and (_05763_, _05762_, _05758_);
  nand (_05764_, _05605_, _00475_);
  nand (_05766_, _05608_, _00434_);
  and (_05767_, _05766_, _05764_);
  nand (_05768_, _05611_, _00311_);
  nand (_05769_, _05613_, _00270_);
  and (_05770_, _05769_, _05768_);
  and (_05771_, _05770_, _05767_);
  and (_05772_, _05771_, _05763_);
  nand (_05773_, _05772_, _05754_);
  nand (_05774_, _05555_, _00570_);
  nand (_05775_, _05559_, _00521_);
  and (_05776_, _05775_, _05774_);
  nand (_05777_, _05564_, _00398_);
  nand (_05778_, _05566_, _00357_);
  and (_05779_, _05778_, _05777_);
  and (_05780_, _05779_, _05776_);
  nand (_05781_, _05571_, _00745_);
  nand (_05782_, _05573_, _00704_);
  and (_05783_, _05782_, _05781_);
  nand (_05784_, _05579_, _00234_);
  nand (_05785_, _05581_, _00193_);
  and (_05786_, _05785_, _05784_);
  and (_05788_, _05786_, _05783_);
  and (_05789_, _05788_, _05780_);
  nand (_05791_, _05589_, _00663_);
  nand (_05792_, _05593_, _00622_);
  and (_05793_, _05792_, _05791_);
  nand (_05795_, _05597_, _00080_);
  nand (_05796_, _05600_, _00121_);
  and (_05797_, _05796_, _05795_);
  and (_05799_, _05797_, _05793_);
  nand (_05800_, _05605_, _00480_);
  nand (_05801_, _05608_, _00439_);
  and (_05803_, _05801_, _05800_);
  nand (_05804_, _05611_, _00316_);
  nand (_05805_, _05613_, _00275_);
  and (_05807_, _05805_, _05804_);
  and (_05808_, _05807_, _05803_);
  and (_05809_, _05808_, _05799_);
  and (_05811_, _05809_, _05789_);
  or (_05812_, _05811_, _05773_);
  not (_05813_, _05812_);
  nand (_05815_, _05555_, _00578_);
  nand (_05816_, _05559_, _00526_);
  and (_05817_, _05816_, _05815_);
  nand (_05819_, _05564_, _00403_);
  nand (_05820_, _05566_, _00362_);
  and (_05821_, _05820_, _05819_);
  and (_05822_, _05821_, _05817_);
  nand (_05823_, _05571_, _00750_);
  nand (_05824_, _05573_, _00709_);
  and (_05825_, _05824_, _05823_);
  nand (_05826_, _05579_, _00239_);
  nand (_05827_, _05581_, _00198_);
  and (_05828_, _05827_, _05826_);
  and (_05829_, _05828_, _05825_);
  and (_05830_, _05829_, _05822_);
  nand (_05831_, _05589_, _00668_);
  nand (_05832_, _05593_, _00627_);
  and (_05833_, _05832_, _05831_);
  nand (_05834_, _05597_, _00085_);
  nand (_05835_, _05600_, _00126_);
  and (_05836_, _05835_, _05834_);
  and (_05837_, _05836_, _05833_);
  nand (_05838_, _05605_, _00485_);
  nand (_05839_, _05608_, _00444_);
  and (_05841_, _05839_, _05838_);
  nand (_05842_, _05611_, _00321_);
  nand (_05844_, _05613_, _00280_);
  and (_05845_, _05844_, _05842_);
  and (_05846_, _05845_, _05841_);
  and (_05848_, _05846_, _05837_);
  nand (_05849_, _05848_, _05830_);
  nand (_05850_, _05555_, _00532_);
  nand (_05852_, _05559_, _00491_);
  and (_05853_, _05852_, _05850_);
  nand (_05854_, _05564_, _00368_);
  nand (_05856_, _05566_, _00327_);
  and (_05857_, _05856_, _05854_);
  and (_05858_, _05857_, _05853_);
  nand (_05860_, _05571_, _00715_);
  nand (_05861_, _05573_, _00674_);
  and (_05862_, _05861_, _05860_);
  nand (_05864_, _05579_, _00204_);
  nand (_05865_, _05581_, _00132_);
  and (_05866_, _05865_, _05864_);
  and (_05868_, _05866_, _05862_);
  and (_05869_, _05868_, _05858_);
  nand (_05870_, _05589_, _00633_);
  nand (_05872_, _05593_, _00588_);
  and (_05873_, _05872_, _05870_);
  nand (_05874_, _05597_, _00050_);
  nand (_05875_, _05600_, _00091_);
  and (_05876_, _05875_, _05874_);
  and (_05877_, _05876_, _05873_);
  nand (_05878_, _05605_, _00450_);
  nand (_05879_, _05608_, _00409_);
  and (_05880_, _05879_, _05878_);
  nand (_05881_, _05611_, _00286_);
  nand (_05882_, _05613_, _00245_);
  and (_05883_, _05882_, _05881_);
  and (_05884_, _05883_, _05880_);
  and (_05885_, _05884_, _05877_);
  and (_05886_, _05885_, _05869_);
  and (_05887_, _05886_, _05849_);
  and (_05888_, _05887_, _05813_);
  and (_05889_, _05888_, _05733_);
  not (_05890_, _05889_);
  and (_05891_, _05772_, _05754_);
  or (_05892_, _05811_, _05891_);
  not (_05893_, _05892_);
  and (_05894_, _05893_, _05887_);
  and (_05895_, _05894_, _05733_);
  nand (_05896_, _05809_, _05789_);
  or (_05897_, _05896_, _05773_);
  or (_05898_, _05886_, _05849_);
  nor (_05899_, _05898_, _05897_);
  and (_05900_, _05899_, _05733_);
  nor (_05901_, _05900_, _05895_);
  and (_05902_, _05901_, _05890_);
  and (_05903_, _05848_, _05830_);
  and (_05904_, _05886_, _05903_);
  not (_05905_, _05897_);
  and (_05906_, _05905_, _05904_);
  and (_05907_, _05733_, _05906_);
  not (_05908_, _05907_);
  or (_05909_, _05896_, _05891_);
  not (_05910_, _05909_);
  and (_05911_, _05910_, _05904_);
  and (_05912_, _05733_, _05911_);
  not (_05913_, _05912_);
  not (_05914_, _05904_);
  or (_05915_, _05892_, _05914_);
  or (_05916_, _05915_, _05732_);
  not (_05917_, _05887_);
  or (_05918_, _05917_, _05909_);
  or (_05919_, _05918_, _05732_);
  and (_05920_, _05919_, _05916_);
  or (_05921_, _05917_, _05897_);
  or (_05922_, _05921_, _05732_);
  or (_05923_, _05812_, _05914_);
  or (_05924_, _05923_, _05732_);
  and (_05925_, _05924_, _05922_);
  and (_05926_, _05925_, _05920_);
  and (_05927_, _05926_, _05913_);
  and (_05928_, _05927_, _05908_);
  and (_05929_, _05928_, _05902_);
  or (_05930_, _05929_, _05550_);
  not (_05931_, _05658_);
  not (_05932_, _05694_);
  and (_05933_, _05730_, _05932_);
  and (_05934_, _05933_, _05931_);
  and (_05935_, _05934_, _05899_);
  and (_05936_, \oc8051_golden_model_1.ACC [0], _05557_);
  not (_05937_, \oc8051_golden_model_1.ACC [1]);
  nor (_05938_, _05588_, _05558_);
  nor (_05939_, _05938_, _05937_);
  and (_05940_, _05938_, _05937_);
  nor (_05941_, _05940_, _05939_);
  and (_05942_, _05941_, _05936_);
  nor (_05943_, _05941_, _05936_);
  nor (_05944_, _05943_, _05942_);
  and (_05945_, _05944_, _05935_);
  or (_05946_, _05898_, _05892_);
  or (_05947_, _05946_, _05732_);
  or (_05948_, _05886_, _05903_);
  or (_05949_, _05948_, _05909_);
  or (_05950_, _05949_, _05732_);
  and (_05951_, _05950_, _05947_);
  or (_05952_, _05948_, _05897_);
  or (_05953_, _05952_, _05732_);
  or (_05954_, _05948_, _05812_);
  or (_05955_, _05954_, _05732_);
  and (_05956_, _05955_, _05953_);
  or (_05957_, _05898_, _05812_);
  or (_05958_, _05957_, _05732_);
  or (_05959_, _05948_, _05892_);
  or (_05960_, _05959_, _05732_);
  and (_05961_, _05960_, _05958_);
  and (_05962_, _05961_, _05956_);
  nand (_05963_, _05962_, _05951_);
  not (_05964_, _05731_);
  not (_05965_, _05657_);
  and (_05966_, _05965_, _05618_);
  and (_05967_, _05966_, _05964_);
  and (_05968_, _05967_, _05899_);
  nor (_05969_, _05898_, _05909_);
  and (_05970_, _05969_, _05733_);
  nor (_05971_, _05970_, _05968_);
  not (_05972_, _05971_);
  or (_05973_, _05972_, _05963_);
  nand (_05974_, _05973_, \oc8051_golden_model_1.PC [1]);
  not (_05975_, _05935_);
  and (_05976_, _05969_, _05934_);
  not (_05977_, _05976_);
  not (_05978_, _05938_);
  or (_05979_, _05963_, _05978_);
  nand (_05980_, _05979_, _05977_);
  and (_05981_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  and (_05982_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_05983_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_05984_, _05983_, _05982_);
  and (_05985_, _05984_, _05981_);
  nor (_05986_, _05984_, _05981_);
  nor (_05987_, _05986_, _05985_);
  nand (_05988_, _05987_, _05976_);
  and (_05989_, _05988_, _05971_);
  nand (_05990_, _05989_, _05980_);
  nand (_05991_, _05990_, _05975_);
  nand (_05992_, _05991_, _05929_);
  and (_05993_, _05992_, _05974_);
  or (_05994_, _05993_, _05945_);
  nand (_05995_, _05994_, _05930_);
  or (_05996_, _05929_, \oc8051_golden_model_1.PC [0]);
  not (_05997_, \oc8051_golden_model_1.ACC [0]);
  and (_05998_, _05997_, \oc8051_golden_model_1.PC [0]);
  nor (_05999_, _05998_, _05936_);
  and (_06000_, _05999_, _05935_);
  nand (_06001_, _05973_, _05557_);
  not (_06002_, _05929_);
  or (_06003_, _05963_, _05557_);
  and (_06004_, _06003_, _05977_);
  nor (_06005_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_06006_, _06005_, _05981_);
  nand (_06007_, _06006_, _05976_);
  nand (_06008_, _06007_, _05971_);
  or (_06009_, _06008_, _06004_);
  and (_06010_, _06009_, _05975_);
  or (_06011_, _06010_, _06002_);
  and (_06012_, _06011_, _06001_);
  or (_06013_, _06012_, _06000_);
  and (_06014_, _06013_, _05996_);
  and (_06015_, _06014_, _05995_);
  and (_06016_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_06017_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_06018_, _06017_, _06016_);
  not (_06019_, _06018_);
  and (_06020_, _06019_, _05973_);
  and (_06021_, _05962_, _05951_);
  and (_06022_, _05551_, \oc8051_golden_model_1.PC [2]);
  nor (_06023_, _05551_, \oc8051_golden_model_1.PC [2]);
  nor (_06024_, _06023_, _06022_);
  nor (_06025_, _06024_, _05976_);
  and (_06026_, _06025_, _06021_);
  nor (_06027_, _05985_, _05982_);
  and (_06028_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06029_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06030_, _06029_, _06028_);
  not (_06031_, _06030_);
  nor (_06032_, _06031_, _06027_);
  and (_06033_, _06031_, _06027_);
  nor (_06034_, _06033_, _06032_);
  not (_06035_, _06034_);
  and (_06036_, _06035_, _05976_);
  or (_06037_, _06036_, _06026_);
  and (_06038_, _06037_, _05971_);
  or (_06039_, _06038_, _05935_);
  or (_06040_, _06039_, _06020_);
  not (_06041_, _05902_);
  nor (_06042_, _05942_, _05939_);
  and (_06043_, _06024_, \oc8051_golden_model_1.ACC [2]);
  nor (_06044_, _06024_, \oc8051_golden_model_1.ACC [2]);
  nor (_06045_, _06044_, _06043_);
  not (_06046_, _06045_);
  nor (_06047_, _06046_, _06042_);
  and (_06048_, _06046_, _06042_);
  nor (_06049_, _06048_, _06047_);
  and (_06050_, _06049_, _05935_);
  nor (_06051_, _06050_, _06041_);
  nand (_06052_, _06051_, _06040_);
  not (_06053_, _05928_);
  nor (_06054_, _06018_, _05902_);
  nor (_06055_, _06054_, _06053_);
  nand (_06056_, _06055_, _06052_);
  nor (_06057_, _06019_, _05928_);
  not (_06058_, _06057_);
  and (_06059_, _06058_, _06056_);
  nor (_06060_, _06047_, _06043_);
  nor (_06061_, _06022_, _05562_);
  nor (_06062_, _06061_, _05564_);
  nor (_06063_, _06062_, \oc8051_golden_model_1.ACC [3]);
  and (_06064_, _06062_, \oc8051_golden_model_1.ACC [3]);
  nor (_06065_, _06064_, _06063_);
  not (_06066_, _06065_);
  and (_06067_, _06066_, _06060_);
  nor (_06068_, _06066_, _06060_);
  nor (_06069_, _06068_, _06067_);
  nor (_06070_, _06069_, _05975_);
  not (_06071_, _06062_);
  or (_06072_, _05963_, _06071_);
  and (_06073_, _05570_, \oc8051_golden_model_1.PC [1]);
  nor (_06074_, _06016_, \oc8051_golden_model_1.PC [3]);
  nor (_06075_, _06074_, _06073_);
  or (_06076_, _06075_, _06021_);
  and (_06077_, _06076_, _06072_);
  nand (_06078_, _06077_, _05977_);
  nor (_06079_, _06032_, _06028_);
  and (_06080_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_06081_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_06082_, _06081_, _06080_);
  not (_06083_, _06082_);
  nor (_06084_, _06083_, _06079_);
  and (_06085_, _06083_, _06079_);
  nor (_06086_, _06085_, _06084_);
  nand (_06087_, _06086_, _05976_);
  and (_06088_, _06087_, _05971_);
  nand (_06089_, _06088_, _06078_);
  or (_06090_, _06075_, _05971_);
  and (_06091_, _06090_, _05975_);
  and (_06092_, _06091_, _06089_);
  or (_06093_, _06092_, _06070_);
  and (_06094_, _06093_, _05929_);
  not (_06095_, _06075_);
  nor (_06096_, _06095_, _05929_);
  nor (_06097_, _06096_, _06094_);
  and (_06098_, _06097_, _06059_);
  and (_06099_, _06098_, _06015_);
  and (_06100_, _06099_, _00101_);
  and (_06101_, _05994_, _05930_);
  nand (_06102_, _06013_, _05996_);
  and (_06103_, _06102_, _06101_);
  and (_06104_, _06098_, _06103_);
  and (_06105_, _06104_, _00149_);
  nor (_06106_, _06105_, _06100_);
  nand (_06107_, _06058_, _06056_);
  or (_06108_, _06096_, _06094_);
  and (_06109_, _06108_, _06107_);
  and (_06110_, _06109_, _06103_);
  and (_06111_, _06110_, _00684_);
  and (_06112_, _06097_, _06107_);
  and (_06113_, _06103_, _06112_);
  and (_06114_, _06113_, _00337_);
  nor (_06115_, _06114_, _06111_);
  and (_06116_, _06115_, _06106_);
  and (_06117_, _06014_, _06101_);
  and (_06118_, _06098_, _06117_);
  and (_06119_, _06118_, _00214_);
  and (_06120_, _06102_, _05995_);
  and (_06121_, _06120_, _06112_);
  and (_06122_, _06121_, _00255_);
  nor (_06123_, _06122_, _06119_);
  and (_06124_, _06108_, _06059_);
  and (_06125_, _06124_, _06117_);
  and (_06126_, _06125_, _00542_);
  and (_06127_, _06120_, _06124_);
  and (_06128_, _06127_, _00419_);
  nor (_06129_, _06128_, _06126_);
  and (_06130_, _06129_, _06123_);
  and (_06131_, _06130_, _06116_);
  and (_06132_, _06120_, _06109_);
  and (_06133_, _06132_, _00602_);
  and (_06134_, _06124_, _06015_);
  and (_06135_, _06134_, _00460_);
  nor (_06136_, _06135_, _06133_);
  and (_06137_, _06109_, _06117_);
  and (_06138_, _06137_, _00725_);
  and (_06139_, _06015_, _06109_);
  and (_06140_, _06139_, _00643_);
  nor (_06141_, _06140_, _06138_);
  and (_06142_, _06141_, _06136_);
  and (_06143_, _06124_, _06103_);
  and (_06144_, _06143_, _00501_);
  and (_06145_, _06098_, _06120_);
  and (_06146_, _06145_, _00060_);
  nor (_06147_, _06146_, _06144_);
  and (_06148_, _06112_, _06117_);
  and (_06149_, _06148_, _00378_);
  and (_06150_, _06015_, _06112_);
  and (_06151_, _06150_, _00296_);
  nor (_06152_, _06151_, _06149_);
  and (_06153_, _06152_, _06147_);
  and (_06154_, _06153_, _06142_);
  and (_06155_, _06154_, _06131_);
  not (_06156_, _06155_);
  nand (_06157_, _06148_, _00368_);
  nand (_06158_, _06113_, _00327_);
  and (_06159_, _06158_, _06157_);
  nand (_06160_, _06137_, _00715_);
  nand (_06161_, _06134_, _00450_);
  and (_06162_, _06161_, _06160_);
  and (_06163_, _06162_, _06159_);
  nand (_06164_, _06125_, _00532_);
  nand (_06165_, _06150_, _00286_);
  and (_06166_, _06165_, _06164_);
  nand (_06167_, _06145_, _00050_);
  nand (_06168_, _06099_, _00091_);
  and (_06169_, _06168_, _06167_);
  and (_06170_, _06169_, _06166_);
  and (_06171_, _06170_, _06163_);
  nand (_06172_, _06132_, _00588_);
  nand (_06173_, _06143_, _00491_);
  and (_06174_, _06173_, _06172_);
  nand (_06175_, _06127_, _00409_);
  nand (_06176_, _06121_, _00245_);
  and (_06177_, _06176_, _06175_);
  and (_06178_, _06177_, _06174_);
  nand (_06179_, _06110_, _00674_);
  nand (_06180_, _06104_, _00132_);
  and (_06181_, _06180_, _06179_);
  nand (_06182_, _06139_, _00633_);
  nand (_06183_, _06118_, _00204_);
  and (_06184_, _06183_, _06182_);
  and (_06185_, _06184_, _06181_);
  and (_06186_, _06185_, _06178_);
  nand (_06187_, _06186_, _06171_);
  and (_06188_, _05967_, _05906_);
  not (_06189_, _06188_);
  nor (_06190_, _06189_, _06187_);
  and (_06191_, _06190_, _06156_);
  and (_06192_, _05657_, _05618_);
  not (_06193_, _05730_);
  and (_06194_, _06193_, _06192_);
  and (_06195_, _06194_, _05906_);
  not (_06196_, _06195_);
  and (_06197_, _06193_, _05694_);
  and (_06198_, _05931_, _06197_);
  and (_06199_, _06198_, _05911_);
  and (_06200_, _06148_, _00393_);
  and (_06201_, _06118_, _00229_);
  nor (_06202_, _06201_, _06200_);
  and (_06203_, _06139_, _00658_);
  and (_06204_, _06127_, _00434_);
  nor (_06205_, _06204_, _06203_);
  and (_06206_, _06205_, _06202_);
  and (_06207_, _06104_, _00182_);
  and (_06208_, _06099_, _00116_);
  nor (_06209_, _06208_, _06207_);
  and (_06210_, _06150_, _00311_);
  and (_06211_, _06121_, _00270_);
  nor (_06212_, _06211_, _06210_);
  and (_06213_, _06212_, _06209_);
  and (_06214_, _06213_, _06206_);
  and (_06215_, _06125_, _00562_);
  and (_06216_, _06143_, _00516_);
  nor (_06217_, _06216_, _06215_);
  and (_06218_, _06137_, _00740_);
  and (_06219_, _06134_, _00475_);
  nor (_06220_, _06219_, _06218_);
  and (_06221_, _06220_, _06217_);
  and (_06222_, _06113_, _00352_);
  and (_06223_, _06145_, _00075_);
  nor (_06224_, _06223_, _06222_);
  and (_06225_, _06110_, _00699_);
  and (_06226_, _06132_, _00617_);
  nor (_06227_, _06226_, _06225_);
  and (_06228_, _06227_, _06224_);
  and (_06229_, _06228_, _06221_);
  and (_06230_, _06229_, _06214_);
  nor (_06231_, _06230_, _06187_);
  and (_06232_, _06231_, _06199_);
  not (_06233_, \oc8051_golden_model_1.SP [1]);
  and (_06234_, _06233_, \oc8051_golden_model_1.SP [0]);
  not (_06235_, \oc8051_golden_model_1.SP [0]);
  and (_06236_, \oc8051_golden_model_1.SP [1], _06235_);
  nor (_06237_, _06236_, _06234_);
  or (_06238_, _06237_, _05916_);
  and (_06239_, _05730_, _05694_);
  and (_06240_, _05931_, _06239_);
  and (_06241_, _06240_, _05969_);
  not (_06242_, _06241_);
  nor (_06243_, _06242_, _06187_);
  not (_06244_, _06230_);
  nand (_06245_, _06244_, _06243_);
  not (_06246_, _05952_);
  and (_06247_, _06246_, _06198_);
  not (_06248_, _06237_);
  and (_06249_, _06248_, _06247_);
  not (_06250_, _05949_);
  and (_06251_, _05967_, _06250_);
  not (_06252_, _06251_);
  nor (_06253_, _06252_, _06187_);
  nand (_06254_, _06253_, _06156_);
  not (_06255_, _05959_);
  and (_06256_, _05966_, _05730_);
  and (_06257_, _06256_, _06255_);
  not (_06258_, _05960_);
  not (_06259_, _05923_);
  and (_06260_, _06240_, _06259_);
  not (_06261_, _06260_);
  nand (_06262_, _06148_, _00388_);
  nand (_06263_, _06104_, _00171_);
  and (_06264_, _06263_, _06262_);
  nand (_06265_, _06139_, _00653_);
  nand (_06266_, _06132_, _00612_);
  and (_06267_, _06266_, _06265_);
  and (_06268_, _06267_, _06264_);
  nand (_06269_, _06113_, _00347_);
  nand (_06270_, _06150_, _00306_);
  and (_06271_, _06270_, _06269_);
  nand (_06272_, _06145_, _00070_);
  nand (_06273_, _06099_, _00111_);
  and (_06274_, _06273_, _06272_);
  and (_06275_, _06274_, _06271_);
  and (_06276_, _06275_, _06268_);
  nand (_06277_, _06125_, _00554_);
  nand (_06278_, _06143_, _00511_);
  and (_06279_, _06278_, _06277_);
  nand (_06280_, _06137_, _00735_);
  nand (_06281_, _06134_, _00470_);
  and (_06282_, _06281_, _06280_);
  and (_06283_, _06282_, _06279_);
  nand (_06284_, _06121_, _00265_);
  nand (_06285_, _06118_, _00224_);
  and (_06286_, _06285_, _06284_);
  nand (_06287_, _06110_, _00694_);
  nand (_06288_, _06127_, _00429_);
  and (_06289_, _06288_, _06287_);
  and (_06290_, _06289_, _06286_);
  and (_06291_, _06290_, _06283_);
  and (_06292_, _06291_, _06276_);
  and (_06293_, _05967_, _06259_);
  and (_06294_, _06293_, _06292_);
  not (_06295_, _06293_);
  and (_06296_, _06150_, _00321_);
  and (_06297_, _06118_, _00239_);
  nor (_06298_, _06297_, _06296_);
  and (_06299_, _06139_, _00668_);
  and (_06300_, _06132_, _00627_);
  nor (_06301_, _06300_, _06299_);
  and (_06302_, _06301_, _06298_);
  and (_06303_, _06104_, _00198_);
  and (_06304_, _06099_, _00126_);
  nor (_06305_, _06304_, _06303_);
  and (_06306_, _06113_, _00362_);
  and (_06307_, _06121_, _00280_);
  nor (_06308_, _06307_, _06306_);
  and (_06309_, _06308_, _06305_);
  and (_06310_, _06309_, _06302_);
  and (_06311_, _06137_, _00750_);
  and (_06312_, _06110_, _00709_);
  nor (_06313_, _06312_, _06311_);
  and (_06314_, _06143_, _00526_);
  and (_06315_, _06127_, _00444_);
  nor (_06316_, _06315_, _06314_);
  and (_06317_, _06316_, _06313_);
  and (_06318_, _06148_, _00403_);
  and (_06319_, _06145_, _00085_);
  nor (_06320_, _06319_, _06318_);
  and (_06321_, _06125_, _00578_);
  and (_06322_, _06134_, _00485_);
  nor (_06323_, _06322_, _06321_);
  and (_06324_, _06323_, _06320_);
  and (_06325_, _06324_, _06317_);
  and (_06326_, _06325_, _06310_);
  nor (_06327_, _06326_, _06187_);
  not (_06328_, _06292_);
  and (_06329_, _06328_, _06187_);
  nor (_06330_, _06329_, _06327_);
  and (_06331_, _06240_, _05894_);
  and (_06332_, _06240_, _05899_);
  nor (_06333_, _06332_, _06331_);
  not (_06334_, _06333_);
  and (_06335_, _06334_, _06330_);
  not (_06336_, _05968_);
  not (_06337_, _05946_);
  and (_06338_, _05967_, _06337_);
  and (_06339_, _06239_, _06192_);
  and (_06340_, _06337_, _06339_);
  nor (_06341_, _06340_, _06338_);
  and (_06342_, _06240_, _05906_);
  nor (_06343_, _06342_, _06199_);
  and (_06344_, _06256_, _06337_);
  not (_06345_, _06344_);
  not (_06346_, _05618_);
  and (_06347_, _05657_, _06346_);
  and (_06348_, _06347_, _06197_);
  and (_06349_, _05964_, _06192_);
  or (_06350_, _06349_, _06348_);
  and (_06351_, _06350_, _06337_);
  and (_06352_, _05933_, _06192_);
  and (_06353_, _06352_, _06337_);
  or (_06354_, _06353_, _06251_);
  nor (_06355_, _06354_, _06351_);
  and (_06356_, _06355_, _06345_);
  and (_06357_, _06197_, _06192_);
  and (_06358_, _06347_, _05730_);
  nor (_06359_, _06358_, _06357_);
  nor (_06360_, _06359_, _05946_);
  and (_06361_, _05964_, _06347_);
  and (_06362_, _06361_, _06337_);
  nor (_06363_, _06362_, _06360_);
  and (_06364_, _06363_, _06356_);
  not (_06365_, _05918_);
  and (_06366_, _05934_, _06365_);
  and (_06367_, _05934_, _05888_);
  nor (_06368_, _06367_, _06366_);
  and (_06369_, _05969_, _06198_);
  not (_06370_, _06369_);
  and (_06371_, _05967_, _05894_);
  and (_06372_, _05966_, _06197_);
  and (_06373_, _06372_, _06337_);
  nor (_06374_, _06373_, _06371_);
  and (_06375_, _06374_, _06370_);
  and (_06376_, _06375_, _06368_);
  and (_06377_, _06259_, _06198_);
  and (_06378_, _06240_, _05911_);
  nor (_06379_, _06378_, _06377_);
  not (_06380_, _05915_);
  and (_06381_, _06380_, _06198_);
  not (_06382_, _05921_);
  and (_06383_, _05934_, _06382_);
  nor (_06384_, _06383_, _06381_);
  and (_06385_, _06384_, _06379_);
  and (_06386_, _06385_, _06376_);
  and (_06387_, _06386_, _06364_);
  and (_06388_, _06387_, _06343_);
  and (_06389_, _06388_, _06341_);
  and (_06390_, _06389_, _06024_);
  nor (_06391_, _06389_, _06019_);
  nor (_06392_, _06391_, _06390_);
  nor (_06393_, _06389_, _06095_);
  and (_06394_, _06389_, _06071_);
  nor (_06395_, _06394_, _06393_);
  nor (_06396_, _06395_, _06392_);
  and (_06397_, _06389_, _05557_);
  nor (_06398_, _06397_, _05550_);
  and (_06399_, _06397_, _05550_);
  nor (_06400_, _06399_, _06398_);
  nor (_06401_, _06389_, _05557_);
  or (_06402_, _06401_, _06397_);
  and (_06403_, _06402_, _06400_);
  and (_06404_, _06403_, _06396_);
  and (_06405_, _06404_, _00735_);
  and (_06406_, _06395_, _06392_);
  and (_06407_, _06406_, _06403_);
  and (_06408_, _06407_, _00224_);
  nor (_06409_, _06408_, _06405_);
  not (_06410_, _06402_);
  and (_06411_, _06410_, _06400_);
  and (_06412_, _06411_, _06396_);
  and (_06413_, _06412_, _00694_);
  nor (_06414_, _06410_, _06400_);
  not (_06415_, _06392_);
  nor (_06416_, _06395_, _06415_);
  and (_06417_, _06416_, _06414_);
  and (_06418_, _06417_, _00470_);
  nor (_06419_, _06418_, _06413_);
  and (_06420_, _06419_, _06409_);
  and (_06421_, _06416_, _06403_);
  and (_06422_, _06421_, _00554_);
  and (_06423_, _06395_, _06415_);
  and (_06424_, _06423_, _06403_);
  and (_06425_, _06424_, _00388_);
  nor (_06426_, _06425_, _06422_);
  and (_06427_, _06423_, _06411_);
  and (_06428_, _06427_, _00347_);
  and (_06429_, _06406_, _06414_);
  and (_06430_, _06429_, _00111_);
  nor (_06431_, _06430_, _06428_);
  and (_06432_, _06431_, _06426_);
  and (_06433_, _06432_, _06420_);
  and (_06434_, _06414_, _06396_);
  and (_06435_, _06434_, _00653_);
  nor (_06436_, _06402_, _06400_);
  and (_06437_, _06436_, _06396_);
  and (_06438_, _06437_, _00612_);
  nor (_06439_, _06438_, _06435_);
  and (_06440_, _06436_, _06416_);
  and (_06441_, _06440_, _00429_);
  and (_06442_, _06423_, _06436_);
  and (_06443_, _06442_, _00265_);
  nor (_06444_, _06443_, _06441_);
  and (_06445_, _06444_, _06439_);
  and (_06446_, _06416_, _06411_);
  and (_06447_, _06446_, _00511_);
  and (_06448_, _06406_, _06411_);
  and (_06449_, _06448_, _00171_);
  nor (_06450_, _06449_, _06447_);
  and (_06451_, _06423_, _06414_);
  and (_06452_, _06451_, _00306_);
  and (_06453_, _06406_, _06436_);
  and (_06454_, _06453_, _00070_);
  nor (_06455_, _06454_, _06452_);
  and (_06456_, _06455_, _06450_);
  and (_06457_, _06456_, _06445_);
  and (_06458_, _06457_, _06433_);
  nor (_06459_, _06458_, _06336_);
  and (_06460_, _06337_, _06198_);
  and (_06461_, _06240_, _06337_);
  nor (_06462_, _06461_, _06460_);
  nor (_06463_, _06338_, _06247_);
  not (_06464_, _06463_);
  and (_06465_, _06464_, _06292_);
  and (_06466_, _05967_, _06246_);
  and (_06467_, _06466_, _06292_);
  and (_06468_, _06250_, _06198_);
  and (_06469_, _06468_, \oc8051_golden_model_1.SP [3]);
  nor (_06470_, _06469_, _06466_);
  not (_06471_, _05954_);
  and (_06472_, _05967_, _06471_);
  nor (_06473_, _06472_, _06251_);
  or (_06474_, _06473_, _06292_);
  and (_06475_, _06240_, _06250_);
  not (_06476_, _06475_);
  nand (_06477_, _06473_, \oc8051_golden_model_1.PSW [3]);
  and (_06478_, _06477_, _06476_);
  and (_06479_, _06478_, _06474_);
  or (_06480_, _06479_, _06468_);
  and (_06481_, _06480_, _06470_);
  or (_06482_, _06481_, _06467_);
  and (_06483_, _06240_, _06246_);
  not (_06484_, _06483_);
  and (_06485_, _06463_, _06484_);
  and (_06486_, _06485_, _06482_);
  or (_06487_, _06486_, _06465_);
  and (_06488_, _06487_, _06462_);
  and (_06489_, _06192_, _05694_);
  not (_06490_, _05957_);
  and (_06491_, _06490_, _06489_);
  not (_06492_, _06491_);
  and (_06493_, _06490_, _06347_);
  and (_06494_, _06192_, _05932_);
  and (_06495_, _06494_, _06490_);
  nor (_06496_, _06495_, _06493_);
  and (_06497_, _06496_, _06492_);
  not (_06498_, _06497_);
  nor (_06499_, _06475_, _06483_);
  nand (_06500_, _06499_, _06462_);
  and (_06501_, _06500_, _06330_);
  or (_06502_, _06501_, _06498_);
  or (_06503_, _06502_, _06488_);
  and (_06504_, _06490_, _06198_);
  and (_06505_, _06240_, _06490_);
  nor (_06506_, _06505_, _06504_);
  or (_06507_, _06497_, _06292_);
  and (_06508_, _06507_, _06506_);
  and (_06509_, _06508_, _06503_);
  and (_06510_, _05969_, _05967_);
  not (_06511_, _06506_);
  and (_06512_, _06511_, _06330_);
  nor (_06513_, _06512_, _06510_);
  not (_06514_, _06513_);
  nor (_06515_, _06514_, _06509_);
  not (_06516_, _06510_);
  nor (_06517_, _06516_, _06292_);
  or (_06518_, _06517_, _06515_);
  and (_06519_, _06518_, _06242_);
  nor (_06520_, _06330_, _06242_);
  or (_06521_, _06520_, _06519_);
  and (_06522_, _06521_, _06336_);
  or (_06523_, _06522_, _06334_);
  nor (_06524_, _06523_, _06459_);
  or (_06525_, _06524_, _06335_);
  and (_06526_, _05967_, _06382_);
  not (_06527_, _06526_);
  and (_06528_, _06240_, _06382_);
  nor (_06529_, _06528_, _06383_);
  and (_06530_, _06529_, _06527_);
  and (_06531_, _05967_, _05888_);
  not (_06532_, _06531_);
  and (_06533_, _06240_, _05888_);
  nor (_06534_, _06533_, _06367_);
  and (_06535_, _06534_, _06532_);
  and (_06536_, _06535_, _06530_);
  and (_06537_, _05967_, _06380_);
  not (_06538_, _06537_);
  and (_06539_, _05967_, _06365_);
  not (_06540_, _06539_);
  and (_06541_, _06240_, _06365_);
  nor (_06542_, _06541_, _06366_);
  and (_06543_, _06542_, _06540_);
  and (_06544_, _06543_, _06538_);
  and (_06545_, _06544_, _06536_);
  nand (_06546_, _06545_, _06525_);
  and (_06547_, _06240_, _06380_);
  nor (_06548_, _06545_, _06328_);
  nor (_06549_, _06548_, _06547_);
  and (_06550_, _06549_, _06546_);
  and (_06551_, _06547_, \oc8051_golden_model_1.SP [3]);
  or (_06552_, _06551_, _06381_);
  nor (_06553_, _06552_, _06550_);
  and (_06554_, _06330_, _06381_);
  or (_06555_, _06554_, _06553_);
  and (_06556_, _06555_, _06295_);
  or (_06557_, _06556_, _06294_);
  nand (_06558_, _06557_, _06261_);
  not (_06559_, \oc8051_golden_model_1.SP [3]);
  and (_06560_, _06260_, _06559_);
  nor (_06561_, _06560_, _06377_);
  nand (_06562_, _06561_, _06558_);
  and (_06563_, _05967_, _05911_);
  not (_06564_, _06377_);
  nor (_06565_, _06564_, _06330_);
  nor (_06566_, _06565_, _06563_);
  nand (_06567_, _06566_, _06562_);
  and (_06568_, _06563_, _06292_);
  nor (_06569_, _06568_, _06199_);
  and (_06570_, _06569_, _06567_);
  not (_06571_, _06199_);
  nor (_06572_, _06330_, _06571_);
  or (_06573_, _06572_, _06570_);
  nand (_06574_, _06573_, _06189_);
  nor (_06575_, _06189_, _06292_);
  not (_06576_, _06575_);
  and (_06577_, _06576_, _06574_);
  and (_06578_, _06137_, _00745_);
  and (_06579_, _06110_, _00704_);
  nor (_06580_, _06579_, _06578_);
  and (_06581_, _06139_, _00663_);
  and (_06582_, _06125_, _00570_);
  nor (_06583_, _06582_, _06581_);
  and (_06584_, _06583_, _06580_);
  and (_06585_, _06148_, _00398_);
  and (_06586_, _06113_, _00357_);
  nor (_06587_, _06586_, _06585_);
  and (_06588_, _06121_, _00275_);
  and (_06589_, _06104_, _00193_);
  nor (_06590_, _06589_, _06588_);
  and (_06591_, _06590_, _06587_);
  and (_06592_, _06591_, _06584_);
  and (_06593_, _06134_, _00480_);
  and (_06594_, _06099_, _00121_);
  nor (_06595_, _06594_, _06593_);
  and (_06596_, _06127_, _00439_);
  and (_06597_, _06118_, _00234_);
  nor (_06598_, _06597_, _06596_);
  and (_06599_, _06598_, _06595_);
  and (_06600_, _06132_, _00622_);
  and (_06601_, _06145_, _00080_);
  nor (_06602_, _06601_, _06600_);
  and (_06603_, _06143_, _00521_);
  and (_06604_, _06150_, _00316_);
  nor (_06605_, _06604_, _06603_);
  and (_06606_, _06605_, _06602_);
  and (_06607_, _06606_, _06599_);
  and (_06608_, _06607_, _06592_);
  nor (_06609_, _06608_, _06187_);
  nor (_06610_, _06381_, _06241_);
  and (_06611_, _06610_, _06499_);
  and (_06612_, _06506_, _06462_);
  nor (_06614_, _06377_, _06199_);
  and (_06615_, _06614_, _06333_);
  and (_06616_, _06615_, _06612_);
  and (_06617_, _06616_, _06611_);
  not (_06618_, _06617_);
  and (_06619_, _06618_, _06609_);
  not (_06620_, _06619_);
  and (_06621_, _06412_, _00689_);
  and (_06622_, _06434_, _00648_);
  nor (_06623_, _06622_, _06621_);
  and (_06624_, _06424_, _00383_);
  and (_06625_, _06407_, _00219_);
  nor (_06626_, _06625_, _06624_);
  and (_06627_, _06626_, _06623_);
  and (_06628_, _06427_, _00342_);
  and (_06629_, _06442_, _00260_);
  nor (_06630_, _06629_, _06628_);
  and (_06631_, _06451_, _00301_);
  and (_06632_, _06453_, _00065_);
  nor (_06633_, _06632_, _06631_);
  and (_06634_, _06633_, _06630_);
  and (_06635_, _06634_, _06627_);
  and (_06636_, _06446_, _00506_);
  and (_06637_, _06440_, _00424_);
  nor (_06638_, _06637_, _06636_);
  and (_06639_, _06404_, _00730_);
  and (_06640_, _06437_, _00607_);
  nor (_06641_, _06640_, _06639_);
  and (_06642_, _06641_, _06638_);
  and (_06643_, _06448_, _00160_);
  and (_06644_, _06429_, _00106_);
  nor (_06645_, _06644_, _06643_);
  and (_06646_, _06421_, _00547_);
  and (_06647_, _06417_, _00465_);
  nor (_06648_, _06647_, _06646_);
  and (_06649_, _06648_, _06645_);
  and (_06650_, _06649_, _06642_);
  and (_06651_, _06650_, _06635_);
  nor (_06652_, _06651_, _06336_);
  and (_06653_, _06194_, _06380_);
  and (_06654_, _06382_, _06192_);
  nor (_06655_, _06654_, _06653_);
  and (_06656_, _05899_, _06357_);
  and (_06657_, _06194_, _06337_);
  nor (_06658_, _06657_, _06656_);
  and (_06659_, _06658_, _06655_);
  and (_06660_, _06194_, _05911_);
  and (_06661_, _06194_, _06259_);
  nor (_06662_, _06661_, _06660_);
  and (_06663_, _06194_, _06365_);
  and (_06664_, _05730_, _06192_);
  not (_06665_, _06664_);
  nor (_06666_, _06665_, _05915_);
  nor (_06667_, _06666_, _06663_);
  and (_06668_, _06667_, _06662_);
  and (_06669_, _06668_, _06659_);
  not (_06670_, \oc8051_golden_model_1.SP [2]);
  nor (_06671_, _06468_, _06260_);
  nor (_06672_, _06671_, _06670_);
  nor (_06673_, _05898_, _05896_);
  and (_06674_, _06673_, _06349_);
  not (_06675_, _06674_);
  and (_06676_, _05969_, _06357_);
  and (_06677_, _06471_, _06357_);
  nor (_06678_, _06677_, _06676_);
  and (_06679_, _06678_, _06675_);
  not (_06680_, _06679_);
  nor (_06681_, _06680_, _06672_);
  and (_06682_, _06681_, _06669_);
  and (_06683_, _06664_, _05888_);
  nor (_06684_, _06665_, _05923_);
  nor (_06685_, _06684_, _06683_);
  and (_06686_, _06664_, _05899_);
  and (_06687_, _06664_, _05906_);
  nor (_06688_, _06687_, _06686_);
  and (_06689_, _06688_, _06685_);
  and (_06690_, _06664_, _05911_);
  and (_06691_, _06664_, _06246_);
  nor (_06692_, _06691_, _06690_);
  and (_06693_, _06194_, _06246_);
  and (_06694_, _06194_, _06250_);
  nor (_06695_, _06694_, _06693_);
  and (_06696_, _06695_, _06692_);
  and (_06697_, _05888_, _06357_);
  and (_06698_, _06349_, _05888_);
  nor (_06699_, _06698_, _06697_);
  and (_06700_, _06699_, _06196_);
  and (_06701_, _06700_, _06696_);
  and (_06702_, _05954_, _05918_);
  nor (_06703_, _06702_, _06665_);
  not (_06704_, _06703_);
  and (_06705_, _06349_, _06471_);
  and (_06706_, _06664_, _06250_);
  nor (_06707_, _06706_, _06705_);
  and (_06708_, _06707_, _06704_);
  and (_06709_, _06547_, \oc8051_golden_model_1.SP [2]);
  not (_06710_, _05969_);
  and (_06711_, _06710_, _05946_);
  nor (_06712_, _06711_, _06665_);
  nor (_06713_, _06712_, _06709_);
  and (_06714_, _06713_, _06708_);
  and (_06715_, _06714_, _06701_);
  and (_06716_, _06715_, _06689_);
  and (_06717_, _06716_, _06682_);
  not (_06718_, _06717_);
  nor (_06719_, _06718_, _06652_);
  and (_06720_, _06132_, _00607_);
  and (_06721_, _06148_, _00383_);
  nor (_06722_, _06721_, _06720_);
  and (_06723_, _06113_, _00342_);
  and (_06724_, _06145_, _00065_);
  nor (_06725_, _06724_, _06723_);
  and (_06726_, _06725_, _06722_);
  and (_06727_, _06134_, _00465_);
  and (_06728_, _06143_, _00506_);
  nor (_06729_, _06728_, _06727_);
  and (_06730_, _06125_, _00547_);
  and (_06731_, _06118_, _00219_);
  nor (_06732_, _06731_, _06730_);
  and (_06733_, _06732_, _06729_);
  and (_06734_, _06733_, _06726_);
  and (_06735_, _06150_, _00301_);
  and (_06736_, _06121_, _00260_);
  nor (_06737_, _06736_, _06735_);
  and (_06738_, _06110_, _00689_);
  and (_06739_, _06099_, _00106_);
  nor (_06740_, _06739_, _06738_);
  and (_06741_, _06740_, _06737_);
  and (_06742_, _06137_, _00730_);
  and (_06743_, _06104_, _00160_);
  nor (_06744_, _06743_, _06742_);
  and (_06745_, _06139_, _00648_);
  and (_06746_, _06127_, _00424_);
  nor (_06747_, _06746_, _06745_);
  and (_06748_, _06747_, _06744_);
  and (_06749_, _06748_, _06741_);
  and (_06750_, _06749_, _06734_);
  not (_06751_, _06750_);
  nor (_06752_, _06510_, _06466_);
  and (_06753_, _06752_, _06463_);
  and (_06754_, _06753_, _06473_);
  nand (_06755_, _06754_, _06497_);
  nor (_06756_, _06563_, _06188_);
  and (_06757_, _06756_, _06295_);
  nand (_06758_, _06757_, _06545_);
  or (_06759_, _06758_, _06755_);
  and (_06760_, _06759_, _06751_);
  not (_06761_, _06760_);
  and (_06762_, _06761_, _06719_);
  and (_06763_, _06762_, _06620_);
  not (_06764_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_06765_, _06292_, _06187_);
  nor (_06766_, _06765_, _06571_);
  nor (_06767_, _06242_, _06765_);
  nor (_06768_, _06506_, _06765_);
  nand (_06769_, _06125_, _00537_);
  nand (_06770_, _06143_, _00496_);
  and (_06771_, _06770_, _06769_);
  nand (_06772_, _06148_, _00373_);
  nand (_06773_, _06113_, _00332_);
  and (_06774_, _06773_, _06772_);
  and (_06775_, _06774_, _06771_);
  nand (_06776_, _06137_, _00720_);
  nand (_06777_, _06110_, _00679_);
  and (_06778_, _06777_, _06776_);
  nand (_06779_, _06118_, _00209_);
  nand (_06780_, _06104_, _00138_);
  and (_06781_, _06780_, _06779_);
  and (_06782_, _06781_, _06778_);
  and (_06783_, _06782_, _06775_);
  nand (_06784_, _06139_, _00638_);
  nand (_06785_, _06132_, _00596_);
  and (_06786_, _06785_, _06784_);
  nand (_06787_, _06145_, _00055_);
  nand (_06788_, _06099_, _00096_);
  and (_06789_, _06788_, _06787_);
  and (_06790_, _06789_, _06786_);
  nand (_06791_, _06134_, _00455_);
  nand (_06792_, _06127_, _00414_);
  and (_06793_, _06792_, _06791_);
  nand (_06794_, _06150_, _00291_);
  nand (_06795_, _06121_, _00250_);
  and (_06796_, _06795_, _06794_);
  and (_06797_, _06796_, _06793_);
  and (_06798_, _06797_, _06790_);
  nand (_06799_, _06798_, _06783_);
  and (_06800_, _06799_, _06338_);
  not (_06801_, _06466_);
  and (_06802_, _06798_, _06783_);
  or (_06803_, _06802_, _06801_);
  and (_06804_, _06799_, _06251_);
  and (_06805_, _06347_, _05694_);
  and (_06806_, _06471_, _06805_);
  not (_06807_, _06806_);
  and (_06808_, _06471_, _06339_);
  nor (_06809_, _06808_, _06677_);
  and (_06810_, _05966_, _06239_);
  and (_06811_, _06810_, _06471_);
  and (_06812_, _06810_, _06255_);
  nor (_06813_, _06812_, _06811_);
  and (_06814_, _06813_, _06809_);
  and (_06815_, _06814_, _06807_);
  and (_06816_, _06250_, _06339_);
  and (_06817_, _06347_, _06239_);
  not (_06818_, _06817_);
  nor (_06819_, _06810_, _06348_);
  nor (_06820_, _05967_, _06357_);
  and (_06821_, _06820_, _06819_);
  and (_06822_, _06821_, _06818_);
  nor (_06823_, _06822_, _05949_);
  nor (_06824_, _06823_, _06816_);
  and (_06825_, _06824_, _06815_);
  or (_06826_, _06825_, _06804_);
  nand (_06827_, _06802_, _06472_);
  and (_06828_, _06827_, _06476_);
  nand (_06829_, _06828_, _06826_);
  or (_06830_, _06476_, _06765_);
  nand (_06831_, _06830_, _06829_);
  and (_06832_, _06246_, _06358_);
  or (_06833_, _06693_, _06691_);
  or (_06834_, _06833_, _06832_);
  and (_06835_, _06834_, _05694_);
  not (_06836_, _06835_);
  and (_06837_, _06468_, _06235_);
  nor (_06838_, _06837_, _06466_);
  and (_06839_, _06810_, _06246_);
  and (_06840_, _06246_, _06348_);
  nor (_06841_, _06840_, _06839_);
  and (_06842_, _06841_, _06838_);
  and (_06843_, _06842_, _06836_);
  nand (_06844_, _06843_, _06831_);
  nand (_06845_, _06844_, _06803_);
  and (_06846_, _06845_, _06484_);
  nor (_06847_, _06484_, _06765_);
  or (_06848_, _06847_, _06846_);
  and (_06849_, _06802_, _06247_);
  not (_06850_, _06341_);
  not (_06851_, _06357_);
  and (_06852_, _06819_, _06818_);
  and (_06853_, _06852_, _06851_);
  nor (_06854_, _06853_, _05946_);
  nor (_06855_, _06854_, _06850_);
  not (_06856_, _06855_);
  nor (_06857_, _06856_, _06849_);
  and (_06858_, _06857_, _06848_);
  or (_06859_, _06858_, _06800_);
  nand (_06860_, _06859_, _06462_);
  nor (_06861_, _06462_, _06765_);
  nor (_06862_, _06861_, _06498_);
  nand (_06863_, _06862_, _06860_);
  and (_06864_, _06802_, _06498_);
  and (_06865_, _06810_, _06490_);
  nor (_06866_, _06865_, _06511_);
  not (_06867_, _06866_);
  nor (_06868_, _06867_, _06864_);
  and (_06869_, _06868_, _06863_);
  nor (_06870_, _06869_, _06768_);
  not (_06871_, _06339_);
  and (_06872_, _06822_, _06871_);
  nor (_06873_, _06872_, _06710_);
  nor (_06874_, _06873_, _06870_);
  and (_06875_, _06799_, _06510_);
  or (_06876_, _06875_, _06874_);
  and (_06877_, _06876_, _06242_);
  nor (_06878_, _06877_, _06767_);
  not (_06879_, _05899_);
  nor (_06880_, _06872_, _06879_);
  nor (_06881_, _06880_, _06878_);
  and (_06882_, _06404_, _00720_);
  and (_06883_, _06407_, _00209_);
  nor (_06884_, _06883_, _06882_);
  and (_06885_, _06412_, _00679_);
  and (_06886_, _06440_, _00414_);
  nor (_06887_, _06886_, _06885_);
  and (_06888_, _06887_, _06884_);
  and (_06889_, _06421_, _00537_);
  and (_06890_, _06424_, _00373_);
  nor (_06891_, _06890_, _06889_);
  and (_06892_, _06427_, _00332_);
  and (_06893_, _06429_, _00096_);
  nor (_06894_, _06893_, _06892_);
  and (_06895_, _06894_, _06891_);
  and (_06896_, _06895_, _06888_);
  and (_06897_, _06434_, _00638_);
  and (_06898_, _06437_, _00596_);
  nor (_06899_, _06898_, _06897_);
  and (_06900_, _06417_, _00455_);
  and (_06901_, _06448_, _00138_);
  nor (_06902_, _06901_, _06900_);
  and (_06903_, _06902_, _06899_);
  and (_06904_, _06446_, _00496_);
  and (_06905_, _06442_, _00250_);
  nor (_06906_, _06905_, _06904_);
  and (_06907_, _06451_, _00291_);
  and (_06908_, _06453_, _00055_);
  nor (_06909_, _06908_, _06907_);
  and (_06910_, _06909_, _06906_);
  and (_06911_, _06910_, _06903_);
  and (_06912_, _06911_, _06896_);
  nor (_06913_, _06912_, _06336_);
  or (_06914_, _06913_, _06881_);
  and (_06915_, _06332_, _06765_);
  and (_06916_, _06810_, _05894_);
  nor (_06917_, _06916_, _06331_);
  not (_06918_, _06917_);
  nor (_06919_, _06918_, _06915_);
  and (_06920_, _06919_, _06914_);
  not (_06921_, _06331_);
  nor (_06922_, _06921_, _06765_);
  nor (_06923_, _06922_, _06920_);
  not (_06924_, _05888_);
  not (_06925_, _06489_);
  and (_06926_, _06852_, _06925_);
  nor (_06927_, _06926_, _06924_);
  nor (_06928_, _06927_, _06923_);
  nor (_06929_, _06799_, _06535_);
  nor (_06930_, _06926_, _05918_);
  nor (_06931_, _06930_, _06929_);
  and (_06932_, _06931_, _06928_);
  nor (_06933_, _06799_, _06543_);
  nor (_06934_, _06926_, _05921_);
  nor (_06935_, _06934_, _06933_);
  and (_06936_, _06935_, _06932_);
  nor (_06937_, _06799_, _06530_);
  nor (_06938_, _06872_, _05915_);
  nor (_06939_, _06938_, _06937_);
  and (_06940_, _06939_, _06936_);
  and (_06941_, _06799_, _06537_);
  or (_06942_, _06941_, _06940_);
  and (_06943_, _06547_, _06235_);
  nor (_06944_, _06943_, _06381_);
  and (_06945_, _06944_, _06942_);
  not (_06946_, _06381_);
  nor (_06947_, _06946_, _06765_);
  nor (_06948_, _06947_, _06945_);
  nor (_06949_, _06872_, _05923_);
  nor (_06950_, _06949_, _06948_);
  and (_06951_, _06799_, _06293_);
  or (_06952_, _06951_, _06950_);
  and (_06953_, _06260_, _06235_);
  nor (_06954_, _06953_, _06377_);
  and (_06955_, _06954_, _06952_);
  nor (_06956_, _06564_, _06765_);
  or (_06957_, _06956_, _06955_);
  and (_06958_, _05911_, _06339_);
  not (_06959_, _06958_);
  and (_06960_, _05911_, _06357_);
  and (_06961_, _05911_, _06805_);
  nor (_06962_, _06961_, _06960_);
  and (_06963_, _06810_, _05911_);
  nor (_06964_, _06963_, _06563_);
  and (_06965_, _06964_, _06962_);
  and (_06966_, _06965_, _06959_);
  and (_06967_, _06966_, _06957_);
  and (_06968_, _06799_, _06563_);
  or (_06969_, _06968_, _06967_);
  and (_06970_, _06969_, _06571_);
  or (_06971_, _06970_, _06766_);
  nand (_06972_, _05657_, _05694_);
  not (_06973_, _06972_);
  and (_06974_, _06973_, _05906_);
  not (_06975_, _06974_);
  and (_06976_, _06810_, _05906_);
  nor (_06977_, _06976_, _06188_);
  and (_06978_, _06977_, _06975_);
  nand (_06979_, _06978_, _06971_);
  and (_06980_, _06799_, _06188_);
  not (_06981_, _06980_);
  nand (_06982_, _06981_, _06979_);
  or (_06983_, _06982_, _06764_);
  and (_06984_, _06231_, _06618_);
  not (_06985_, _06984_);
  and (_06986_, _06156_, _06759_);
  not (_06987_, _06986_);
  and (_06988_, _06429_, _00101_);
  and (_06989_, _06448_, _00149_);
  nor (_06990_, _06989_, _06988_);
  and (_06991_, _06437_, _00602_);
  and (_06992_, _06427_, _00337_);
  nor (_06993_, _06992_, _06991_);
  and (_06994_, _06993_, _06990_);
  and (_06995_, _06421_, _00542_);
  and (_06996_, _06417_, _00460_);
  nor (_06997_, _06996_, _06995_);
  and (_06998_, _06451_, _00296_);
  and (_06999_, _06453_, _00060_);
  nor (_07000_, _06999_, _06998_);
  and (_07001_, _07000_, _06997_);
  and (_07002_, _07001_, _06994_);
  and (_07003_, _06404_, _00725_);
  and (_07004_, _06412_, _00684_);
  nor (_07005_, _07004_, _07003_);
  and (_07006_, _06434_, _00643_);
  and (_07007_, _06440_, _00419_);
  nor (_07008_, _07007_, _07006_);
  and (_07009_, _07008_, _07005_);
  and (_07010_, _06446_, _00501_);
  and (_07011_, _06407_, _00214_);
  nor (_07012_, _07011_, _07010_);
  and (_07013_, _06424_, _00378_);
  and (_07014_, _06442_, _00255_);
  nor (_07015_, _07014_, _07013_);
  and (_07016_, _07015_, _07012_);
  and (_07017_, _07016_, _07009_);
  and (_07018_, _07017_, _07002_);
  nor (_07019_, _07018_, _06336_);
  and (_07020_, _06382_, _06358_);
  and (_07021_, _06250_, _06358_);
  nor (_07022_, _07021_, _07020_);
  nor (_07023_, _06706_, _06666_);
  and (_07024_, _07023_, _07022_);
  and (_07025_, _06704_, _06692_);
  and (_07026_, _07025_, _07024_);
  nor (_07027_, _06547_, _06260_);
  nor (_07028_, _07027_, _06233_);
  not (_07029_, _07028_);
  and (_07030_, _05899_, _06358_);
  not (_07031_, _07030_);
  nor (_07032_, _06665_, _05921_);
  and (_07033_, _06365_, _06358_);
  nor (_07034_, _07033_, _07032_);
  and (_07035_, _07034_, _07031_);
  and (_07036_, _07035_, _07029_);
  and (_07037_, _07036_, _07026_);
  and (_07038_, _06711_, _06924_);
  nor (_07039_, _06712_, _06358_);
  nor (_07040_, _07039_, _07038_);
  not (_07041_, _07040_);
  and (_07042_, _06468_, \oc8051_golden_model_1.SP [1]);
  not (_07043_, _06358_);
  and (_07044_, _05952_, _05923_);
  nor (_07045_, _07044_, _07043_);
  nor (_07046_, _07045_, _07042_);
  and (_07047_, _05954_, _05915_);
  nor (_07048_, _07047_, _07043_);
  not (_07049_, _07048_);
  and (_07050_, _05911_, _06358_);
  not (_07051_, _07050_);
  and (_07052_, _06817_, _05906_);
  and (_07053_, _05933_, _06347_);
  and (_07054_, _07053_, _05906_);
  nor (_07055_, _07054_, _07052_);
  and (_07056_, _07055_, _07051_);
  and (_07057_, _07056_, _07049_);
  and (_07058_, _07057_, _07046_);
  and (_07059_, _07058_, _06689_);
  and (_07060_, _07059_, _07041_);
  and (_07061_, _07060_, _07037_);
  not (_07062_, _07061_);
  nor (_07063_, _07062_, _07019_);
  and (_07064_, _07063_, _06987_);
  and (_07065_, _07064_, _06985_);
  not (_07066_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_07067_, _06981_, _06979_);
  or (_07068_, _07067_, _07066_);
  and (_07069_, _07068_, _07065_);
  nand (_07070_, _07069_, _06983_);
  not (_07071_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_07072_, _07067_, _07071_);
  not (_07073_, _07065_);
  not (_07074_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_07075_, _06982_, _07074_);
  and (_07076_, _07075_, _07073_);
  nand (_07077_, _07076_, _07072_);
  nand (_07078_, _07077_, _07070_);
  nand (_07079_, _07078_, _06763_);
  not (_07080_, _06763_);
  not (_07081_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_07082_, _07067_, _07081_);
  not (_07083_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_07084_, _06982_, _07083_);
  and (_07085_, _07084_, _07073_);
  nand (_07086_, _07085_, _07082_);
  not (_07087_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_07088_, _06982_, _07087_);
  not (_07089_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_07090_, _07067_, _07089_);
  and (_07091_, _07090_, _07065_);
  nand (_07092_, _07091_, _07088_);
  nand (_07093_, _07092_, _07086_);
  nand (_07094_, _07093_, _07080_);
  nand (_07095_, _07094_, _07079_);
  nand (_07096_, _07095_, _06577_);
  not (_07097_, _06577_);
  nand (_07098_, _06982_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_07099_, _07067_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_07100_, _07099_, _07073_);
  nand (_07101_, _07100_, _07098_);
  nand (_07102_, _07067_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_07103_, _06982_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_07104_, _07103_, _07065_);
  nand (_07105_, _07104_, _07102_);
  nand (_07106_, _07105_, _07101_);
  nand (_07107_, _07106_, _06763_);
  nand (_07108_, _06982_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_07109_, _07067_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_07110_, _07109_, _07073_);
  nand (_07111_, _07110_, _07108_);
  nand (_07112_, _07067_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_07113_, _06982_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_07114_, _07113_, _07065_);
  nand (_07115_, _07114_, _07112_);
  nand (_07116_, _07115_, _07111_);
  nand (_07117_, _07116_, _07080_);
  nand (_07118_, _07117_, _07107_);
  nand (_07119_, _07118_, _07097_);
  nand (_07120_, _07119_, _07096_);
  and (_07121_, _07120_, _06258_);
  or (_07122_, _07121_, _06257_);
  and (_07123_, _06352_, _06471_);
  not (_07124_, _07123_);
  nor (_07125_, _07124_, _06187_);
  and (_07126_, _07125_, _06155_);
  or (_07127_, _07126_, _07122_);
  and (_07128_, _06237_, _06705_);
  and (_07129_, _06347_, _06193_);
  and (_07130_, _07129_, _06250_);
  or (_07131_, _07130_, _06694_);
  or (_07132_, _07131_, _07128_);
  or (_07133_, _07132_, _07127_);
  and (_07134_, _06256_, _06250_);
  and (_07135_, _07120_, _07134_);
  or (_07136_, _07135_, _06253_);
  or (_07137_, _07136_, _07133_);
  and (_07138_, _07137_, _06254_);
  nor (_07139_, _06476_, _06187_);
  and (_07140_, _06230_, _07139_);
  or (_07141_, _07140_, _07138_);
  not (_07142_, _06468_);
  nor (_07143_, _07142_, _06187_);
  nor (_07144_, _06248_, _05950_);
  or (_07145_, _07144_, _07143_);
  or (_07146_, _07145_, _07141_);
  nand (_07147_, _07143_, _06156_);
  and (_07148_, _07147_, _07146_);
  and (_07149_, _07129_, _06246_);
  or (_07150_, _07149_, _06693_);
  or (_07151_, _07150_, _07148_);
  nor (_07152_, _06801_, _06187_);
  and (_07153_, _06256_, _06246_);
  and (_07154_, _07120_, _07153_);
  or (_07155_, _07154_, _07152_);
  or (_07156_, _07155_, _07151_);
  nand (_07157_, _07152_, _06156_);
  and (_07158_, _07157_, _07156_);
  nor (_07159_, _06484_, _06187_);
  and (_07160_, _06230_, _07159_);
  or (_07161_, _07160_, _06247_);
  nor (_07162_, _07161_, _07158_);
  nor (_07163_, _07162_, _06249_);
  not (_07164_, _06461_);
  nor (_07165_, _07164_, _06187_);
  and (_07166_, _06230_, _07165_);
  or (_07167_, _07166_, _07163_);
  nor (_07168_, _06248_, _05947_);
  and (_07169_, _07129_, _06490_);
  and (_07170_, _06194_, _06490_);
  or (_07171_, _07170_, _07169_);
  or (_07172_, _07171_, _07168_);
  or (_07173_, _07172_, _07167_);
  and (_07174_, _06256_, _06490_);
  and (_07175_, _07120_, _07174_);
  or (_07176_, _07175_, _06243_);
  or (_07177_, _07176_, _07173_);
  and (_07178_, _07177_, _06245_);
  or (_07179_, _07178_, _05970_);
  nand (_07180_, _06248_, _05970_);
  and (_07181_, _07180_, _07179_);
  and (_07182_, _06256_, _05899_);
  not (_07183_, _07182_);
  nor (_07184_, _07183_, _06187_);
  not (_07185_, _07184_);
  nor (_07186_, _06187_, _06336_);
  and (_07187_, _05899_, _05657_);
  not (_07188_, _07187_);
  nor (_07189_, _07188_, _06187_);
  nor (_07190_, _07189_, _07186_);
  and (_07191_, _07190_, _07185_);
  nor (_07192_, _07191_, _06156_);
  and (_07193_, _06194_, _05894_);
  and (_07194_, _07129_, _05894_);
  or (_07195_, _07194_, _07193_);
  or (_07196_, _07195_, _07192_);
  or (_07197_, _07196_, _07181_);
  not (_07198_, _06371_);
  nor (_07199_, _07198_, _06187_);
  and (_07200_, _06256_, _05894_);
  and (_07201_, _07120_, _07200_);
  or (_07202_, _07201_, _07199_);
  or (_07203_, _07202_, _07197_);
  nand (_07204_, _07199_, _06156_);
  and (_07205_, _07204_, _07203_);
  or (_07206_, _07205_, _05895_);
  nand (_07207_, _06248_, _05895_);
  and (_07208_, _07207_, _07206_);
  not (_07209_, _05919_);
  not (_07210_, _06541_);
  nor (_07211_, _07210_, _06187_);
  not (_07212_, _07211_);
  not (_07213_, _06366_);
  nor (_07214_, _07213_, _06187_);
  not (_07215_, _07214_);
  not (_07216_, _06533_);
  nor (_07217_, _07216_, _06187_);
  not (_07218_, _06367_);
  nor (_07219_, _07218_, _06187_);
  nor (_07220_, _07219_, _07217_);
  and (_07221_, _07220_, _07215_);
  and (_07222_, _07221_, _07212_);
  nor (_07223_, _07222_, _06156_);
  or (_07224_, _07223_, _07209_);
  or (_07225_, _07224_, _07208_);
  or (_07226_, _06237_, _05919_);
  and (_07227_, _07226_, _07225_);
  not (_07228_, _05916_);
  not (_07229_, _06528_);
  nor (_07230_, _07229_, _06187_);
  not (_07231_, _06383_);
  nor (_07232_, _07231_, _06187_);
  nor (_07233_, _07232_, _07230_);
  nor (_07234_, _07233_, _06156_);
  or (_07235_, _07234_, _07228_);
  or (_07236_, _07235_, _07227_);
  and (_07237_, _07236_, _06238_);
  and (_07238_, _07129_, _05911_);
  or (_07239_, _07238_, _06660_);
  nor (_07240_, _07239_, _07237_);
  not (_07241_, _06563_);
  nor (_07242_, _07241_, _06187_);
  and (_07243_, _06256_, _05911_);
  and (_07244_, _07120_, _07243_);
  nor (_07245_, _07244_, _07242_);
  and (_07246_, _07245_, _07240_);
  and (_07247_, _07242_, _06156_);
  nor (_07248_, _07247_, _07246_);
  nor (_07249_, _06187_, _06571_);
  nor (_07250_, _06378_, _05912_);
  nor (_07251_, _06248_, _07250_);
  nor (_07252_, _07251_, _07249_);
  not (_07253_, _07252_);
  nor (_07254_, _07253_, _07248_);
  nor (_07255_, _07254_, _06232_);
  and (_07256_, _07129_, _05906_);
  nor (_07257_, _07256_, _07255_);
  and (_07258_, _07257_, _06196_);
  and (_07259_, _06256_, _05906_);
  and (_07260_, _07120_, _07259_);
  nor (_07261_, _07260_, _06190_);
  and (_07262_, _07261_, _07258_);
  nor (_07263_, _07262_, _06191_);
  not (_07264_, _07263_);
  not (_07265_, _07249_);
  nor (_07266_, _05916_, \oc8051_golden_model_1.SP [0]);
  nor (_07267_, _07191_, _06799_);
  nor (_07268_, _05947_, _06235_);
  nor (_07269_, _07164_, _06765_);
  not (_07270_, _07165_);
  and (_07271_, _06705_, _06235_);
  not (_07272_, _06705_);
  not (_07273_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_07274_, _06982_, _07273_);
  not (_07275_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_07276_, _07067_, _07275_);
  and (_07277_, _07276_, _07065_);
  nand (_07278_, _07277_, _07274_);
  not (_07279_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_07280_, _07067_, _07279_);
  not (_07281_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_07282_, _06982_, _07281_);
  and (_07283_, _07282_, _07073_);
  nand (_07284_, _07283_, _07280_);
  nand (_07285_, _07284_, _07278_);
  nand (_07286_, _07285_, _06763_);
  not (_07287_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_07288_, _07067_, _07287_);
  not (_07289_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_07290_, _06982_, _07289_);
  and (_07291_, _07290_, _07073_);
  nand (_07292_, _07291_, _07288_);
  not (_07293_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_07294_, _06982_, _07293_);
  not (_07295_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_07296_, _07067_, _07295_);
  and (_07297_, _07296_, _07065_);
  nand (_07298_, _07297_, _07294_);
  nand (_07299_, _07298_, _07292_);
  nand (_07300_, _07299_, _07080_);
  nand (_07301_, _07300_, _07286_);
  nand (_07302_, _07301_, _06577_);
  nand (_07303_, _06982_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_07304_, _07067_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_07305_, _07304_, _07073_);
  nand (_07306_, _07305_, _07303_);
  nand (_07307_, _07067_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_07308_, _06982_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_07309_, _07308_, _07065_);
  nand (_07310_, _07309_, _07307_);
  nand (_07311_, _07310_, _07306_);
  nand (_07312_, _07311_, _06763_);
  nand (_07313_, _06982_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_07314_, _07067_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_07315_, _07314_, _07073_);
  nand (_07316_, _07315_, _07313_);
  nand (_07317_, _07067_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand (_07318_, _06982_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_07319_, _07318_, _07065_);
  nand (_07320_, _07319_, _07317_);
  nand (_07321_, _07320_, _07316_);
  nand (_07322_, _07321_, _07080_);
  nand (_07323_, _07322_, _07312_);
  nand (_07324_, _07323_, _07097_);
  and (_07325_, _07324_, _07302_);
  and (_07326_, _07325_, _06258_);
  nor (_07327_, _06372_, _05733_);
  and (_07328_, _07327_, _06819_);
  nor (_07329_, _07328_, _05959_);
  not (_07330_, _07329_);
  nor (_07331_, _07330_, _07326_);
  and (_07332_, _07125_, _06802_);
  nor (_07333_, _07332_, _07331_);
  and (_07334_, _07333_, _07272_);
  nor (_07335_, _07334_, _07271_);
  nor (_07336_, _05949_, _06972_);
  nor (_07337_, _07336_, _07335_);
  not (_07338_, _07134_);
  nor (_07339_, _07338_, _07325_);
  nor (_07340_, _07339_, _06253_);
  and (_07341_, _07340_, _07337_);
  and (_07342_, _06253_, _06799_);
  nor (_07343_, _07342_, _07341_);
  nor (_07344_, _07343_, _07139_);
  not (_07345_, _07344_);
  and (_07346_, _07345_, _06830_);
  nor (_07347_, _05950_, _06235_);
  nor (_07348_, _07347_, _07346_);
  nor (_07349_, _05952_, _06972_);
  and (_07350_, _07143_, _06802_);
  nor (_07351_, _07350_, _07349_);
  and (_07352_, _07351_, _07348_);
  not (_07353_, _07153_);
  nor (_07354_, _07353_, _07325_);
  not (_07355_, _07354_);
  and (_07356_, _07355_, _07352_);
  and (_07357_, _07152_, _06802_);
  nor (_07358_, _07357_, _07159_);
  and (_07359_, _07358_, _07356_);
  nor (_07360_, _07359_, _06847_);
  nor (_07361_, _07360_, _06247_);
  and (_07362_, _06247_, _06235_);
  or (_07363_, _07362_, _07361_);
  and (_07364_, _07363_, _07270_);
  nor (_07365_, _07364_, _07269_);
  nor (_07366_, _05957_, _06972_);
  or (_07367_, _07366_, _07365_);
  nor (_07368_, _07367_, _07268_);
  not (_07369_, _07174_);
  nor (_07370_, _07369_, _07325_);
  nor (_07371_, _07370_, _06243_);
  and (_07372_, _07371_, _07368_);
  nor (_07373_, _07372_, _06767_);
  nor (_07374_, _07373_, _05970_);
  and (_07375_, _05970_, _06235_);
  nor (_07376_, _07375_, _07374_);
  and (_07377_, _05894_, _06973_);
  or (_07378_, _07377_, _07376_);
  nor (_07379_, _07378_, _07267_);
  not (_07380_, _07325_);
  and (_07381_, _07200_, _07380_);
  not (_07382_, _07381_);
  and (_07383_, _07382_, _07379_);
  and (_07384_, _07199_, _06802_);
  nor (_07385_, _07384_, _05895_);
  and (_07386_, _07385_, _07383_);
  and (_07387_, _05895_, _06235_);
  nor (_07388_, _07387_, _07386_);
  nor (_07389_, _07222_, _06799_);
  nor (_07390_, _07389_, _07209_);
  not (_07391_, _07390_);
  nor (_07392_, _07391_, _07388_);
  nor (_07393_, _05919_, \oc8051_golden_model_1.SP [0]);
  nor (_07394_, _07393_, _07392_);
  nor (_07395_, _06529_, _06187_);
  and (_07396_, _07395_, _06802_);
  or (_07397_, _07396_, _07228_);
  nor (_07398_, _07397_, _07394_);
  nor (_07399_, _07398_, _07266_);
  and (_07400_, _06962_, _06959_);
  not (_07401_, _07400_);
  nor (_07402_, _07401_, _07399_);
  not (_07403_, _07243_);
  nor (_07404_, _07403_, _07325_);
  nor (_07405_, _07404_, _07242_);
  and (_07406_, _07405_, _07402_);
  and (_07407_, _07242_, _06799_);
  nor (_07408_, _07407_, _07406_);
  nor (_07409_, _07250_, _06235_);
  nor (_07410_, _07409_, _07408_);
  and (_07411_, _07410_, _07265_);
  nor (_07412_, _07411_, _06766_);
  nor (_07413_, _07412_, _06974_);
  not (_07414_, _07259_);
  nor (_07415_, _07414_, _07325_);
  nor (_07416_, _07415_, _06190_);
  and (_07417_, _07416_, _07413_);
  and (_07418_, _06190_, _06799_);
  nor (_07419_, _07418_, _07417_);
  not (_07420_, _00000_);
  nor (_07421_, _07152_, _07143_);
  nor (_07422_, _06253_, _07139_);
  and (_07423_, _07422_, _07421_);
  nor (_07424_, _07199_, _07159_);
  nor (_07425_, _07200_, _06495_);
  and (_07426_, _07425_, _06707_);
  and (_07427_, _07250_, _05920_);
  and (_07428_, _07427_, _07426_);
  nor (_07429_, _07021_, _06840_);
  nor (_07430_, _06976_, _06832_);
  and (_07431_, _07430_, _07429_);
  nor (_07432_, _07243_, _06247_);
  and (_07433_, _06192_, _05906_);
  nor (_07434_, _07433_, _06660_);
  and (_07435_, _07434_, _07432_);
  and (_07436_, _07435_, _07431_);
  and (_07437_, _07436_, _07428_);
  and (_07438_, _05894_, _06358_);
  not (_07439_, _07438_);
  nor (_07440_, _07129_, _06256_);
  nor (_07441_, _07440_, _05959_);
  nor (_07442_, _07441_, _07169_);
  and (_07443_, _07442_, _07439_);
  and (_07444_, _06493_, _05730_);
  not (_07445_, _07444_);
  and (_07446_, _07445_, _07056_);
  and (_07447_, _07446_, _06696_);
  and (_07448_, _07447_, _07443_);
  and (_07449_, _07448_, _07437_);
  nor (_07450_, _06352_, _06361_);
  and (_07451_, _06361_, _06246_);
  nor (_07452_, _07451_, _05894_);
  nor (_07453_, _07452_, _07450_);
  not (_07454_, _07453_);
  and (_07455_, _05966_, _05933_);
  and (_07456_, _07455_, _05906_);
  nor (_07457_, _07256_, _07456_);
  and (_07458_, _06349_, _05894_);
  and (_07459_, _05894_, _06489_);
  nor (_07460_, _07459_, _07458_);
  and (_07461_, _07460_, _07457_);
  and (_07462_, _07461_, _07454_);
  not (_07463_, _07238_);
  nor (_07464_, _07130_, _06491_);
  and (_07465_, _07464_, _07463_);
  nor (_07466_, _07174_, _07153_);
  and (_07467_, _05894_, _06348_);
  nor (_07468_, _07467_, _07134_);
  and (_07469_, _07468_, _07466_);
  and (_07470_, _07469_, _07465_);
  not (_07471_, _05947_);
  or (_07472_, _05970_, _07471_);
  not (_07473_, _07472_);
  not (_07474_, _05950_);
  nor (_07475_, _07474_, _05895_);
  and (_07476_, _07475_, _07473_);
  and (_07477_, _06372_, _06255_);
  and (_07478_, _05967_, _06255_);
  nor (_07479_, _07478_, _07477_);
  nand (_07480_, _07479_, _05960_);
  not (_07481_, _07480_);
  and (_07482_, _07481_, _07476_);
  and (_07483_, _07482_, _07470_);
  and (_07484_, _07483_, _07462_);
  and (_07485_, _07484_, _07449_);
  and (_07486_, _07485_, _07212_);
  and (_07487_, _07486_, _07424_);
  and (_07488_, _07487_, _07423_);
  nor (_07489_, _07242_, _07249_);
  and (_07490_, _05899_, _06347_);
  nor (_07491_, _07490_, _06656_);
  or (_07492_, _06494_, _06339_);
  and (_07493_, _07492_, _05899_);
  not (_07494_, _07493_);
  nor (_07495_, _07182_, _07123_);
  and (_07496_, _07495_, _07494_);
  and (_07497_, _07496_, _07491_);
  nor (_07498_, _07497_, _06187_);
  nor (_07499_, _07498_, _06190_);
  and (_07500_, _07499_, _07489_);
  nor (_07501_, _07165_, _06243_);
  nor (_07502_, _07395_, _07186_);
  and (_07503_, _07502_, _07501_);
  and (_07504_, _07503_, _07500_);
  and (_07505_, _07504_, _07221_);
  and (_07506_, _07505_, _07488_);
  nor (_07507_, _07506_, _07420_);
  not (_07508_, _07507_);
  nor (_07509_, _07508_, _07419_);
  and (_07510_, _07509_, _07264_);
  and (_07511_, _06609_, _06199_);
  and (_07512_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_07513_, _07512_, \oc8051_golden_model_1.SP [2]);
  nor (_07514_, _07512_, \oc8051_golden_model_1.SP [2]);
  nor (_07515_, _07514_, _07513_);
  not (_07516_, _07515_);
  nor (_07517_, _07516_, _05916_);
  and (_07518_, _07199_, _06751_);
  nor (_07519_, _07191_, _06751_);
  and (_07520_, _05894_, _06347_);
  and (_07521_, _06609_, _06241_);
  and (_07522_, _07515_, _06247_);
  not (_07523_, _06247_);
  and (_07524_, _06609_, _06475_);
  and (_07525_, _06253_, _06751_);
  not (_07526_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_07527_, _06982_, _07526_);
  not (_07528_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_07529_, _07067_, _07528_);
  and (_07530_, _07529_, _07065_);
  nand (_07531_, _07530_, _07527_);
  not (_07532_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_07533_, _07067_, _07532_);
  not (_07534_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_07535_, _06982_, _07534_);
  and (_07536_, _07535_, _07073_);
  nand (_07537_, _07536_, _07533_);
  nand (_07538_, _07537_, _07531_);
  nand (_07539_, _07538_, _06763_);
  not (_07540_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_07541_, _07067_, _07540_);
  not (_07542_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_07543_, _06982_, _07542_);
  and (_07544_, _07543_, _07073_);
  nand (_07545_, _07544_, _07541_);
  not (_07546_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_07547_, _06982_, _07546_);
  not (_07548_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_07549_, _07067_, _07548_);
  and (_07550_, _07549_, _07065_);
  nand (_07551_, _07550_, _07547_);
  nand (_07552_, _07551_, _07545_);
  nand (_07553_, _07552_, _07080_);
  nand (_07554_, _07553_, _07539_);
  nand (_07555_, _07554_, _06577_);
  nand (_07556_, _06982_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_07557_, _07067_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_07558_, _07557_, _07073_);
  nand (_07559_, _07558_, _07556_);
  nand (_07560_, _07067_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_07561_, _06982_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_07562_, _07561_, _07065_);
  nand (_07563_, _07562_, _07560_);
  nand (_07564_, _07563_, _07559_);
  nand (_07565_, _07564_, _06763_);
  nand (_07566_, _06982_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_07567_, _07067_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_07568_, _07567_, _07073_);
  nand (_07569_, _07568_, _07566_);
  nand (_07570_, _07067_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_07571_, _06982_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_07572_, _07571_, _07065_);
  nand (_07573_, _07572_, _07570_);
  nand (_07574_, _07573_, _07569_);
  nand (_07575_, _07574_, _07080_);
  nand (_07576_, _07575_, _07565_);
  nand (_07577_, _07576_, _07097_);
  nand (_07578_, _07577_, _07555_);
  nor (_07579_, _07578_, _05960_);
  nor (_07580_, _07579_, _07481_);
  and (_07581_, _07125_, _06750_);
  or (_07582_, _07581_, _07580_);
  and (_07583_, _07516_, _06705_);
  and (_07584_, _06250_, _06347_);
  nor (_07585_, _07584_, _07583_);
  not (_07586_, _07585_);
  nor (_07587_, _07586_, _07582_);
  and (_07588_, _07578_, _07134_);
  nor (_07589_, _07588_, _06253_);
  and (_07590_, _07589_, _07587_);
  nor (_07591_, _07590_, _07525_);
  nor (_07592_, _07591_, _07139_);
  nor (_07593_, _07592_, _07524_);
  nor (_07594_, _07515_, _05950_);
  nor (_07595_, _07594_, _07593_);
  and (_07596_, _06246_, _06347_);
  and (_07597_, _07143_, _06750_);
  nor (_07598_, _07597_, _07596_);
  and (_07599_, _07598_, _07595_);
  and (_07600_, _07578_, _07153_);
  nor (_07601_, _07600_, _07152_);
  and (_07602_, _07601_, _07599_);
  and (_07603_, _07152_, _06751_);
  nor (_07604_, _07603_, _07602_);
  and (_07605_, _06608_, _07159_);
  nor (_07606_, _07605_, _07604_);
  and (_07607_, _07606_, _07523_);
  nor (_07608_, _07607_, _07522_);
  and (_07609_, _07165_, _06608_);
  or (_07610_, _07609_, _07608_);
  nor (_07611_, _07515_, _05947_);
  nor (_07612_, _07611_, _06493_);
  not (_07613_, _07612_);
  nor (_07614_, _07613_, _07610_);
  and (_07615_, _07578_, _07174_);
  nor (_07616_, _07615_, _06243_);
  and (_07617_, _07616_, _07614_);
  nor (_07618_, _07617_, _07521_);
  nor (_07619_, _07618_, _05970_);
  and (_07620_, _07515_, _05970_);
  nor (_07621_, _07620_, _07619_);
  or (_07622_, _07621_, _07520_);
  nor (_07623_, _07622_, _07519_);
  and (_07624_, _07578_, _07200_);
  nor (_07625_, _07624_, _07199_);
  and (_07626_, _07625_, _07623_);
  nor (_07627_, _07626_, _07518_);
  nor (_07628_, _07627_, _05895_);
  and (_07629_, _07515_, _05895_);
  nor (_07630_, _07629_, _07628_);
  nor (_07631_, _07222_, _06751_);
  nor (_07632_, _07631_, _07209_);
  not (_07633_, _07632_);
  nor (_07634_, _07633_, _07630_);
  nor (_07635_, _07516_, _05919_);
  nor (_07636_, _07635_, _07634_);
  and (_07637_, _07395_, _06750_);
  or (_07638_, _07637_, _07228_);
  nor (_07639_, _07638_, _07636_);
  nor (_07640_, _07639_, _07517_);
  and (_07641_, _05911_, _06347_);
  nor (_07642_, _07641_, _07640_);
  and (_07643_, _07578_, _07243_);
  nor (_07644_, _07643_, _07242_);
  and (_07645_, _07644_, _07642_);
  and (_07646_, _07242_, _06751_);
  nor (_07647_, _07646_, _07645_);
  nor (_07648_, _07515_, _07250_);
  nor (_07649_, _07648_, _07249_);
  not (_07650_, _07649_);
  nor (_07651_, _07650_, _07647_);
  nor (_07652_, _07651_, _07511_);
  and (_07653_, _06347_, _05906_);
  nor (_07654_, _07653_, _07652_);
  and (_07655_, _07578_, _07259_);
  nor (_07656_, _07655_, _06190_);
  and (_07657_, _07656_, _07654_);
  and (_07658_, _06190_, _06751_);
  nor (_07659_, _07658_, _07657_);
  not (_07660_, _07659_);
  not (_07661_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_07662_, _06982_, _07661_);
  not (_07663_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_07664_, _07067_, _07663_);
  and (_07665_, _07664_, _07065_);
  nand (_07666_, _07665_, _07662_);
  not (_07667_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_07668_, _07067_, _07667_);
  not (_07669_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_07670_, _06982_, _07669_);
  and (_07671_, _07670_, _07073_);
  nand (_07672_, _07671_, _07668_);
  nand (_07673_, _07672_, _07666_);
  nand (_07674_, _07673_, _06763_);
  not (_07675_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_07676_, _07067_, _07675_);
  not (_07677_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_07678_, _06982_, _07677_);
  and (_07679_, _07678_, _07073_);
  nand (_07680_, _07679_, _07676_);
  not (_07681_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_07682_, _06982_, _07681_);
  not (_07683_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_07684_, _07067_, _07683_);
  and (_07685_, _07684_, _07065_);
  nand (_07686_, _07685_, _07682_);
  nand (_07687_, _07686_, _07680_);
  nand (_07688_, _07687_, _07080_);
  nand (_07689_, _07688_, _07674_);
  nand (_07690_, _07689_, _06577_);
  nand (_07691_, _06982_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_07692_, _07067_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_07693_, _07692_, _07073_);
  nand (_07694_, _07693_, _07691_);
  nand (_07695_, _07067_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_07696_, _06982_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_07697_, _07696_, _07065_);
  nand (_07698_, _07697_, _07695_);
  nand (_07699_, _07698_, _07694_);
  nand (_07700_, _07699_, _06763_);
  nand (_07701_, _06982_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_07702_, _07067_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_07703_, _07702_, _07073_);
  nand (_07704_, _07703_, _07701_);
  nand (_07705_, _07067_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_07706_, _06982_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_07707_, _07706_, _07065_);
  nand (_07708_, _07707_, _07705_);
  nand (_07709_, _07708_, _07704_);
  nand (_07710_, _07709_, _07080_);
  nand (_07711_, _07710_, _07700_);
  nand (_07712_, _07711_, _07097_);
  nand (_07713_, _07712_, _07690_);
  and (_07714_, _07713_, _07243_);
  and (_07715_, _06327_, _06241_);
  and (_07716_, _07713_, _07174_);
  nor (_07717_, _07513_, \oc8051_golden_model_1.SP [3]);
  and (_07718_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_07719_, _07718_, \oc8051_golden_model_1.SP [3]);
  and (_07720_, _07719_, \oc8051_golden_model_1.SP [0]);
  nor (_07721_, _07720_, _07717_);
  not (_07722_, _07721_);
  nor (_07723_, _07722_, _05947_);
  and (_07724_, _06253_, _06328_);
  and (_07725_, _07713_, _07134_);
  and (_07726_, _07721_, _06705_);
  and (_07727_, _07713_, _06258_);
  not (_07728_, \oc8051_golden_model_1.PSW [3]);
  and (_07729_, _05960_, _07728_);
  nor (_07730_, _07729_, _07125_);
  not (_07731_, _07730_);
  nor (_07732_, _07731_, _07727_);
  and (_07733_, _07125_, _06328_);
  nor (_07734_, _07733_, _07732_);
  nor (_07735_, _07734_, _06705_);
  or (_07736_, _07735_, _07134_);
  nor (_07737_, _07736_, _07726_);
  or (_07738_, _07737_, _06253_);
  nor (_07739_, _07738_, _07725_);
  nor (_07740_, _07739_, _07724_);
  nor (_07741_, _07740_, _07139_);
  not (_07742_, _06326_);
  and (_07743_, _07742_, _07139_);
  or (_07744_, _07743_, _07474_);
  nor (_07745_, _07744_, _07741_);
  nor (_07746_, _07721_, _05950_);
  nor (_07747_, _07746_, _07143_);
  not (_07748_, _07747_);
  nor (_07749_, _07748_, _07745_);
  and (_07750_, _07143_, _06328_);
  nor (_07751_, _07750_, _07153_);
  not (_07752_, _07751_);
  nor (_07753_, _07752_, _07749_);
  and (_07754_, _07713_, _07153_);
  nor (_07755_, _07754_, _07152_);
  not (_07756_, _07755_);
  nor (_07757_, _07756_, _07753_);
  and (_07758_, _07152_, _06328_);
  or (_07759_, _07758_, _07159_);
  nor (_07760_, _07759_, _07757_);
  and (_07761_, _06326_, _07159_);
  nor (_07762_, _07761_, _07760_);
  and (_07763_, _07762_, _07523_);
  and (_07764_, _07721_, _06247_);
  nor (_07765_, _07764_, _07763_);
  nor (_07766_, _07765_, _07165_);
  nor (_07767_, _07270_, _06330_);
  or (_07768_, _07767_, _07766_);
  and (_07769_, _07768_, _05947_);
  or (_07770_, _07769_, _07174_);
  nor (_07771_, _07770_, _07723_);
  or (_07772_, _07771_, _06243_);
  nor (_07773_, _07772_, _07716_);
  nor (_07774_, _07773_, _07715_);
  nor (_07775_, _07774_, _05970_);
  and (_07776_, _07721_, _05970_);
  not (_07777_, _07776_);
  and (_07778_, _07777_, _07191_);
  not (_07779_, _07778_);
  nor (_07780_, _07779_, _07775_);
  nor (_07781_, _07191_, _06328_);
  nor (_07782_, _07781_, _07780_);
  nor (_07783_, _07782_, _07200_);
  and (_07784_, _07713_, _07200_);
  nor (_07785_, _07784_, _07199_);
  not (_07786_, _07785_);
  nor (_07787_, _07786_, _07783_);
  nor (_07788_, _07198_, _06765_);
  nor (_07789_, _07788_, _07787_);
  nor (_07790_, _07789_, _05895_);
  and (_07791_, _07721_, _05895_);
  not (_07792_, _07791_);
  and (_07793_, _07792_, _07222_);
  not (_07794_, _07793_);
  nor (_07795_, _07794_, _07790_);
  nor (_07796_, _07222_, _06328_);
  nor (_07797_, _07796_, _07209_);
  not (_07798_, _07797_);
  nor (_07799_, _07798_, _07795_);
  nor (_07800_, _07722_, _05919_);
  or (_07801_, _07800_, _07395_);
  nor (_07802_, _07801_, _07799_);
  and (_07803_, _07395_, _06292_);
  or (_07804_, _07803_, _07228_);
  nor (_07805_, _07804_, _07802_);
  nor (_07806_, _07722_, _05916_);
  nor (_07807_, _07806_, _07243_);
  not (_07808_, _07807_);
  nor (_07809_, _07808_, _07805_);
  or (_07810_, _07809_, _07242_);
  nor (_07811_, _07810_, _07714_);
  not (_07812_, _07250_);
  and (_07813_, _07242_, _06328_);
  nor (_07814_, _07813_, _07812_);
  not (_07815_, _07814_);
  nor (_07816_, _07815_, _07811_);
  nor (_07817_, _07721_, _07250_);
  nor (_07818_, _07817_, _07249_);
  not (_07819_, _07818_);
  nor (_07820_, _07819_, _07816_);
  and (_07821_, _07249_, _07742_);
  nor (_07822_, _07821_, _07259_);
  not (_07823_, _07822_);
  nor (_07824_, _07823_, _07820_);
  and (_07825_, _07713_, _07259_);
  nor (_07826_, _07825_, _06190_);
  not (_07827_, _07826_);
  nor (_07828_, _07827_, _07824_);
  and (_07829_, _06190_, _06328_);
  nor (_07830_, _07829_, _07828_);
  nor (_07831_, _07830_, _07508_);
  and (_07832_, _07831_, _07660_);
  and (_07833_, _07832_, _07510_);
  or (_07834_, _07833_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_07835_, _07718_, _06235_);
  or (_07836_, _07515_, _06236_);
  and (_07837_, _07836_, _07835_);
  and (_07838_, _07719_, _06235_);
  and (_07839_, _07835_, _07722_);
  nor (_07840_, _07839_, _07838_);
  and (_07841_, _07272_, _05920_);
  and (_07842_, _07841_, _07250_);
  and (_07843_, _07842_, _07476_);
  nor (_07844_, _07843_, _07420_);
  and (_07845_, _07844_, _07840_);
  and (_07846_, _07845_, _07837_);
  and (_07847_, _07846_, _06234_);
  not (_07848_, _07847_);
  and (_07849_, _07848_, _07834_);
  not (_07850_, _07833_);
  and (_07851_, _06155_, _06799_);
  and (_07852_, _06750_, _06328_);
  and (_07853_, _07852_, _07851_);
  and (_07854_, _06326_, _06187_);
  and (_07855_, _06244_, _06608_);
  and (_07856_, _07855_, _07854_);
  and (_07857_, _07856_, _07853_);
  and (_07858_, _07857_, \oc8051_golden_model_1.SBUF [7]);
  not (_07859_, _07858_);
  and (_07860_, _06155_, _06802_);
  and (_07861_, _07860_, _07852_);
  not (_07862_, _06608_);
  and (_07863_, _06230_, _07862_);
  and (_07864_, _07863_, _07854_);
  and (_07865_, _07864_, _07861_);
  and (_07866_, _07865_, \oc8051_golden_model_1.IE [7]);
  and (_07867_, _06750_, _06292_);
  and (_07868_, _07867_, _07860_);
  nor (_07869_, _06230_, _06608_);
  and (_07870_, _07869_, _07854_);
  and (_07871_, _07870_, _07868_);
  and (_07872_, _07871_, \oc8051_golden_model_1.P3 [7]);
  nor (_07873_, _07872_, _07866_);
  and (_07874_, _07873_, _07859_);
  and (_07875_, _06230_, _06608_);
  and (_07876_, _07875_, _07854_);
  nor (_07877_, _06750_, _06292_);
  and (_07878_, _07877_, _07851_);
  and (_07879_, _07878_, _07876_);
  and (_07880_, _07879_, \oc8051_golden_model_1.TH1 [7]);
  and (_07881_, _07864_, _07868_);
  and (_07882_, _07881_, \oc8051_golden_model_1.P2 [7]);
  nor (_07883_, _07882_, _07880_);
  and (_07884_, _07883_, _07874_);
  and (_07885_, _07876_, _07853_);
  and (_07886_, _07885_, \oc8051_golden_model_1.TMOD [7]);
  not (_07887_, _07886_);
  and (_07888_, _07877_, _07860_);
  and (_07889_, _07888_, _07876_);
  and (_07890_, _07889_, \oc8051_golden_model_1.TH0 [7]);
  nor (_07891_, _06155_, _06799_);
  and (_07892_, _07891_, _07852_);
  and (_07893_, _07892_, _07876_);
  and (_07894_, _07893_, \oc8051_golden_model_1.TL0 [7]);
  nor (_07895_, _07894_, _07890_);
  and (_07896_, _07895_, _07887_);
  and (_07897_, _07876_, _07861_);
  and (_07898_, _07897_, \oc8051_golden_model_1.TCON [7]);
  and (_07899_, _07876_, _07868_);
  and (_07900_, _07899_, \oc8051_golden_model_1.P0 [7]);
  nor (_07901_, _07900_, _07898_);
  and (_07902_, _07901_, _07896_);
  and (_07903_, _07902_, _07884_);
  not (_07904_, _06187_);
  nor (_07905_, _06326_, _07904_);
  and (_07906_, _07905_, _07855_);
  and (_07907_, _07906_, _07868_);
  and (_07908_, _07907_, \oc8051_golden_model_1.PSW [7]);
  not (_07909_, _07908_);
  and (_07910_, _07905_, _07869_);
  and (_07911_, _07910_, _07868_);
  and (_07912_, _07911_, \oc8051_golden_model_1.B [7]);
  and (_07913_, _07863_, _07905_);
  and (_07914_, _07913_, _07868_);
  and (_07915_, _07914_, \oc8051_golden_model_1.ACC [7]);
  nor (_07916_, _07915_, _07912_);
  and (_07917_, _07916_, _07909_);
  and (_07918_, _07870_, _07861_);
  and (_07919_, _07918_, \oc8051_golden_model_1.IP [7]);
  and (_07920_, _07876_, _06292_);
  nor (_07921_, _06155_, _06802_);
  and (_07922_, _07921_, _06751_);
  and (_07923_, _07922_, _07920_);
  and (_07924_, _07923_, \oc8051_golden_model_1.PCON [7]);
  nor (_07925_, _07924_, _07919_);
  and (_07926_, _07925_, _07917_);
  and (_07927_, _07867_, _07851_);
  and (_07928_, _07927_, _07876_);
  and (_07929_, _07928_, \oc8051_golden_model_1.SP [7]);
  not (_07930_, _07929_);
  and (_07931_, _07891_, _06750_);
  and (_07932_, _07931_, _07920_);
  and (_07933_, _07932_, \oc8051_golden_model_1.DPL [7]);
  and (_07934_, _07921_, _07867_);
  and (_07935_, _07934_, _07876_);
  and (_07936_, _07935_, \oc8051_golden_model_1.DPH [7]);
  nor (_07937_, _07936_, _07933_);
  and (_07938_, _07937_, _07930_);
  and (_07939_, _07876_, _07852_);
  and (_07940_, _07921_, _07939_);
  and (_07941_, _07940_, \oc8051_golden_model_1.TL1 [7]);
  not (_07942_, _07941_);
  and (_07943_, _07861_, _07856_);
  and (_07944_, _07943_, \oc8051_golden_model_1.SCON [7]);
  and (_07945_, _07868_, _07856_);
  and (_07946_, _07945_, \oc8051_golden_model_1.P1 [7]);
  nor (_07947_, _07946_, _07944_);
  and (_07948_, _07947_, _07942_);
  and (_07949_, _07948_, _07938_);
  and (_07950_, _07949_, _07926_);
  and (_07951_, _07950_, _07903_);
  not (_07952_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_07953_, _06982_, _07952_);
  not (_07954_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_07955_, _07067_, _07954_);
  and (_07956_, _07955_, _07065_);
  nand (_07957_, _07956_, _07953_);
  not (_07958_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_07959_, _07067_, _07958_);
  not (_07960_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_07961_, _06982_, _07960_);
  and (_07962_, _07961_, _07073_);
  nand (_07963_, _07962_, _07959_);
  nand (_07964_, _07963_, _07957_);
  nand (_07965_, _07964_, _06763_);
  not (_07966_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_07967_, _07067_, _07966_);
  not (_07968_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_07969_, _06982_, _07968_);
  and (_07970_, _07969_, _07073_);
  nand (_07971_, _07970_, _07967_);
  not (_07972_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_07973_, _06982_, _07972_);
  not (_07974_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_07975_, _07067_, _07974_);
  and (_07976_, _07975_, _07065_);
  nand (_07977_, _07976_, _07973_);
  nand (_07978_, _07977_, _07971_);
  nand (_07979_, _07978_, _07080_);
  nand (_07980_, _07979_, _07965_);
  nand (_07981_, _07980_, _06577_);
  nand (_07982_, _06982_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_07983_, _07067_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_07984_, _07983_, _07073_);
  nand (_07985_, _07984_, _07982_);
  nand (_07986_, _07067_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_07987_, _06982_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_07988_, _07987_, _07065_);
  nand (_07989_, _07988_, _07986_);
  nand (_07990_, _07989_, _07985_);
  nand (_07991_, _07990_, _06763_);
  nand (_07992_, _06982_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_07993_, _07067_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_07994_, _07993_, _07073_);
  nand (_07995_, _07994_, _07992_);
  nand (_07996_, _07067_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_07997_, _06982_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_07998_, _07997_, _07065_);
  nand (_07999_, _07998_, _07996_);
  nand (_08000_, _07999_, _07995_);
  nand (_08001_, _08000_, _07080_);
  nand (_08002_, _08001_, _07991_);
  nand (_08003_, _08002_, _07097_);
  nand (_08004_, _08003_, _07981_);
  or (_08005_, _08004_, _06187_);
  and (_08006_, _08005_, _07951_);
  not (_08007_, _08006_);
  and (_08008_, _07857_, \oc8051_golden_model_1.SBUF [6]);
  not (_08009_, _08008_);
  and (_08010_, _07865_, \oc8051_golden_model_1.IE [6]);
  and (_08011_, _07871_, \oc8051_golden_model_1.P3 [6]);
  nor (_08012_, _08011_, _08010_);
  and (_08013_, _08012_, _08009_);
  and (_08014_, _07881_, \oc8051_golden_model_1.P2 [6]);
  and (_08015_, _07940_, \oc8051_golden_model_1.TL1 [6]);
  nor (_08016_, _08015_, _08014_);
  and (_08017_, _08016_, _08013_);
  and (_08018_, _07897_, \oc8051_golden_model_1.TCON [6]);
  not (_08019_, _08018_);
  and (_08020_, _07889_, \oc8051_golden_model_1.TH0 [6]);
  and (_08021_, _07893_, \oc8051_golden_model_1.TL0 [6]);
  nor (_08022_, _08021_, _08020_);
  and (_08023_, _08022_, _08019_);
  and (_08024_, _07885_, \oc8051_golden_model_1.TMOD [6]);
  and (_08025_, _07928_, \oc8051_golden_model_1.SP [6]);
  nor (_08026_, _08025_, _08024_);
  and (_08027_, _08026_, _08023_);
  and (_08028_, _08027_, _08017_);
  and (_08029_, _07918_, \oc8051_golden_model_1.IP [6]);
  not (_08030_, _08029_);
  and (_08031_, _07911_, \oc8051_golden_model_1.B [6]);
  and (_08032_, _07914_, \oc8051_golden_model_1.ACC [6]);
  nor (_08033_, _08032_, _08031_);
  and (_08034_, _08033_, _08030_);
  and (_08035_, _07907_, \oc8051_golden_model_1.PSW [6]);
  and (_08036_, _07923_, \oc8051_golden_model_1.PCON [6]);
  nor (_08037_, _08036_, _08035_);
  and (_08038_, _08037_, _08034_);
  and (_08039_, _07899_, \oc8051_golden_model_1.P0 [6]);
  not (_08040_, _08039_);
  and (_08041_, _07932_, \oc8051_golden_model_1.DPL [6]);
  and (_08042_, _07935_, \oc8051_golden_model_1.DPH [6]);
  nor (_08043_, _08042_, _08041_);
  and (_08044_, _08043_, _08040_);
  and (_08045_, _07879_, \oc8051_golden_model_1.TH1 [6]);
  not (_08046_, _08045_);
  and (_08047_, _07945_, \oc8051_golden_model_1.P1 [6]);
  and (_08048_, _07943_, \oc8051_golden_model_1.SCON [6]);
  nor (_08049_, _08048_, _08047_);
  and (_08050_, _08049_, _08046_);
  and (_08051_, _08050_, _08044_);
  and (_08052_, _08051_, _08038_);
  and (_08053_, _08052_, _08028_);
  not (_08054_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_08055_, _06982_, _08054_);
  not (_08056_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_08057_, _07067_, _08056_);
  and (_08058_, _08057_, _07065_);
  nand (_08059_, _08058_, _08055_);
  not (_08060_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_08061_, _07067_, _08060_);
  not (_08062_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_08063_, _06982_, _08062_);
  and (_08064_, _08063_, _07073_);
  nand (_08065_, _08064_, _08061_);
  nand (_08066_, _08065_, _08059_);
  nand (_08067_, _08066_, _06763_);
  not (_08068_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_08069_, _07067_, _08068_);
  not (_08070_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_08071_, _06982_, _08070_);
  and (_08072_, _08071_, _07073_);
  nand (_08073_, _08072_, _08069_);
  not (_08074_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_08075_, _06982_, _08074_);
  not (_08076_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_08077_, _07067_, _08076_);
  and (_08078_, _08077_, _07065_);
  nand (_08079_, _08078_, _08075_);
  nand (_08080_, _08079_, _08073_);
  nand (_08081_, _08080_, _07080_);
  nand (_08082_, _08081_, _08067_);
  nand (_08083_, _08082_, _06577_);
  nand (_08084_, _06982_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_08085_, _07067_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_08086_, _08085_, _07073_);
  nand (_08087_, _08086_, _08084_);
  nand (_08088_, _07067_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_08089_, _06982_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_08090_, _08089_, _07065_);
  nand (_08091_, _08090_, _08088_);
  nand (_08092_, _08091_, _08087_);
  nand (_08093_, _08092_, _06763_);
  nand (_08094_, _06982_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_08095_, _07067_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_08096_, _08095_, _07073_);
  nand (_08097_, _08096_, _08094_);
  nand (_08098_, _07067_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_08099_, _06982_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_08100_, _08099_, _07065_);
  nand (_08101_, _08100_, _08098_);
  nand (_08102_, _08101_, _08097_);
  nand (_08103_, _08102_, _07080_);
  nand (_08104_, _08103_, _08093_);
  nand (_08105_, _08104_, _07097_);
  nand (_08106_, _08105_, _08083_);
  or (_08107_, _08106_, _06187_);
  and (_08108_, _08107_, _08053_);
  not (_08109_, _08108_);
  and (_08110_, _07907_, \oc8051_golden_model_1.PSW [5]);
  and (_08111_, _07911_, \oc8051_golden_model_1.B [5]);
  nor (_08112_, _08111_, _08110_);
  and (_08113_, _07881_, \oc8051_golden_model_1.P2 [5]);
  and (_08114_, _07865_, \oc8051_golden_model_1.IE [5]);
  nor (_08115_, _08114_, _08113_);
  and (_08116_, _08115_, _08112_);
  and (_08117_, _07918_, \oc8051_golden_model_1.IP [5]);
  and (_08118_, _07914_, \oc8051_golden_model_1.ACC [5]);
  nor (_08119_, _08118_, _08117_);
  and (_08120_, _07889_, \oc8051_golden_model_1.TH0 [5]);
  and (_08121_, _07871_, \oc8051_golden_model_1.P3 [5]);
  nor (_08122_, _08121_, _08120_);
  and (_08123_, _08122_, _08119_);
  and (_08124_, _07945_, \oc8051_golden_model_1.P1 [5]);
  and (_08125_, _07943_, \oc8051_golden_model_1.SCON [5]);
  nor (_08126_, _08125_, _08124_);
  and (_08127_, _07879_, \oc8051_golden_model_1.TH1 [5]);
  and (_08128_, _07857_, \oc8051_golden_model_1.SBUF [5]);
  nor (_08129_, _08128_, _08127_);
  and (_08130_, _08129_, _08126_);
  and (_08131_, _08130_, _08123_);
  and (_08132_, _08131_, _08116_);
  and (_08133_, _07932_, \oc8051_golden_model_1.DPL [5]);
  and (_08134_, _07851_, _06750_);
  and (_08135_, _07920_, _08134_);
  and (_08136_, _08135_, \oc8051_golden_model_1.SP [5]);
  nor (_08137_, _08136_, _08133_);
  and (_08138_, _07899_, \oc8051_golden_model_1.P0 [5]);
  and (_08139_, _07939_, _07891_);
  and (_08140_, _08139_, \oc8051_golden_model_1.TL0 [5]);
  nor (_08141_, _08140_, _08138_);
  and (_08142_, _08141_, _08137_);
  and (_08143_, _07923_, \oc8051_golden_model_1.PCON [5]);
  not (_08144_, _08143_);
  and (_08145_, _07897_, \oc8051_golden_model_1.TCON [5]);
  and (_08146_, _07885_, \oc8051_golden_model_1.TMOD [5]);
  nor (_08147_, _08146_, _08145_);
  and (_08148_, _08147_, _08144_);
  and (_08149_, _07940_, \oc8051_golden_model_1.TL1 [5]);
  and (_08150_, _07921_, _06750_);
  and (_08151_, _08150_, _07920_);
  and (_08152_, _08151_, \oc8051_golden_model_1.DPH [5]);
  nor (_08153_, _08152_, _08149_);
  and (_08154_, _08153_, _08148_);
  and (_08155_, _08154_, _08142_);
  and (_08156_, _08155_, _08132_);
  not (_08157_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_08158_, _06982_, _08157_);
  not (_08159_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_08160_, _07067_, _08159_);
  and (_08161_, _08160_, _07065_);
  nand (_08162_, _08161_, _08158_);
  not (_08163_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_08164_, _07067_, _08163_);
  not (_08165_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_08166_, _06982_, _08165_);
  and (_08167_, _08166_, _07073_);
  nand (_08168_, _08167_, _08164_);
  nand (_08169_, _08168_, _08162_);
  nand (_08170_, _08169_, _06763_);
  not (_08171_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_08172_, _07067_, _08171_);
  not (_08173_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_08174_, _06982_, _08173_);
  and (_08175_, _08174_, _07073_);
  nand (_08176_, _08175_, _08172_);
  not (_08177_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_08178_, _06982_, _08177_);
  not (_08179_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_08180_, _07067_, _08179_);
  and (_08181_, _08180_, _07065_);
  nand (_08182_, _08181_, _08178_);
  nand (_08183_, _08182_, _08176_);
  nand (_08184_, _08183_, _07080_);
  nand (_08185_, _08184_, _08170_);
  nand (_08186_, _08185_, _06577_);
  nand (_08187_, _06982_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_08188_, _07067_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_08189_, _08188_, _07073_);
  nand (_08190_, _08189_, _08187_);
  nand (_08191_, _07067_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_08192_, _06982_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_08193_, _08192_, _07065_);
  nand (_08194_, _08193_, _08191_);
  nand (_08195_, _08194_, _08190_);
  nand (_08196_, _08195_, _06763_);
  nand (_08197_, _06982_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_08198_, _07067_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_08199_, _08198_, _07073_);
  nand (_08200_, _08199_, _08197_);
  nand (_08201_, _07067_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_08202_, _06982_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_08203_, _08202_, _07065_);
  nand (_08204_, _08203_, _08201_);
  nand (_08205_, _08204_, _08200_);
  nand (_08206_, _08205_, _07080_);
  nand (_08207_, _08206_, _08196_);
  nand (_08208_, _08207_, _07097_);
  nand (_08209_, _08208_, _08186_);
  or (_08210_, _08209_, _06187_);
  and (_08211_, _08210_, _08156_);
  not (_08212_, _08211_);
  and (_08213_, _07943_, \oc8051_golden_model_1.SCON [3]);
  and (_08214_, _07881_, \oc8051_golden_model_1.P2 [3]);
  nor (_08215_, _08214_, _08213_);
  and (_08216_, _07865_, \oc8051_golden_model_1.IE [3]);
  and (_08217_, _07911_, \oc8051_golden_model_1.B [3]);
  nor (_08218_, _08217_, _08216_);
  and (_08219_, _08218_, _08215_);
  and (_08220_, _07889_, \oc8051_golden_model_1.TH0 [3]);
  and (_08221_, _07907_, \oc8051_golden_model_1.PSW [3]);
  nor (_08222_, _08221_, _08220_);
  and (_08223_, _07871_, \oc8051_golden_model_1.P3 [3]);
  and (_08224_, _07914_, \oc8051_golden_model_1.ACC [3]);
  nor (_08225_, _08224_, _08223_);
  and (_08226_, _08225_, _08222_);
  and (_08227_, _07879_, \oc8051_golden_model_1.TH1 [3]);
  and (_08228_, _07945_, \oc8051_golden_model_1.P1 [3]);
  nor (_08229_, _08228_, _08227_);
  and (_08230_, _07857_, \oc8051_golden_model_1.SBUF [3]);
  and (_08231_, _07918_, \oc8051_golden_model_1.IP [3]);
  nor (_08232_, _08231_, _08230_);
  and (_08233_, _08232_, _08229_);
  and (_08234_, _08233_, _08226_);
  and (_08235_, _08234_, _08219_);
  and (_08236_, _07932_, \oc8051_golden_model_1.DPL [3]);
  and (_08237_, _07935_, \oc8051_golden_model_1.DPH [3]);
  nor (_08238_, _08237_, _08236_);
  and (_08239_, _08135_, \oc8051_golden_model_1.SP [3]);
  and (_08240_, _08139_, \oc8051_golden_model_1.TL0 [3]);
  nor (_08241_, _08240_, _08239_);
  and (_08242_, _08241_, _08238_);
  and (_08243_, _07923_, \oc8051_golden_model_1.PCON [3]);
  not (_08244_, _08243_);
  and (_08245_, _07897_, \oc8051_golden_model_1.TCON [3]);
  and (_08246_, _07885_, \oc8051_golden_model_1.TMOD [3]);
  nor (_08247_, _08246_, _08245_);
  and (_08248_, _08247_, _08244_);
  and (_08249_, _07899_, \oc8051_golden_model_1.P0 [3]);
  and (_08250_, _07940_, \oc8051_golden_model_1.TL1 [3]);
  nor (_08251_, _08250_, _08249_);
  and (_08252_, _08251_, _08248_);
  and (_08253_, _08252_, _08242_);
  and (_08254_, _08253_, _08235_);
  or (_08255_, _07713_, _06187_);
  and (_08256_, _08255_, _08254_);
  not (_08257_, _08256_);
  and (_08258_, _07907_, \oc8051_golden_model_1.PSW [1]);
  and (_08259_, _07914_, \oc8051_golden_model_1.ACC [1]);
  nor (_08260_, _08259_, _08258_);
  and (_08261_, _07881_, \oc8051_golden_model_1.P2 [1]);
  and (_08262_, _07871_, \oc8051_golden_model_1.P3 [1]);
  nor (_08263_, _08262_, _08261_);
  and (_08264_, _08263_, _08260_);
  and (_08265_, _07857_, \oc8051_golden_model_1.SBUF [1]);
  and (_08266_, _07918_, \oc8051_golden_model_1.IP [1]);
  nor (_08267_, _08266_, _08265_);
  and (_08268_, _07885_, \oc8051_golden_model_1.TMOD [1]);
  and (_08269_, _07889_, \oc8051_golden_model_1.TH0 [1]);
  nor (_08270_, _08269_, _08268_);
  and (_08271_, _08270_, _08267_);
  and (_08272_, _07943_, \oc8051_golden_model_1.SCON [1]);
  and (_08273_, _07865_, \oc8051_golden_model_1.IE [1]);
  nor (_08274_, _08273_, _08272_);
  and (_08275_, _07897_, \oc8051_golden_model_1.TCON [1]);
  and (_08276_, _07911_, \oc8051_golden_model_1.B [1]);
  nor (_08277_, _08276_, _08275_);
  and (_08278_, _08277_, _08274_);
  and (_08279_, _08278_, _08271_);
  and (_08280_, _08279_, _08264_);
  and (_08281_, _07932_, \oc8051_golden_model_1.DPL [1]);
  and (_08282_, _08151_, \oc8051_golden_model_1.DPH [1]);
  nor (_08283_, _08282_, _08281_);
  and (_08284_, _08135_, \oc8051_golden_model_1.SP [1]);
  and (_08285_, _08139_, \oc8051_golden_model_1.TL0 [1]);
  nor (_08286_, _08285_, _08284_);
  and (_08287_, _08286_, _08283_);
  and (_08288_, _07940_, \oc8051_golden_model_1.TL1 [1]);
  not (_08289_, _08288_);
  and (_08290_, _07879_, \oc8051_golden_model_1.TH1 [1]);
  and (_08291_, _07945_, \oc8051_golden_model_1.P1 [1]);
  nor (_08292_, _08291_, _08290_);
  and (_08293_, _08292_, _08289_);
  and (_08294_, _07899_, \oc8051_golden_model_1.P0 [1]);
  and (_08295_, _07923_, \oc8051_golden_model_1.PCON [1]);
  nor (_08296_, _08295_, _08294_);
  and (_08297_, _08296_, _08293_);
  and (_08298_, _08297_, _08287_);
  and (_08299_, _08298_, _08280_);
  or (_08300_, _07120_, _06187_);
  and (_08301_, _08300_, _08299_);
  not (_08302_, _08301_);
  and (_08303_, _07881_, \oc8051_golden_model_1.P2 [0]);
  not (_08304_, _08303_);
  and (_08305_, _07857_, \oc8051_golden_model_1.SBUF [0]);
  not (_08306_, _08305_);
  and (_08307_, _07865_, \oc8051_golden_model_1.IE [0]);
  and (_08308_, _07871_, \oc8051_golden_model_1.P3 [0]);
  nor (_08309_, _08308_, _08307_);
  and (_08310_, _08309_, _08306_);
  and (_08311_, _08310_, _08304_);
  and (_08312_, _07932_, \oc8051_golden_model_1.DPL [0]);
  and (_08313_, _07935_, \oc8051_golden_model_1.DPH [0]);
  nor (_08314_, _08313_, _08312_);
  and (_08315_, _07928_, \oc8051_golden_model_1.SP [0]);
  not (_08316_, _08315_);
  and (_08317_, _08316_, _08314_);
  and (_08318_, _07945_, \oc8051_golden_model_1.P1 [0]);
  and (_08319_, _07943_, \oc8051_golden_model_1.SCON [0]);
  nor (_08320_, _08319_, _08318_);
  and (_08321_, _07879_, \oc8051_golden_model_1.TH1 [0]);
  and (_08322_, _07940_, \oc8051_golden_model_1.TL1 [0]);
  nor (_08323_, _08322_, _08321_);
  and (_08324_, _08323_, _08320_);
  and (_08325_, _08324_, _08317_);
  and (_08326_, _08325_, _08311_);
  and (_08327_, _07907_, \oc8051_golden_model_1.PSW [0]);
  not (_08328_, _08327_);
  and (_08329_, _07914_, \oc8051_golden_model_1.ACC [0]);
  and (_08330_, _07911_, \oc8051_golden_model_1.B [0]);
  nor (_08331_, _08330_, _08329_);
  and (_08332_, _08331_, _08328_);
  and (_08333_, _07918_, \oc8051_golden_model_1.IP [0]);
  and (_08334_, _07923_, \oc8051_golden_model_1.PCON [0]);
  nor (_08335_, _08334_, _08333_);
  and (_08336_, _08335_, _08332_);
  and (_08337_, _07885_, \oc8051_golden_model_1.TMOD [0]);
  not (_08338_, _08337_);
  and (_08339_, _07889_, \oc8051_golden_model_1.TH0 [0]);
  and (_08340_, _07893_, \oc8051_golden_model_1.TL0 [0]);
  nor (_08341_, _08340_, _08339_);
  and (_08342_, _08341_, _08338_);
  and (_08343_, _07899_, \oc8051_golden_model_1.P0 [0]);
  and (_08344_, _07897_, \oc8051_golden_model_1.TCON [0]);
  nor (_08345_, _08344_, _08343_);
  and (_08346_, _08345_, _08342_);
  and (_08347_, _08346_, _08336_);
  and (_08348_, _08347_, _08326_);
  not (_08349_, _08348_);
  and (_08350_, _07325_, _07904_);
  or (_08351_, _08350_, _08349_);
  and (_08352_, _08351_, _08302_);
  and (_08353_, _07907_, \oc8051_golden_model_1.PSW [2]);
  and (_08354_, _07914_, \oc8051_golden_model_1.ACC [2]);
  nor (_08355_, _08354_, _08353_);
  and (_08356_, _07885_, \oc8051_golden_model_1.TMOD [2]);
  and (_08357_, _07918_, \oc8051_golden_model_1.IP [2]);
  nor (_08358_, _08357_, _08356_);
  and (_08359_, _08358_, _08355_);
  and (_08360_, _07945_, \oc8051_golden_model_1.P1 [2]);
  and (_08361_, _07871_, \oc8051_golden_model_1.P3 [2]);
  nor (_08362_, _08361_, _08360_);
  and (_08363_, _07889_, \oc8051_golden_model_1.TH0 [2]);
  and (_08364_, _07911_, \oc8051_golden_model_1.B [2]);
  nor (_08365_, _08364_, _08363_);
  and (_08366_, _08365_, _08362_);
  and (_08367_, _07943_, \oc8051_golden_model_1.SCON [2]);
  and (_08368_, _07881_, \oc8051_golden_model_1.P2 [2]);
  nor (_08369_, _08368_, _08367_);
  and (_08370_, _07879_, \oc8051_golden_model_1.TH1 [2]);
  and (_08371_, _07865_, \oc8051_golden_model_1.IE [2]);
  nor (_08372_, _08371_, _08370_);
  and (_08373_, _08372_, _08369_);
  and (_08374_, _08373_, _08366_);
  and (_08375_, _08374_, _08359_);
  and (_08376_, _07932_, \oc8051_golden_model_1.DPL [2]);
  and (_08377_, _08135_, \oc8051_golden_model_1.SP [2]);
  nor (_08378_, _08377_, _08376_);
  and (_08379_, _07940_, \oc8051_golden_model_1.TL1 [2]);
  and (_08380_, _08139_, \oc8051_golden_model_1.TL0 [2]);
  nor (_08381_, _08380_, _08379_);
  and (_08382_, _08381_, _08378_);
  and (_08383_, _07923_, \oc8051_golden_model_1.PCON [2]);
  not (_08384_, _08383_);
  and (_08385_, _07897_, \oc8051_golden_model_1.TCON [2]);
  and (_08386_, _07857_, \oc8051_golden_model_1.SBUF [2]);
  nor (_08387_, _08386_, _08385_);
  and (_08388_, _08387_, _08384_);
  and (_08389_, _07899_, \oc8051_golden_model_1.P0 [2]);
  and (_08390_, _08151_, \oc8051_golden_model_1.DPH [2]);
  nor (_08391_, _08390_, _08389_);
  and (_08392_, _08391_, _08388_);
  and (_08393_, _08392_, _08382_);
  and (_08394_, _08393_, _08375_);
  or (_08395_, _07578_, _06187_);
  and (_08396_, _08395_, _08394_);
  not (_08397_, _08396_);
  and (_08398_, _08397_, _08352_);
  and (_08399_, _08398_, _08257_);
  and (_08400_, _07865_, \oc8051_golden_model_1.IE [4]);
  and (_08401_, _07907_, \oc8051_golden_model_1.PSW [4]);
  nor (_08402_, _08401_, _08400_);
  and (_08403_, _07945_, \oc8051_golden_model_1.P1 [4]);
  and (_08404_, _07911_, \oc8051_golden_model_1.B [4]);
  nor (_08405_, _08404_, _08403_);
  and (_08406_, _08405_, _08402_);
  and (_08407_, _07897_, \oc8051_golden_model_1.TCON [4]);
  and (_08408_, _07914_, \oc8051_golden_model_1.ACC [4]);
  nor (_08409_, _08408_, _08407_);
  and (_08410_, _07885_, \oc8051_golden_model_1.TMOD [4]);
  and (_08411_, _07871_, \oc8051_golden_model_1.P3 [4]);
  nor (_08412_, _08411_, _08410_);
  and (_08413_, _08412_, _08409_);
  and (_08414_, _07943_, \oc8051_golden_model_1.SCON [4]);
  and (_08415_, _07918_, \oc8051_golden_model_1.IP [4]);
  nor (_08416_, _08415_, _08414_);
  and (_08417_, _07879_, \oc8051_golden_model_1.TH1 [4]);
  and (_08418_, _07881_, \oc8051_golden_model_1.P2 [4]);
  nor (_08419_, _08418_, _08417_);
  and (_08420_, _08419_, _08416_);
  and (_08421_, _08420_, _08413_);
  and (_08422_, _08421_, _08406_);
  and (_08423_, _07932_, \oc8051_golden_model_1.DPL [4]);
  and (_08424_, _07940_, \oc8051_golden_model_1.TL1 [4]);
  nor (_08425_, _08424_, _08423_);
  and (_08426_, _07923_, \oc8051_golden_model_1.PCON [4]);
  and (_08427_, _08139_, \oc8051_golden_model_1.TL0 [4]);
  nor (_08428_, _08427_, _08426_);
  and (_08429_, _08428_, _08425_);
  and (_08430_, _07899_, \oc8051_golden_model_1.P0 [4]);
  and (_08431_, _07928_, \oc8051_golden_model_1.SP [4]);
  nor (_08432_, _08431_, _08430_);
  and (_08433_, _08151_, \oc8051_golden_model_1.DPH [4]);
  not (_08434_, _08433_);
  and (_08435_, _07889_, \oc8051_golden_model_1.TH0 [4]);
  and (_08436_, _07857_, \oc8051_golden_model_1.SBUF [4]);
  nor (_08437_, _08436_, _08435_);
  and (_08438_, _08437_, _08434_);
  and (_08439_, _08438_, _08432_);
  and (_08440_, _08439_, _08429_);
  and (_08441_, _08440_, _08422_);
  not (_08442_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_08443_, _06982_, _08442_);
  not (_08444_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_08445_, _07067_, _08444_);
  and (_08446_, _08445_, _07065_);
  nand (_08447_, _08446_, _08443_);
  not (_08448_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_08449_, _07067_, _08448_);
  not (_08450_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_08451_, _06982_, _08450_);
  and (_08452_, _08451_, _07073_);
  nand (_08453_, _08452_, _08449_);
  nand (_08454_, _08453_, _08447_);
  nand (_08455_, _08454_, _06763_);
  not (_08456_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_08457_, _07067_, _08456_);
  not (_08458_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_08459_, _06982_, _08458_);
  and (_08460_, _08459_, _07073_);
  nand (_08461_, _08460_, _08457_);
  not (_08462_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_08463_, _06982_, _08462_);
  not (_08464_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_08465_, _07067_, _08464_);
  and (_08466_, _08465_, _07065_);
  nand (_08467_, _08466_, _08463_);
  nand (_08468_, _08467_, _08461_);
  nand (_08469_, _08468_, _07080_);
  nand (_08470_, _08469_, _08455_);
  nand (_08471_, _08470_, _06577_);
  nand (_08472_, _06982_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_08473_, _07067_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_08474_, _08473_, _07073_);
  nand (_08475_, _08474_, _08472_);
  nand (_08476_, _07067_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_08477_, _06982_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_08478_, _08477_, _07065_);
  nand (_08479_, _08478_, _08476_);
  nand (_08480_, _08479_, _08475_);
  nand (_08481_, _08480_, _06763_);
  nand (_08482_, _06982_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_08483_, _07067_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_08484_, _08483_, _07073_);
  nand (_08485_, _08484_, _08482_);
  nand (_08486_, _07067_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_08487_, _06982_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_08488_, _08487_, _07065_);
  nand (_08489_, _08488_, _08486_);
  nand (_08490_, _08489_, _08485_);
  nand (_08491_, _08490_, _07080_);
  nand (_08492_, _08491_, _08481_);
  nand (_08493_, _08492_, _07097_);
  nand (_08494_, _08493_, _08471_);
  or (_08495_, _08494_, _06187_);
  and (_08496_, _08495_, _08441_);
  not (_08497_, _08496_);
  and (_08498_, _08497_, _08399_);
  and (_08499_, _08498_, _08212_);
  and (_08500_, _08499_, _08109_);
  nor (_08501_, _08500_, _08007_);
  and (_08502_, _08500_, _08007_);
  nor (_08503_, _08502_, _08501_);
  and (_08504_, _08503_, _06190_);
  not (_08505_, _06378_);
  not (_08506_, \oc8051_golden_model_1.ACC [7]);
  nor (_08507_, _08006_, _08506_);
  and (_08508_, _08006_, _08506_);
  nor (_08509_, _08508_, _08507_);
  and (_08510_, _08509_, _07217_);
  not (_08511_, _07217_);
  not (_08512_, _07189_);
  and (_08513_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_08514_, _08513_, \oc8051_golden_model_1.PC [6]);
  and (_08515_, _08514_, _06073_);
  and (_08516_, _08515_, \oc8051_golden_model_1.PC [7]);
  nor (_08517_, _08515_, \oc8051_golden_model_1.PC [7]);
  nor (_08518_, _08517_, _08516_);
  and (_08519_, _08518_, _05970_);
  not (_08520_, _07139_);
  not (_08521_, _07922_);
  and (_08522_, _07920_, \oc8051_golden_model_1.P0 [7]);
  not (_08523_, _06330_);
  not (_08524_, _06765_);
  or (_08525_, _06609_, _08524_);
  nor (_08526_, _08525_, _06231_);
  and (_08527_, _08526_, _08523_);
  and (_08528_, _08527_, _07876_);
  and (_08529_, _08528_, \oc8051_golden_model_1.TCON [7]);
  and (_08530_, _08526_, _06330_);
  and (_08531_, _08530_, _07856_);
  and (_08532_, _08531_, \oc8051_golden_model_1.P1 [7]);
  and (_08533_, _08527_, _07856_);
  and (_08534_, _08533_, \oc8051_golden_model_1.SCON [7]);
  and (_08535_, _08530_, _07864_);
  and (_08536_, _08535_, \oc8051_golden_model_1.P2 [7]);
  and (_08537_, _08527_, _07864_);
  and (_08538_, _08537_, \oc8051_golden_model_1.IE [7]);
  and (_08539_, _08530_, _07870_);
  and (_08540_, _08539_, \oc8051_golden_model_1.P3 [7]);
  and (_08541_, _08527_, _07870_);
  and (_08542_, _08541_, \oc8051_golden_model_1.IP [7]);
  and (_08543_, _07906_, _08530_);
  and (_08544_, _08543_, \oc8051_golden_model_1.PSW [7]);
  and (_08545_, _08530_, _07913_);
  and (_08546_, _08545_, \oc8051_golden_model_1.ACC [7]);
  and (_08547_, _08530_, _07910_);
  and (_08548_, _08547_, \oc8051_golden_model_1.B [7]);
  or (_08549_, _08548_, _08546_);
  or (_08550_, _08549_, _08544_);
  or (_08551_, _08550_, _08542_);
  or (_08552_, _08551_, _08540_);
  or (_08553_, _08552_, _08538_);
  or (_08554_, _08553_, _08536_);
  or (_08555_, _08554_, _08534_);
  or (_08556_, _08555_, _08532_);
  or (_08557_, _08556_, _08529_);
  nor (_08558_, _08557_, _08522_);
  and (_08559_, _08558_, _08005_);
  nand (_08560_, _08559_, _08521_);
  or (_08561_, _08560_, _08520_);
  not (_08562_, _08004_);
  and (_08563_, _08494_, _08209_);
  and (_08564_, _07578_, _07713_);
  and (_08565_, _07120_, _07380_);
  and (_08566_, _08565_, _08564_);
  and (_08567_, _08566_, _08563_);
  and (_08568_, _08567_, _08106_);
  nor (_08569_, _08568_, _08562_);
  and (_08570_, _08568_, _08562_);
  nor (_08571_, _08570_, _08569_);
  nor (_08572_, _05949_, _05965_);
  not (_08573_, _08572_);
  or (_08574_, _08573_, _08571_);
  nor (_08575_, _06705_, _08506_);
  and (_08576_, _06250_, _06348_);
  and (_08577_, _06250_, _06192_);
  or (_08578_, _08577_, _08576_);
  or (_08579_, _08578_, _08575_);
  and (_08580_, _08518_, _06705_);
  not (_08581_, _06197_);
  and (_08582_, _07584_, _08581_);
  or (_08583_, _08582_, _08580_);
  or (_08584_, _08583_, _08579_);
  and (_08585_, _08584_, _08574_);
  or (_08586_, _08585_, _07134_);
  not (_08587_, _07027_);
  nor (_08588_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_08589_, _08588_, _06670_);
  nor (_08590_, _08589_, _06559_);
  nor (_08591_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_08592_, _08591_, _06559_);
  and (_08593_, _08592_, _06235_);
  nor (_08594_, _08593_, _08590_);
  and (_08595_, _08594_, _08587_);
  and (_08596_, _07174_, _06292_);
  and (_08597_, _07713_, _07369_);
  nor (_08598_, _08597_, _08596_);
  nor (_08599_, _08598_, _08587_);
  nor (_08600_, _08599_, _08595_);
  or (_08601_, _07174_, _07325_);
  and (_08602_, _07174_, _06802_);
  nor (_08603_, _08602_, _08587_);
  nand (_08604_, _08603_, _08601_);
  nor (_08605_, _07027_, \oc8051_golden_model_1.SP [0]);
  not (_08606_, _08605_);
  and (_08607_, _08606_, _08604_);
  nor (_08608_, _07578_, _07174_);
  nor (_08609_, _07369_, _06750_);
  nor (_08610_, _08609_, _08587_);
  not (_08611_, _08610_);
  nor (_08612_, _08611_, _08608_);
  nor (_08613_, _08588_, _06670_);
  nor (_08614_, _08613_, _08589_);
  and (_08615_, _08614_, _08587_);
  nor (_08616_, _08615_, _08612_);
  not (_08617_, _08616_);
  nand (_08618_, _08617_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor (_08619_, _07369_, _06155_);
  nor (_08620_, _07120_, _07174_);
  or (_08621_, _08620_, _08619_);
  nand (_08622_, _08621_, _07027_);
  nor (_08623_, _06248_, _07027_);
  not (_08624_, _08623_);
  and (_08625_, _08624_, _08622_);
  and (_08626_, _08616_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_08627_, _08626_, _08625_);
  and (_08628_, _08627_, _08618_);
  nand (_08629_, _08617_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_08630_, _08616_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_08631_, _08630_, _08625_);
  and (_08632_, _08631_, _08629_);
  or (_08633_, _08632_, _08628_);
  and (_08634_, _08633_, _08607_);
  not (_08635_, _08607_);
  nand (_08636_, _08617_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_08637_, _08616_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor (_08638_, _08637_, _08625_);
  and (_08639_, _08638_, _08636_);
  nand (_08640_, _08617_, \oc8051_golden_model_1.IRAM[9] [7]);
  nand (_08641_, _08616_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_08642_, _08641_, _08625_);
  and (_08643_, _08642_, _08640_);
  or (_08644_, _08643_, _08639_);
  and (_08645_, _08644_, _08635_);
  or (_08646_, _08645_, _08634_);
  nand (_08647_, _08646_, _08600_);
  not (_08648_, _08600_);
  nand (_08649_, _08607_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor (_08650_, _08607_, _07966_);
  nor (_08651_, _08650_, _08625_);
  nand (_08652_, _08651_, _08649_);
  nand (_08653_, _08607_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_08654_, _08607_, _07974_);
  and (_08655_, _08654_, _08625_);
  nand (_08656_, _08655_, _08653_);
  nand (_08657_, _08656_, _08652_);
  nand (_08658_, _08657_, _08616_);
  nand (_08659_, _08607_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor (_08660_, _08607_, _07958_);
  nor (_08661_, _08660_, _08625_);
  nand (_08662_, _08661_, _08659_);
  nand (_08663_, _08607_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_08664_, _08607_, _07954_);
  and (_08665_, _08664_, _08625_);
  nand (_08666_, _08665_, _08663_);
  nand (_08667_, _08666_, _08662_);
  nand (_08668_, _08667_, _08617_);
  nand (_08669_, _08668_, _08658_);
  nand (_08670_, _08669_, _08648_);
  and (_08671_, _08670_, _08647_);
  or (_08672_, _08671_, _07338_);
  and (_08673_, _08672_, _08586_);
  or (_08674_, _08673_, _06253_);
  not (_08675_, _06253_);
  and (_08676_, _08496_, _08211_);
  not (_08677_, _08351_);
  and (_08678_, _08677_, _08301_);
  and (_08679_, _08396_, _08256_);
  and (_08680_, _08679_, _08678_);
  and (_08681_, _08680_, _08676_);
  and (_08682_, _08681_, _08108_);
  nor (_08683_, _08682_, _08007_);
  and (_08684_, _08682_, _08007_);
  nor (_08685_, _08684_, _08683_);
  or (_08686_, _08685_, _08675_);
  and (_08687_, _08686_, _08674_);
  or (_08688_, _08687_, _07139_);
  and (_08689_, _08688_, _08561_);
  or (_08690_, _08689_, _07474_);
  nor (_08691_, _08518_, _05950_);
  nor (_08692_, _08691_, _07143_);
  and (_08693_, _08692_, _08690_);
  and (_08694_, _08562_, _07143_);
  or (_08695_, _08694_, _07159_);
  or (_08696_, _08695_, _08693_);
  not (_08697_, _07159_);
  nor (_08698_, _08559_, _07922_);
  or (_08699_, _08698_, _08697_);
  and (_08700_, _08699_, _08696_);
  or (_08701_, _08700_, _06247_);
  nand (_08702_, _08006_, _06247_);
  and (_08703_, _08702_, _07270_);
  and (_08704_, _08703_, _08701_);
  nor (_08705_, _08559_, _08521_);
  not (_08706_, _08705_);
  and (_08707_, _08706_, _08560_);
  and (_08708_, _08707_, _07165_);
  or (_08709_, _08708_, _08704_);
  and (_08710_, _08709_, _05947_);
  not (_08711_, _08518_);
  or (_08712_, _08711_, _05947_);
  nand (_08713_, _08712_, _06497_);
  or (_08714_, _08713_, _08710_);
  nand (_08715_, _08006_, _06498_);
  and (_08716_, _08715_, _07369_);
  and (_08717_, _08716_, _08714_);
  nand (_08718_, _08671_, _07904_);
  nand (_08719_, _08718_, _07951_);
  and (_08720_, _08719_, _07174_);
  or (_08721_, _08720_, _06243_);
  or (_08722_, _08721_, _08717_);
  not (_08723_, _05970_);
  not (_08724_, _06243_);
  and (_08725_, _07922_, \oc8051_golden_model_1.PSW [7]);
  or (_08726_, _08725_, _08698_);
  or (_08727_, _08726_, _08724_);
  and (_08728_, _08727_, _08723_);
  and (_08729_, _08728_, _08722_);
  or (_08730_, _08729_, _08519_);
  and (_08731_, _08730_, _08512_);
  nor (_08732_, _08004_, _08512_);
  or (_08733_, _08732_, _07184_);
  or (_08734_, _08733_, _08731_);
  not (_08735_, _07186_);
  or (_08736_, _08671_, _07185_);
  and (_08737_, _08736_, _08735_);
  and (_08738_, _08737_, _08734_);
  and (_08739_, _06404_, _00715_);
  and (_08740_, _06421_, _00532_);
  nor (_08741_, _08740_, _08739_);
  and (_08742_, _06451_, _00286_);
  and (_08743_, _06429_, _00091_);
  nor (_08744_, _08743_, _08742_);
  and (_08745_, _08744_, _08741_);
  and (_08746_, _06412_, _00674_);
  and (_08747_, _06434_, _00633_);
  nor (_08748_, _08747_, _08746_);
  and (_08749_, _06446_, _00491_);
  and (_08750_, _06417_, _00450_);
  nor (_08751_, _08750_, _08749_);
  and (_08752_, _08751_, _08748_);
  and (_08753_, _08752_, _08745_);
  and (_08754_, _06442_, _00245_);
  and (_08755_, _06407_, _00204_);
  nor (_08756_, _08755_, _08754_);
  and (_08757_, _06424_, _00368_);
  and (_08758_, _06427_, _00327_);
  nor (_08759_, _08758_, _08757_);
  and (_08760_, _08759_, _08756_);
  and (_08761_, _06437_, _00588_);
  and (_08762_, _06440_, _00409_);
  nor (_08763_, _08762_, _08761_);
  and (_08764_, _06453_, _00050_);
  and (_08765_, _06448_, _00132_);
  nor (_08766_, _08765_, _08764_);
  and (_08767_, _08766_, _08763_);
  and (_08768_, _08767_, _08760_);
  and (_08769_, _08768_, _08753_);
  not (_08770_, _08769_);
  nor (_08771_, _08770_, _08004_);
  and (_08772_, _06453_, _00085_);
  and (_08773_, _06448_, _00198_);
  nor (_08774_, _08773_, _08772_);
  and (_08775_, _06437_, _00627_);
  and (_08776_, _06427_, _00362_);
  nor (_08777_, _08776_, _08775_);
  and (_08778_, _08777_, _08774_);
  and (_08779_, _06421_, _00578_);
  and (_08780_, _06417_, _00485_);
  nor (_08781_, _08780_, _08779_);
  and (_08782_, _06451_, _00321_);
  and (_08783_, _06407_, _00239_);
  nor (_08784_, _08783_, _08782_);
  and (_08785_, _08784_, _08781_);
  and (_08786_, _08785_, _08778_);
  and (_08787_, _06404_, _00750_);
  and (_08788_, _06412_, _00709_);
  nor (_08789_, _08788_, _08787_);
  and (_08790_, _06434_, _00668_);
  and (_08791_, _06440_, _00444_);
  nor (_08792_, _08791_, _08790_);
  and (_08793_, _08792_, _08789_);
  and (_08794_, _06446_, _00526_);
  and (_08795_, _06429_, _00126_);
  nor (_08796_, _08795_, _08794_);
  and (_08797_, _06424_, _00403_);
  and (_08798_, _06442_, _00280_);
  nor (_08799_, _08798_, _08797_);
  and (_08800_, _08799_, _08796_);
  and (_08801_, _08800_, _08793_);
  and (_08802_, _08801_, _08786_);
  and (_08803_, _08802_, _08770_);
  and (_08804_, _06404_, _00740_);
  and (_08805_, _06442_, _00270_);
  nor (_08806_, _08805_, _08804_);
  and (_08807_, _06434_, _00658_);
  and (_08808_, _06417_, _00475_);
  nor (_08809_, _08808_, _08807_);
  and (_08810_, _08809_, _08806_);
  and (_08811_, _06429_, _00116_);
  and (_08812_, _06448_, _00182_);
  nor (_08813_, _08812_, _08811_);
  and (_08814_, _06421_, _00562_);
  and (_08815_, _06407_, _00229_);
  nor (_08816_, _08815_, _08814_);
  and (_08817_, _08816_, _08813_);
  and (_08818_, _08817_, _08810_);
  and (_08819_, _06412_, _00699_);
  and (_08820_, _06437_, _00617_);
  nor (_08821_, _08820_, _08819_);
  and (_08822_, _06440_, _00434_);
  and (_08823_, _06427_, _00352_);
  nor (_08824_, _08823_, _08822_);
  and (_08825_, _08824_, _08821_);
  and (_08826_, _06446_, _00516_);
  and (_08827_, _06424_, _00393_);
  nor (_08828_, _08827_, _08826_);
  and (_08829_, _06451_, _00311_);
  and (_08830_, _06453_, _00075_);
  nor (_08831_, _08830_, _08829_);
  and (_08832_, _08831_, _08828_);
  and (_08833_, _08832_, _08825_);
  and (_08834_, _08833_, _08818_);
  and (_08835_, _06448_, _00193_);
  and (_08836_, _06429_, _00121_);
  nor (_08837_, _08836_, _08835_);
  and (_08838_, _06404_, _00745_);
  and (_08839_, _06421_, _00570_);
  nor (_08840_, _08839_, _08838_);
  and (_08841_, _08840_, _08837_);
  and (_08842_, _06446_, _00521_);
  and (_08843_, _06417_, _00480_);
  nor (_08844_, _08843_, _08842_);
  and (_08845_, _06412_, _00704_);
  and (_08846_, _06437_, _00622_);
  nor (_08847_, _08846_, _08845_);
  and (_08848_, _08847_, _08844_);
  and (_08849_, _08848_, _08841_);
  and (_08850_, _06442_, _00275_);
  and (_08851_, _06407_, _00234_);
  nor (_08852_, _08851_, _08850_);
  and (_08853_, _06427_, _00357_);
  and (_08855_, _06453_, _00080_);
  nor (_08856_, _08855_, _08853_);
  and (_08857_, _08856_, _08852_);
  and (_08858_, _06434_, _00663_);
  and (_08859_, _06440_, _00439_);
  nor (_08860_, _08859_, _08858_);
  and (_08861_, _06424_, _00398_);
  and (_08862_, _06451_, _00316_);
  nor (_08863_, _08862_, _08861_);
  and (_08864_, _08863_, _08860_);
  and (_08866_, _08864_, _08857_);
  and (_08867_, _08866_, _08849_);
  and (_08868_, _08867_, _08834_);
  and (_08869_, _08868_, _08803_);
  not (_08870_, _07018_);
  and (_08871_, _08870_, _06912_);
  not (_08872_, _06458_);
  and (_08873_, _06651_, _08872_);
  and (_08874_, _08873_, _08871_);
  and (_08875_, _08874_, _08869_);
  and (_08877_, _08875_, \oc8051_golden_model_1.TL0 [7]);
  nor (_08878_, _08867_, _08834_);
  and (_08879_, _07018_, _06912_);
  and (_08880_, _06651_, _06458_);
  and (_08881_, _08880_, _08879_);
  nor (_08882_, _08802_, _08769_);
  and (_08883_, _08882_, _08881_);
  and (_08884_, _08883_, _08878_);
  and (_08885_, _08884_, \oc8051_golden_model_1.B [7]);
  or (_08886_, _08885_, _08877_);
  not (_08888_, _08867_);
  and (_08889_, _08888_, _08834_);
  and (_08890_, _08889_, _08883_);
  and (_08891_, _08890_, \oc8051_golden_model_1.ACC [7]);
  not (_08892_, _08834_);
  and (_08893_, _08867_, _08892_);
  and (_08894_, _08893_, _08883_);
  and (_08895_, _08894_, \oc8051_golden_model_1.PSW [7]);
  or (_08896_, _08895_, _08891_);
  or (_08897_, _08896_, _08886_);
  and (_08899_, _08879_, _08873_);
  and (_08900_, _08899_, _08869_);
  and (_08901_, _08900_, \oc8051_golden_model_1.TCON [7]);
  and (_08902_, _08893_, _08803_);
  and (_08903_, _08902_, _08881_);
  and (_08904_, _08903_, \oc8051_golden_model_1.P1 [7]);
  or (_08905_, _08904_, _08901_);
  and (_08906_, _08881_, _08869_);
  and (_08907_, _08906_, \oc8051_golden_model_1.P0 [7]);
  not (_08908_, _06912_);
  and (_08910_, _07018_, _08908_);
  and (_08911_, _08910_, _08873_);
  and (_08912_, _08911_, _08869_);
  and (_08913_, _08912_, \oc8051_golden_model_1.TMOD [7]);
  or (_08914_, _08913_, _08907_);
  or (_08915_, _08914_, _08905_);
  and (_08916_, _08878_, _08803_);
  and (_08917_, _08916_, _08881_);
  and (_08918_, _08917_, \oc8051_golden_model_1.P3 [7]);
  and (_08919_, _08916_, _08899_);
  and (_08921_, _08919_, \oc8051_golden_model_1.IP [7]);
  or (_08922_, _08921_, _08918_);
  and (_08923_, _08889_, _08803_);
  and (_08924_, _08923_, _08881_);
  and (_08925_, _08924_, \oc8051_golden_model_1.P2 [7]);
  and (_08926_, _08923_, _08899_);
  and (_08927_, _08926_, \oc8051_golden_model_1.IE [7]);
  or (_08928_, _08927_, _08925_);
  or (_08929_, _08928_, _08922_);
  and (_08930_, _08902_, _08899_);
  and (_08931_, _08930_, \oc8051_golden_model_1.SCON [7]);
  and (_08932_, _08911_, _08902_);
  and (_08933_, _08932_, \oc8051_golden_model_1.SBUF [7]);
  or (_08934_, _08933_, _08931_);
  or (_08935_, _08934_, _08929_);
  or (_08936_, _08935_, _08915_);
  or (_08937_, _08936_, _08897_);
  nor (_08938_, _07018_, _06912_);
  and (_08939_, _08938_, _08869_);
  and (_08940_, _08939_, _08873_);
  and (_08941_, _08940_, \oc8051_golden_model_1.TL1 [7]);
  and (_08942_, _08880_, _08869_);
  and (_08943_, _08942_, _08871_);
  and (_08944_, _08943_, \oc8051_golden_model_1.DPL [7]);
  not (_08945_, _06651_);
  and (_08946_, _08945_, _06458_);
  and (_08947_, _08946_, _08939_);
  and (_08948_, _08947_, \oc8051_golden_model_1.PCON [7]);
  or (_08949_, _08948_, _08944_);
  or (_08950_, _08949_, _08941_);
  nor (_08951_, _06651_, _06458_);
  and (_08952_, _08951_, _08869_);
  and (_08953_, _08952_, _08879_);
  and (_08954_, _08953_, \oc8051_golden_model_1.TH0 [7]);
  and (_08955_, _08952_, _08910_);
  and (_08956_, _08955_, \oc8051_golden_model_1.TH1 [7]);
  or (_08957_, _08956_, _08954_);
  and (_08958_, _08939_, _08880_);
  and (_08959_, _08958_, \oc8051_golden_model_1.DPH [7]);
  and (_08960_, _08910_, _08942_);
  and (_08961_, _08960_, \oc8051_golden_model_1.SP [7]);
  or (_08962_, _08961_, _08959_);
  or (_08963_, _08962_, _08957_);
  or (_08964_, _08963_, _08950_);
  or (_08965_, _08964_, _08937_);
  or (_08966_, _08965_, _08771_);
  and (_08967_, _08966_, _07186_);
  and (_08968_, _06352_, _05894_);
  not (_08969_, _08968_);
  nor (_08970_, _07200_, _07520_);
  and (_08971_, _08970_, _08969_);
  and (_08972_, _08971_, _07460_);
  not (_08973_, _08972_);
  or (_08974_, _08973_, _08967_);
  or (_08975_, _08974_, _08738_);
  nor (_08976_, _08972_, _06187_);
  nor (_08977_, _08976_, _07199_);
  and (_08978_, _08977_, _08975_);
  and (_08979_, _08770_, _07199_);
  or (_08980_, _08979_, _05895_);
  or (_08981_, _08980_, _08978_);
  and (_08982_, _08711_, _05895_);
  nor (_08983_, _08982_, _07219_);
  and (_08984_, _08983_, _08981_);
  nand (_08985_, _08769_, _08006_);
  nor (_08986_, _08769_, _08006_);
  not (_08987_, _08986_);
  and (_08988_, _08987_, _08985_);
  and (_08989_, _08988_, _07219_);
  or (_08990_, _08989_, _08984_);
  and (_08991_, _08990_, _08511_);
  or (_08992_, _08991_, _08510_);
  and (_08993_, _08992_, _07215_);
  and (_08994_, _08986_, _07214_);
  or (_08995_, _08994_, _08993_);
  and (_08996_, _08995_, _07212_);
  and (_08997_, _08507_, _07211_);
  or (_08998_, _08997_, _07209_);
  or (_08999_, _08998_, _08996_);
  nor (_09000_, _08518_, _05919_);
  nor (_09001_, _09000_, _07232_);
  and (_09002_, _09001_, _08999_);
  and (_09003_, _08985_, _07232_);
  or (_09004_, _09003_, _07230_);
  or (_09005_, _09004_, _09002_);
  nand (_09006_, _08508_, _07230_);
  and (_09007_, _09006_, _05916_);
  and (_09008_, _09007_, _09005_);
  or (_09009_, _08711_, _05916_);
  or (_09010_, _07050_, _06960_);
  and (_09011_, _07492_, _05911_);
  nor (_09012_, _09011_, _09010_);
  nand (_09013_, _09012_, _09009_);
  or (_09014_, _09013_, _09008_);
  nor (_09015_, _09012_, _08571_);
  nor (_09016_, _09015_, _07238_);
  and (_09017_, _09016_, _09014_);
  and (_09018_, _08571_, _07238_);
  or (_09019_, _09018_, _07243_);
  or (_09020_, _09019_, _09017_);
  not (_09021_, _07242_);
  not (_09022_, _08671_);
  nand (_09023_, _08617_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_09024_, _08616_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_09025_, _09024_, _08625_);
  and (_09026_, _09025_, _09023_);
  nand (_09027_, _08617_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_09028_, _08616_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_09029_, _09028_, _08625_);
  and (_09030_, _09029_, _09027_);
  or (_09031_, _09030_, _09026_);
  and (_09032_, _09031_, _08607_);
  nand (_09033_, _08617_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_09034_, _08616_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_09035_, _09034_, _08625_);
  and (_09036_, _09035_, _09033_);
  nand (_09037_, _08617_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_09038_, _08616_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_09039_, _09038_, _08625_);
  and (_09040_, _09039_, _09037_);
  or (_09041_, _09040_, _09036_);
  and (_09042_, _09041_, _08635_);
  or (_09043_, _09042_, _09032_);
  nand (_09044_, _09043_, _08600_);
  nand (_09045_, _08607_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor (_09046_, _08607_, _08068_);
  nor (_09047_, _09046_, _08625_);
  nand (_09048_, _09047_, _09045_);
  nand (_09049_, _08607_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_09050_, _08607_, _08076_);
  and (_09051_, _09050_, _08625_);
  nand (_09052_, _09051_, _09049_);
  nand (_09053_, _09052_, _09048_);
  nand (_09054_, _09053_, _08616_);
  nand (_09055_, _08607_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor (_09056_, _08607_, _08060_);
  nor (_09057_, _09056_, _08625_);
  nand (_09058_, _09057_, _09055_);
  nand (_09059_, _08607_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_09060_, _08607_, _08056_);
  and (_09061_, _09060_, _08625_);
  nand (_09062_, _09061_, _09059_);
  nand (_09063_, _09062_, _09058_);
  nand (_09064_, _09063_, _08617_);
  nand (_09065_, _09064_, _09054_);
  nand (_09066_, _09065_, _08648_);
  and (_09067_, _09066_, _09044_);
  not (_09068_, _09067_);
  nand (_09069_, _08617_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_09070_, _08616_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_09071_, _09070_, _08625_);
  and (_09072_, _09071_, _09069_);
  nand (_09073_, _08617_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_09074_, _08616_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_09075_, _09074_, _08625_);
  and (_09076_, _09075_, _09073_);
  or (_09077_, _09076_, _09072_);
  and (_09078_, _09077_, _08607_);
  nand (_09079_, _08617_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_09080_, _08616_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_09081_, _09080_, _08625_);
  and (_09082_, _09081_, _09079_);
  nand (_09083_, _08617_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_09084_, _08616_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_09085_, _09084_, _08625_);
  and (_09086_, _09085_, _09083_);
  or (_09087_, _09086_, _09082_);
  and (_09088_, _09087_, _08635_);
  or (_09089_, _09088_, _09078_);
  nand (_09090_, _09089_, _08600_);
  nand (_09091_, _08607_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_09092_, _08607_, _08171_);
  nor (_09093_, _09092_, _08625_);
  nand (_09094_, _09093_, _09091_);
  nand (_09095_, _08607_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_09096_, _08607_, _08179_);
  and (_09097_, _09096_, _08625_);
  nand (_09098_, _09097_, _09095_);
  nand (_09099_, _09098_, _09094_);
  nand (_09100_, _09099_, _08616_);
  nand (_09101_, _08607_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor (_09102_, _08607_, _08163_);
  nor (_09103_, _09102_, _08625_);
  nand (_09104_, _09103_, _09101_);
  nand (_09105_, _08607_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_09106_, _08607_, _08159_);
  and (_09107_, _09106_, _08625_);
  nand (_09108_, _09107_, _09105_);
  nand (_09109_, _09108_, _09104_);
  nand (_09110_, _09109_, _08617_);
  nand (_09111_, _09110_, _09100_);
  nand (_09112_, _09111_, _08648_);
  and (_09113_, _09112_, _09090_);
  not (_09114_, _09113_);
  nand (_09115_, _08617_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_09116_, _08616_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_09117_, _09116_, _08625_);
  and (_09118_, _09117_, _09115_);
  nand (_09119_, _08617_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_09120_, _08616_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_09121_, _09120_, _08625_);
  and (_09122_, _09121_, _09119_);
  or (_09123_, _09122_, _09118_);
  and (_09124_, _09123_, _08607_);
  nand (_09125_, _08617_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_09126_, _08616_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_09127_, _09126_, _08625_);
  and (_09128_, _09127_, _09125_);
  nand (_09129_, _08617_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_09130_, _08616_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_09131_, _09130_, _08625_);
  and (_09132_, _09131_, _09129_);
  or (_09133_, _09132_, _09128_);
  and (_09134_, _09133_, _08635_);
  or (_09135_, _09134_, _09124_);
  nand (_09136_, _09135_, _08600_);
  nand (_09137_, _08607_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor (_09138_, _08607_, _08456_);
  nor (_09139_, _09138_, _08625_);
  nand (_09140_, _09139_, _09137_);
  nand (_09141_, _08607_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_09142_, _08607_, _08464_);
  and (_09143_, _09142_, _08625_);
  nand (_09144_, _09143_, _09141_);
  nand (_09145_, _09144_, _09140_);
  nand (_09146_, _09145_, _08616_);
  nand (_09147_, _08607_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor (_09148_, _08607_, _08448_);
  nor (_09149_, _09148_, _08625_);
  nand (_09150_, _09149_, _09147_);
  nand (_09151_, _08607_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_09152_, _08607_, _08444_);
  and (_09153_, _09152_, _08625_);
  nand (_09154_, _09153_, _09151_);
  nand (_09155_, _09154_, _09150_);
  nand (_09156_, _09155_, _08617_);
  nand (_09157_, _09156_, _09146_);
  nand (_09158_, _09157_, _08648_);
  and (_09159_, _09158_, _09136_);
  not (_09160_, _09159_);
  nand (_09161_, _08617_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_09162_, _08616_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor (_09163_, _09162_, _08625_);
  and (_09164_, _09163_, _09161_);
  nand (_09165_, _08617_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_09166_, _08616_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_09167_, _09166_, _08625_);
  and (_09168_, _09167_, _09165_);
  or (_09169_, _09168_, _09164_);
  and (_09170_, _09169_, _08607_);
  nand (_09171_, _08617_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_09172_, _08616_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_09173_, _09172_, _08625_);
  and (_09174_, _09173_, _09171_);
  nand (_09175_, _08617_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_09176_, _08616_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_09177_, _09176_, _08625_);
  and (_09178_, _09177_, _09175_);
  or (_09179_, _09178_, _09174_);
  and (_09180_, _09179_, _08635_);
  or (_09181_, _09180_, _09170_);
  nand (_09182_, _09181_, _08600_);
  nand (_09183_, _08607_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_09184_, _08607_, _07675_);
  nor (_09185_, _09184_, _08625_);
  nand (_09186_, _09185_, _09183_);
  nand (_09187_, _08607_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_09188_, _08607_, _07683_);
  and (_09189_, _09188_, _08625_);
  nand (_09190_, _09189_, _09187_);
  nand (_09191_, _09190_, _09186_);
  nand (_09192_, _09191_, _08616_);
  nand (_09193_, _08607_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor (_09194_, _08607_, _07667_);
  nor (_09195_, _09194_, _08625_);
  nand (_09196_, _09195_, _09193_);
  nand (_09197_, _08607_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_09198_, _08607_, _07663_);
  and (_09199_, _09198_, _08625_);
  nand (_09200_, _09199_, _09197_);
  nand (_09201_, _09200_, _09196_);
  nand (_09202_, _09201_, _08617_);
  nand (_09203_, _09202_, _09192_);
  nand (_09204_, _09203_, _08648_);
  and (_09205_, _09204_, _09182_);
  not (_09206_, _09205_);
  nand (_09207_, _08617_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_09208_, _08616_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_09209_, _09208_, _08625_);
  and (_09210_, _09209_, _09207_);
  nand (_09211_, _08617_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_09212_, _08616_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_09213_, _09212_, _08625_);
  and (_09214_, _09213_, _09211_);
  or (_09215_, _09214_, _09210_);
  and (_09216_, _09215_, _08607_);
  nand (_09217_, _08617_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_09218_, _08616_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_09219_, _09218_, _08625_);
  and (_09220_, _09219_, _09217_);
  nand (_09221_, _08617_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_09222_, _08616_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_09223_, _09222_, _08625_);
  and (_09224_, _09223_, _09221_);
  or (_09225_, _09224_, _09220_);
  and (_09226_, _09225_, _08635_);
  or (_09227_, _09226_, _09216_);
  nand (_09228_, _09227_, _08600_);
  nand (_09229_, _08607_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_09230_, _08607_, _07540_);
  nor (_09231_, _09230_, _08625_);
  nand (_09232_, _09231_, _09229_);
  nand (_09233_, _08607_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_09234_, _08607_, _07548_);
  and (_09235_, _09234_, _08625_);
  nand (_09236_, _09235_, _09233_);
  nand (_09237_, _09236_, _09232_);
  nand (_09238_, _09237_, _08616_);
  nand (_09239_, _08607_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_09240_, _08607_, _07532_);
  nor (_09241_, _09240_, _08625_);
  nand (_09242_, _09241_, _09239_);
  nand (_09243_, _08607_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_09244_, _08607_, _07528_);
  and (_09245_, _09244_, _08625_);
  nand (_09246_, _09245_, _09243_);
  nand (_09247_, _09246_, _09242_);
  nand (_09248_, _09247_, _08617_);
  nand (_09249_, _09248_, _09238_);
  nand (_09250_, _09249_, _08648_);
  and (_09251_, _09250_, _09228_);
  not (_09252_, _09251_);
  nand (_09253_, _08617_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_09254_, _08616_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor (_09255_, _09254_, _08625_);
  and (_09256_, _09255_, _09253_);
  nand (_09257_, _08617_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_09258_, _08616_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_09259_, _09258_, _08625_);
  and (_09260_, _09259_, _09257_);
  or (_09261_, _09260_, _09256_);
  and (_09262_, _09261_, _08607_);
  nand (_09263_, _08617_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_09264_, _08616_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_09265_, _09264_, _08625_);
  and (_09266_, _09265_, _09263_);
  nand (_09267_, _08617_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_09268_, _08616_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_09269_, _09268_, _08625_);
  and (_09270_, _09269_, _09267_);
  or (_09271_, _09270_, _09266_);
  and (_09272_, _09271_, _08635_);
  or (_09273_, _09272_, _09262_);
  nand (_09274_, _09273_, _08600_);
  nand (_09275_, _08607_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_09276_, _08607_, _07081_);
  nor (_09277_, _09276_, _08625_);
  nand (_09278_, _09277_, _09275_);
  nand (_09279_, _08607_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_09280_, _08607_, _07089_);
  and (_09281_, _09280_, _08625_);
  nand (_09282_, _09281_, _09279_);
  nand (_09283_, _09282_, _09278_);
  nand (_09284_, _09283_, _08616_);
  nand (_09285_, _08607_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor (_09286_, _08607_, _07071_);
  nor (_09287_, _09286_, _08625_);
  nand (_09288_, _09287_, _09285_);
  nand (_09289_, _08607_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_09290_, _08607_, _07066_);
  and (_09291_, _09290_, _08625_);
  nand (_09292_, _09291_, _09289_);
  nand (_09293_, _09292_, _09288_);
  nand (_09294_, _09293_, _08617_);
  nand (_09295_, _09294_, _09284_);
  nand (_09296_, _09295_, _08648_);
  and (_09297_, _09296_, _09274_);
  nand (_09298_, _08617_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_09299_, _08616_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor (_09300_, _09299_, _08625_);
  and (_09301_, _09300_, _09298_);
  nand (_09302_, _08617_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_09303_, _08616_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_09304_, _09303_, _08625_);
  and (_09305_, _09304_, _09302_);
  or (_09306_, _09305_, _09301_);
  and (_09307_, _09306_, _08607_);
  nand (_09308_, _08617_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_09309_, _08616_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_09310_, _09309_, _08625_);
  and (_09311_, _09310_, _09308_);
  nand (_09312_, _08617_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_09313_, _08616_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_09314_, _09313_, _08625_);
  and (_09315_, _09314_, _09312_);
  or (_09316_, _09315_, _09311_);
  and (_09317_, _09316_, _08635_);
  or (_09318_, _09317_, _09307_);
  nand (_09319_, _09318_, _08600_);
  nand (_09320_, _08607_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_09321_, _08607_, _07287_);
  nor (_09322_, _09321_, _08625_);
  nand (_09323_, _09322_, _09320_);
  nand (_09324_, _08607_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_09325_, _08607_, _07295_);
  and (_09326_, _09325_, _08625_);
  nand (_09327_, _09326_, _09324_);
  nand (_09328_, _09327_, _09323_);
  nand (_09329_, _09328_, _08616_);
  nand (_09330_, _08607_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_09331_, _08607_, _07279_);
  nor (_09332_, _09331_, _08625_);
  nand (_09333_, _09332_, _09330_);
  nand (_09334_, _08607_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_09335_, _08607_, _07275_);
  and (_09336_, _09335_, _08625_);
  nand (_09337_, _09336_, _09334_);
  nand (_09338_, _09337_, _09333_);
  nand (_09339_, _09338_, _08617_);
  nand (_09340_, _09339_, _09329_);
  nand (_09341_, _09340_, _08648_);
  and (_09342_, _09341_, _09319_);
  nor (_09343_, _09342_, _09297_);
  and (_09344_, _09343_, _09252_);
  and (_09345_, _09344_, _09206_);
  and (_09346_, _09345_, _09160_);
  and (_09347_, _09346_, _09114_);
  and (_09348_, _09347_, _09068_);
  nor (_09349_, _09348_, _09022_);
  and (_09350_, _09348_, _09022_);
  or (_09351_, _09350_, _09349_);
  or (_09352_, _09351_, _07403_);
  and (_09353_, _09352_, _09021_);
  and (_09354_, _09353_, _09020_);
  and (_09355_, _08685_, _07242_);
  or (_09356_, _09355_, _09354_);
  and (_09357_, _09356_, _08505_);
  nor (_09358_, _05592_, _05552_);
  and (_09359_, _09358_, \oc8051_golden_model_1.PC [3]);
  and (_09360_, _09359_, _08514_);
  and (_09361_, _09360_, \oc8051_golden_model_1.PC [7]);
  nor (_09362_, _09360_, \oc8051_golden_model_1.PC [7]);
  nor (_09363_, _09362_, _09361_);
  and (_09364_, _09363_, _06378_);
  or (_09365_, _09364_, _09357_);
  and (_09366_, _09365_, _05913_);
  and (_09367_, _08518_, _05912_);
  or (_09368_, _09367_, _09366_);
  and (_09369_, _09368_, _07265_);
  and (_09370_, _08698_, _07249_);
  nor (_09371_, _07653_, _07433_);
  not (_09372_, _09371_);
  nor (_09373_, _09372_, _09370_);
  not (_09374_, _09373_);
  nor (_09375_, _09374_, _09369_);
  not (_09376_, _08106_);
  not (_09377_, _08209_);
  not (_09378_, _08494_);
  not (_09379_, _07713_);
  not (_09380_, _07578_);
  not (_09381_, _07120_);
  and (_09382_, _09381_, _07325_);
  and (_09383_, _09382_, _09380_);
  and (_09384_, _09383_, _09379_);
  and (_09385_, _09384_, _09378_);
  and (_09386_, _09385_, _09377_);
  and (_09387_, _09386_, _09376_);
  and (_09388_, _09387_, _08562_);
  nor (_09389_, _09387_, _08562_);
  nor (_09390_, _09389_, _09388_);
  nor (_09391_, _09390_, _09371_);
  nor (_09392_, _09391_, _09375_);
  nor (_09393_, _09392_, _07259_);
  and (_09394_, _09342_, _09297_);
  and (_09395_, _09394_, _09251_);
  and (_09396_, _09395_, _09205_);
  and (_09397_, _09396_, _09159_);
  and (_09398_, _09397_, _09113_);
  and (_09399_, _09398_, _09067_);
  nor (_09400_, _09399_, _09022_);
  and (_09401_, _09399_, _09022_);
  or (_09402_, _09401_, _09400_);
  nor (_09403_, _09402_, _07414_);
  nor (_09404_, _09403_, _06190_);
  not (_09405_, _09404_);
  nor (_09406_, _09405_, _09393_);
  nor (_09407_, _09406_, _08504_);
  nor (_09408_, _09407_, _07508_);
  or (_09409_, _09408_, _07850_);
  and (_09410_, _09409_, _07849_);
  and (_09411_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_09412_, _09411_, \oc8051_golden_model_1.PC [10]);
  and (_09413_, _09412_, _09361_);
  and (_09414_, _09413_, \oc8051_golden_model_1.PC [11]);
  and (_09415_, _09414_, \oc8051_golden_model_1.PC [12]);
  and (_09416_, _09415_, \oc8051_golden_model_1.PC [13]);
  and (_09417_, _09416_, \oc8051_golden_model_1.PC [14]);
  nor (_09418_, _09417_, \oc8051_golden_model_1.PC [15]);
  and (_09419_, _09361_, \oc8051_golden_model_1.PC [8]);
  and (_09420_, _09419_, \oc8051_golden_model_1.PC [9]);
  and (_09421_, _09420_, \oc8051_golden_model_1.PC [10]);
  and (_09422_, _09421_, \oc8051_golden_model_1.PC [11]);
  and (_09423_, _09422_, \oc8051_golden_model_1.PC [12]);
  and (_09424_, _09423_, \oc8051_golden_model_1.PC [13]);
  and (_09425_, _09424_, \oc8051_golden_model_1.PC [14]);
  and (_09426_, _09425_, \oc8051_golden_model_1.PC [15]);
  nor (_09427_, _09426_, _09418_);
  or (_09428_, _09427_, _08505_);
  and (_09429_, _09412_, _08516_);
  and (_09430_, _09429_, \oc8051_golden_model_1.PC [11]);
  and (_09431_, _09430_, \oc8051_golden_model_1.PC [12]);
  and (_09432_, _09431_, \oc8051_golden_model_1.PC [13]);
  and (_09433_, _09432_, \oc8051_golden_model_1.PC [14]);
  nor (_09434_, _09433_, \oc8051_golden_model_1.PC [15]);
  and (_09435_, _08516_, \oc8051_golden_model_1.PC [8]);
  and (_09436_, _09435_, \oc8051_golden_model_1.PC [9]);
  and (_09437_, _09436_, \oc8051_golden_model_1.PC [10]);
  and (_09438_, _09437_, \oc8051_golden_model_1.PC [11]);
  and (_09439_, _09438_, \oc8051_golden_model_1.PC [12]);
  and (_09440_, _09439_, \oc8051_golden_model_1.PC [13]);
  and (_09441_, _09440_, \oc8051_golden_model_1.PC [14]);
  and (_09442_, _09441_, \oc8051_golden_model_1.PC [15]);
  nor (_09443_, _09442_, _09434_);
  or (_09444_, _09443_, _06378_);
  and (_09445_, _09444_, _09428_);
  and (_09446_, _09445_, _07844_);
  and (_09447_, _09446_, _07847_);
  or (_41177_, _09447_, _09410_);
  not (_09448_, \oc8051_golden_model_1.B [7]);
  nor (_09449_, _01452_, _09448_);
  nor (_09450_, _07911_, _09448_);
  and (_09451_, _08509_, _07911_);
  or (_09452_, _09451_, _09450_);
  and (_09453_, _09452_, _06533_);
  not (_09454_, _07911_);
  nor (_09455_, _08004_, _09454_);
  or (_09456_, _09455_, _09450_);
  or (_09457_, _09456_, _07188_);
  or (_09458_, _09456_, _07142_);
  and (_09459_, _08685_, _07911_);
  or (_09460_, _09459_, _09450_);
  or (_09461_, _09460_, _06252_);
  and (_09462_, _07911_, \oc8051_golden_model_1.ACC [7]);
  or (_09463_, _09462_, _09450_);
  and (_09464_, _09463_, _07123_);
  nor (_09465_, _07123_, _09448_);
  or (_09466_, _09465_, _06251_);
  or (_09467_, _09466_, _09464_);
  and (_09468_, _09467_, _06476_);
  and (_09469_, _09468_, _09461_);
  nor (_09471_, _08547_, _09448_);
  and (_09472_, _08560_, _08547_);
  or (_09473_, _09472_, _09471_);
  and (_09474_, _09473_, _06475_);
  or (_09475_, _09474_, _06468_);
  or (_09476_, _09475_, _09469_);
  and (_09477_, _09476_, _09458_);
  or (_09478_, _09477_, _06466_);
  or (_09479_, _09463_, _06801_);
  and (_09480_, _09479_, _06484_);
  and (_09481_, _09480_, _09478_);
  and (_09482_, _08698_, _08547_);
  or (_09483_, _09482_, _09471_);
  and (_09484_, _09483_, _06483_);
  or (_09485_, _09484_, _09481_);
  and (_09486_, _09485_, _07164_);
  and (_09487_, _06372_, _06490_);
  or (_09488_, _09471_, _08706_);
  and (_09489_, _09488_, _06461_);
  and (_09490_, _09489_, _09473_);
  or (_09492_, _09490_, _09487_);
  or (_09493_, _09492_, _09486_);
  not (_09494_, _09487_);
  and (_09495_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_09496_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_09497_, _09496_, _09495_);
  and (_09498_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and (_09499_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and (_09500_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_09501_, _09500_, _09499_);
  nor (_09502_, _09501_, _09497_);
  and (_09503_, _09502_, _09498_);
  nor (_09504_, _09503_, _09497_);
  and (_09505_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_09506_, _09505_, _09499_);
  and (_09507_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_09508_, _09507_, _09495_);
  nor (_09509_, _09508_, _09506_);
  not (_09510_, _09509_);
  nor (_09511_, _09510_, _09504_);
  and (_09512_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_09513_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and (_09514_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and (_09515_, _09514_, _09513_);
  nor (_09516_, _09514_, _09513_);
  nor (_09517_, _09516_, _09515_);
  and (_09518_, _09517_, _09512_);
  nor (_09519_, _09517_, _09512_);
  nor (_09520_, _09519_, _09518_);
  and (_09521_, _09510_, _09504_);
  nor (_09522_, _09521_, _09511_);
  and (_09523_, _09522_, _09520_);
  nor (_09524_, _09523_, _09511_);
  not (_09525_, _09499_);
  and (_09526_, _09505_, _09525_);
  and (_09527_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and (_09528_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_09529_, _09528_, _09513_);
  and (_09530_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  and (_09531_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_09532_, _09531_, _09530_);
  nor (_09533_, _09532_, _09529_);
  and (_09534_, _09533_, _09527_);
  nor (_09535_, _09533_, _09527_);
  nor (_09536_, _09535_, _09534_);
  and (_09537_, _09536_, _09526_);
  nor (_09538_, _09536_, _09526_);
  nor (_09539_, _09538_, _09537_);
  not (_09540_, _09539_);
  nor (_09541_, _09540_, _09524_);
  and (_09542_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_09543_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and (_09544_, _09543_, _09542_);
  nor (_09545_, _09518_, _09515_);
  and (_09546_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and (_09547_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_09548_, _09547_, _09546_);
  nor (_09549_, _09547_, _09546_);
  nor (_09550_, _09549_, _09548_);
  not (_09551_, _09550_);
  nor (_09552_, _09551_, _09545_);
  and (_09553_, _09551_, _09545_);
  nor (_09554_, _09553_, _09552_);
  and (_09555_, _09554_, _09544_);
  nor (_09556_, _09554_, _09544_);
  nor (_09557_, _09556_, _09555_);
  and (_09558_, _09540_, _09524_);
  nor (_09559_, _09558_, _09541_);
  and (_09560_, _09559_, _09557_);
  nor (_09561_, _09560_, _09541_);
  nor (_09562_, _09534_, _09529_);
  and (_09563_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and (_09564_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and (_09565_, _09564_, _09563_);
  nor (_09566_, _09564_, _09563_);
  nor (_09567_, _09566_, _09565_);
  not (_09568_, _09567_);
  nor (_09569_, _09568_, _09562_);
  and (_09570_, _09568_, _09562_);
  nor (_09571_, _09570_, _09569_);
  and (_09572_, _09571_, _09548_);
  nor (_09573_, _09571_, _09548_);
  nor (_09574_, _09573_, _09572_);
  nor (_09575_, _09537_, _09506_);
  and (_09576_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  and (_09577_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_09578_, _09577_, _09528_);
  nor (_09579_, _09577_, _09528_);
  nor (_09580_, _09579_, _09578_);
  and (_09581_, _09580_, _09576_);
  nor (_09582_, _09580_, _09576_);
  nor (_09583_, _09582_, _09581_);
  not (_09584_, _09583_);
  nor (_09585_, _09584_, _09575_);
  and (_09586_, _09584_, _09575_);
  nor (_09587_, _09586_, _09585_);
  and (_09588_, _09587_, _09574_);
  nor (_09589_, _09587_, _09574_);
  nor (_09590_, _09589_, _09588_);
  not (_09591_, _09590_);
  nor (_09592_, _09591_, _09561_);
  nor (_09593_, _09555_, _09552_);
  not (_09594_, _09593_);
  and (_09595_, _09591_, _09561_);
  nor (_09596_, _09595_, _09592_);
  and (_09597_, _09596_, _09594_);
  nor (_09598_, _09597_, _09592_);
  nor (_09599_, _09572_, _09569_);
  not (_09600_, _09599_);
  nor (_09601_, _09588_, _09585_);
  not (_09602_, _09601_);
  and (_09603_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_09604_, _09603_, _09528_);
  and (_09605_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_09606_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_09607_, _09606_, _09605_);
  nor (_09608_, _09607_, _09604_);
  nor (_09609_, _09581_, _09578_);
  and (_09610_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and (_09611_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and (_09612_, _09611_, _09610_);
  nor (_09613_, _09611_, _09610_);
  nor (_09614_, _09613_, _09612_);
  not (_09615_, _09614_);
  nor (_09616_, _09615_, _09609_);
  and (_09617_, _09615_, _09609_);
  nor (_09618_, _09617_, _09616_);
  and (_09619_, _09618_, _09565_);
  nor (_09620_, _09618_, _09565_);
  nor (_09621_, _09620_, _09619_);
  and (_09622_, _09621_, _09608_);
  nor (_09623_, _09621_, _09608_);
  nor (_09624_, _09623_, _09622_);
  and (_09625_, _09624_, _09602_);
  nor (_09626_, _09624_, _09602_);
  nor (_09627_, _09626_, _09625_);
  and (_09628_, _09627_, _09600_);
  nor (_09629_, _09627_, _09600_);
  nor (_09630_, _09629_, _09628_);
  not (_09631_, _09630_);
  nor (_09632_, _09631_, _09598_);
  nor (_09633_, _09628_, _09625_);
  nor (_09634_, _09619_, _09616_);
  not (_09635_, _09634_);
  and (_09636_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and (_09637_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_09638_, _09637_, _09636_);
  nor (_09639_, _09637_, _09636_);
  nor (_09640_, _09639_, _09638_);
  and (_09641_, _09640_, _09604_);
  nor (_09642_, _09640_, _09604_);
  nor (_09643_, _09642_, _09641_);
  and (_09644_, _09643_, _09612_);
  nor (_09645_, _09643_, _09612_);
  nor (_09647_, _09645_, _09644_);
  and (_09648_, _09647_, _09603_);
  nor (_09650_, _09647_, _09603_);
  nor (_09651_, _09650_, _09648_);
  and (_09653_, _09651_, _09622_);
  nor (_09654_, _09651_, _09622_);
  nor (_09656_, _09654_, _09653_);
  and (_09657_, _09656_, _09635_);
  nor (_09659_, _09656_, _09635_);
  nor (_09660_, _09659_, _09657_);
  not (_09662_, _09660_);
  nor (_09663_, _09662_, _09633_);
  and (_09665_, _09662_, _09633_);
  nor (_09666_, _09665_, _09663_);
  and (_09668_, _09666_, _09632_);
  nor (_09669_, _09657_, _09653_);
  nor (_09671_, _09644_, _09641_);
  not (_09672_, _09671_);
  and (_09674_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and (_09675_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_09677_, _09675_, _09674_);
  nor (_09678_, _09675_, _09674_);
  nor (_09680_, _09678_, _09677_);
  and (_09681_, _09680_, _09638_);
  nor (_09683_, _09680_, _09638_);
  nor (_09684_, _09683_, _09681_);
  and (_09685_, _09684_, _09648_);
  nor (_09686_, _09684_, _09648_);
  nor (_09687_, _09686_, _09685_);
  and (_09688_, _09687_, _09672_);
  nor (_09689_, _09687_, _09672_);
  nor (_09690_, _09689_, _09688_);
  not (_09691_, _09690_);
  nor (_09692_, _09691_, _09669_);
  and (_09693_, _09691_, _09669_);
  nor (_09694_, _09693_, _09692_);
  and (_09695_, _09694_, _09663_);
  nor (_09696_, _09694_, _09663_);
  nor (_09697_, _09696_, _09695_);
  and (_09698_, _09697_, _09668_);
  nor (_09699_, _09697_, _09668_);
  nor (_09700_, _09699_, _09698_);
  and (_09701_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and (_09702_, _09701_, _09499_);
  and (_09703_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and (_09704_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor (_09705_, _09704_, _09496_);
  nor (_09706_, _09705_, _09702_);
  and (_09707_, _09706_, _09703_);
  nor (_09708_, _09707_, _09702_);
  not (_09709_, _09708_);
  nor (_09710_, _09502_, _09498_);
  nor (_09711_, _09710_, _09503_);
  and (_09712_, _09711_, _09709_);
  and (_09713_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_09714_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and (_09715_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_09716_, _09715_, _09714_);
  nor (_09717_, _09715_, _09714_);
  nor (_09718_, _09717_, _09716_);
  and (_09719_, _09718_, _09713_);
  nor (_09720_, _09718_, _09713_);
  nor (_09721_, _09720_, _09719_);
  nor (_09722_, _09711_, _09709_);
  nor (_09723_, _09722_, _09712_);
  and (_09724_, _09723_, _09721_);
  nor (_09725_, _09724_, _09712_);
  nor (_09726_, _09522_, _09520_);
  nor (_09727_, _09726_, _09523_);
  not (_09728_, _09727_);
  nor (_09729_, _09728_, _09725_);
  and (_09730_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_09731_, _09730_, _09543_);
  nor (_09732_, _09719_, _09716_);
  nor (_09733_, _09543_, _09542_);
  nor (_09734_, _09733_, _09544_);
  not (_09735_, _09734_);
  nor (_09736_, _09735_, _09732_);
  and (_09737_, _09735_, _09732_);
  nor (_09738_, _09737_, _09736_);
  and (_09739_, _09738_, _09731_);
  nor (_09740_, _09738_, _09731_);
  nor (_09742_, _09740_, _09739_);
  and (_09744_, _09728_, _09725_);
  nor (_09745_, _09744_, _09729_);
  and (_09747_, _09745_, _09742_);
  nor (_09748_, _09747_, _09729_);
  nor (_09750_, _09559_, _09557_);
  nor (_09751_, _09750_, _09560_);
  not (_09753_, _09751_);
  nor (_09754_, _09753_, _09748_);
  nor (_09756_, _09739_, _09736_);
  not (_09757_, _09756_);
  and (_09759_, _09753_, _09748_);
  nor (_09760_, _09759_, _09754_);
  and (_09762_, _09760_, _09757_);
  nor (_09763_, _09762_, _09754_);
  nor (_09765_, _09596_, _09594_);
  nor (_09766_, _09765_, _09597_);
  not (_09768_, _09766_);
  nor (_09769_, _09768_, _09763_);
  and (_09771_, _09631_, _09598_);
  nor (_09772_, _09771_, _09632_);
  and (_09774_, _09772_, _09769_);
  nor (_09775_, _09666_, _09632_);
  nor (_09777_, _09775_, _09668_);
  nand (_09778_, _09777_, _09774_);
  and (_09779_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and (_09780_, _09779_, _09701_);
  and (_09781_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_09782_, _09779_, _09701_);
  nor (_09783_, _09782_, _09780_);
  and (_09784_, _09783_, _09781_);
  nor (_09785_, _09784_, _09780_);
  not (_09786_, _09785_);
  nor (_09787_, _09706_, _09703_);
  nor (_09788_, _09787_, _09707_);
  and (_09789_, _09788_, _09786_);
  and (_09790_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and (_09791_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_09792_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_09793_, _09792_, _09791_);
  nor (_09794_, _09792_, _09791_);
  nor (_09795_, _09794_, _09793_);
  and (_09796_, _09795_, _09790_);
  nor (_09797_, _09795_, _09790_);
  nor (_09798_, _09797_, _09796_);
  nor (_09799_, _09788_, _09786_);
  nor (_09800_, _09799_, _09789_);
  and (_09801_, _09800_, _09798_);
  nor (_09802_, _09801_, _09789_);
  not (_09803_, _09802_);
  nor (_09804_, _09723_, _09721_);
  nor (_09805_, _09804_, _09724_);
  and (_09806_, _09805_, _09803_);
  nor (_09807_, _09796_, _09793_);
  and (_09808_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and (_09809_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor (_09810_, _09809_, _09808_);
  nor (_09811_, _09810_, _09731_);
  not (_09812_, _09811_);
  nor (_09813_, _09812_, _09807_);
  and (_09814_, _09812_, _09807_);
  nor (_09815_, _09814_, _09813_);
  nor (_09816_, _09805_, _09803_);
  nor (_09817_, _09816_, _09806_);
  and (_09818_, _09817_, _09815_);
  nor (_09819_, _09818_, _09806_);
  nor (_09820_, _09745_, _09742_);
  nor (_09821_, _09820_, _09747_);
  not (_09822_, _09821_);
  nor (_09823_, _09822_, _09819_);
  and (_09824_, _09822_, _09819_);
  nor (_09825_, _09824_, _09823_);
  and (_09826_, _09825_, _09813_);
  nor (_09827_, _09826_, _09823_);
  nor (_09828_, _09760_, _09757_);
  nor (_09829_, _09828_, _09762_);
  not (_09830_, _09829_);
  nor (_09831_, _09830_, _09827_);
  and (_09832_, _09768_, _09763_);
  nor (_09833_, _09832_, _09769_);
  and (_09834_, _09833_, _09831_);
  nor (_09835_, _09772_, _09769_);
  nor (_09836_, _09835_, _09774_);
  and (_09837_, _09836_, _09834_);
  nor (_09838_, _09836_, _09834_);
  nor (_09839_, _09838_, _09837_);
  and (_09840_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and (_09841_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_09842_, _09841_, _09840_);
  and (_09843_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_09844_, _09841_, _09840_);
  nor (_09845_, _09844_, _09842_);
  and (_09846_, _09845_, _09843_);
  nor (_09847_, _09846_, _09842_);
  not (_09848_, _09847_);
  nor (_09849_, _09783_, _09781_);
  nor (_09850_, _09849_, _09784_);
  and (_09851_, _09850_, _09848_);
  and (_09852_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_09853_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_09854_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and (_09855_, _09854_, _09853_);
  nor (_09856_, _09854_, _09853_);
  nor (_09857_, _09856_, _09855_);
  and (_09858_, _09857_, _09852_);
  nor (_09859_, _09857_, _09852_);
  nor (_09860_, _09859_, _09858_);
  nor (_09861_, _09850_, _09848_);
  nor (_09862_, _09861_, _09851_);
  and (_09863_, _09862_, _09860_);
  nor (_09864_, _09863_, _09851_);
  not (_09865_, _09864_);
  nor (_09866_, _09800_, _09798_);
  nor (_09867_, _09866_, _09801_);
  and (_09868_, _09867_, _09865_);
  not (_09869_, _09730_);
  nor (_09870_, _09858_, _09855_);
  nor (_09871_, _09870_, _09869_);
  and (_09872_, _09870_, _09869_);
  nor (_09873_, _09872_, _09871_);
  nor (_09874_, _09867_, _09865_);
  nor (_09875_, _09874_, _09868_);
  and (_09876_, _09875_, _09873_);
  nor (_09877_, _09876_, _09868_);
  not (_09878_, _09877_);
  nor (_09879_, _09817_, _09815_);
  nor (_09880_, _09879_, _09818_);
  and (_09881_, _09880_, _09878_);
  nor (_09882_, _09880_, _09878_);
  nor (_09883_, _09882_, _09881_);
  and (_09884_, _09883_, _09871_);
  nor (_09885_, _09884_, _09881_);
  nor (_09886_, _09825_, _09813_);
  nor (_09887_, _09886_, _09826_);
  not (_09888_, _09887_);
  nor (_09889_, _09888_, _09885_);
  and (_09890_, _09830_, _09827_);
  nor (_09891_, _09890_, _09831_);
  and (_09892_, _09891_, _09889_);
  nor (_09893_, _09833_, _09831_);
  nor (_09894_, _09893_, _09834_);
  nand (_09895_, _09894_, _09892_);
  or (_09896_, _09894_, _09892_);
  and (_09897_, _09896_, _09895_);
  and (_09898_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_09899_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_09900_, _09899_, _09898_);
  and (_09901_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor (_09902_, _09899_, _09898_);
  nor (_09903_, _09902_, _09900_);
  and (_09904_, _09903_, _09901_);
  nor (_09905_, _09904_, _09900_);
  not (_09906_, _09905_);
  nor (_09907_, _09845_, _09843_);
  nor (_09908_, _09907_, _09846_);
  and (_09909_, _09908_, _09906_);
  and (_09910_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_09911_, _09910_, _09854_);
  and (_09912_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and (_09913_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_09914_, _09913_, _09912_);
  nor (_09915_, _09914_, _09911_);
  nor (_09916_, _09908_, _09906_);
  nor (_09917_, _09916_, _09909_);
  and (_09918_, _09917_, _09915_);
  nor (_09919_, _09918_, _09909_);
  not (_09920_, _09919_);
  nor (_09921_, _09862_, _09860_);
  nor (_09922_, _09921_, _09863_);
  and (_09923_, _09922_, _09920_);
  nor (_09924_, _09922_, _09920_);
  nor (_09925_, _09924_, _09923_);
  and (_09926_, _09925_, _09911_);
  nor (_09927_, _09926_, _09923_);
  not (_09928_, _09927_);
  nor (_09929_, _09875_, _09873_);
  nor (_09930_, _09929_, _09876_);
  and (_09931_, _09930_, _09928_);
  nor (_09932_, _09883_, _09871_);
  nor (_09933_, _09932_, _09884_);
  and (_09934_, _09933_, _09931_);
  and (_09935_, _09888_, _09885_);
  nor (_09936_, _09935_, _09889_);
  and (_09937_, _09936_, _09934_);
  nor (_09938_, _09891_, _09889_);
  nor (_09939_, _09938_, _09892_);
  nor (_09940_, _09939_, _09937_);
  and (_09941_, _09939_, _09937_);
  not (_09942_, _09941_);
  and (_09943_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_09944_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and (_09945_, _09944_, _09943_);
  and (_09946_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_09947_, _09944_, _09943_);
  nor (_09948_, _09947_, _09945_);
  and (_09949_, _09948_, _09946_);
  nor (_09950_, _09949_, _09945_);
  not (_09951_, _09950_);
  nor (_09952_, _09903_, _09901_);
  nor (_09953_, _09952_, _09904_);
  and (_09954_, _09953_, _09951_);
  nor (_09955_, _09953_, _09951_);
  nor (_09956_, _09955_, _09954_);
  and (_09957_, _09956_, _09910_);
  nor (_09958_, _09957_, _09954_);
  not (_09959_, _09958_);
  nor (_09960_, _09917_, _09915_);
  nor (_09961_, _09960_, _09918_);
  and (_09962_, _09961_, _09959_);
  nor (_09963_, _09925_, _09911_);
  nor (_09964_, _09963_, _09926_);
  and (_09965_, _09964_, _09962_);
  nor (_09966_, _09930_, _09928_);
  nor (_09967_, _09966_, _09931_);
  and (_09968_, _09967_, _09965_);
  nor (_09969_, _09933_, _09931_);
  nor (_09970_, _09969_, _09934_);
  and (_09971_, _09970_, _09968_);
  nor (_09972_, _09936_, _09934_);
  nor (_09973_, _09972_, _09937_);
  and (_09974_, _09973_, _09971_);
  and (_09975_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and (_09976_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and (_09977_, _09976_, _09975_);
  nor (_09978_, _09948_, _09946_);
  nor (_09979_, _09978_, _09949_);
  and (_09980_, _09979_, _09977_);
  nor (_09981_, _09956_, _09910_);
  nor (_09982_, _09981_, _09957_);
  and (_09983_, _09982_, _09980_);
  nor (_09984_, _09961_, _09959_);
  nor (_09985_, _09984_, _09962_);
  and (_09986_, _09985_, _09983_);
  nor (_09987_, _09964_, _09962_);
  nor (_09988_, _09987_, _09965_);
  and (_09989_, _09988_, _09986_);
  nor (_09990_, _09967_, _09965_);
  nor (_09991_, _09990_, _09968_);
  and (_09992_, _09991_, _09989_);
  nor (_09993_, _09970_, _09968_);
  nor (_09994_, _09993_, _09971_);
  and (_09995_, _09994_, _09992_);
  nor (_09996_, _09973_, _09971_);
  nor (_09997_, _09996_, _09974_);
  and (_09998_, _09997_, _09995_);
  nor (_09999_, _09998_, _09974_);
  and (_10000_, _09999_, _09942_);
  nor (_10001_, _10000_, _09940_);
  nand (_10002_, _10001_, _09897_);
  and (_10003_, _10002_, _09895_);
  not (_10004_, _10003_);
  and (_10005_, _10004_, _09839_);
  or (_10006_, _10005_, _09837_);
  or (_10007_, _09777_, _09774_);
  and (_10008_, _10007_, _09778_);
  nand (_10009_, _10008_, _10006_);
  and (_10010_, _10009_, _09778_);
  not (_10011_, _10010_);
  and (_10012_, _10011_, _09700_);
  or (_10013_, _10012_, _09698_);
  and (_10014_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not (_10015_, _10014_);
  nor (_10016_, _10015_, _09637_);
  nor (_10017_, _10016_, _09681_);
  nor (_10018_, _09688_, _09685_);
  nor (_10019_, _10018_, _10017_);
  and (_10020_, _10018_, _10017_);
  nor (_10021_, _10020_, _10019_);
  nor (_10022_, _09695_, _09692_);
  not (_10023_, _10022_);
  and (_10024_, _10023_, _10021_);
  nor (_10025_, _10023_, _10021_);
  nor (_10026_, _10025_, _10024_);
  and (_10027_, _10026_, _10013_);
  or (_10028_, _10019_, _09677_);
  or (_10029_, _10028_, _10024_);
  or (_10030_, _10029_, _10027_);
  or (_10031_, _10030_, _09494_);
  and (_10032_, _10031_, _06242_);
  and (_10033_, _10032_, _09493_);
  and (_10034_, _08726_, _08547_);
  or (_10035_, _10034_, _09471_);
  and (_10036_, _10035_, _06241_);
  or (_10037_, _10036_, _07187_);
  or (_10038_, _10037_, _10033_);
  and (_10039_, _10038_, _09457_);
  or (_10040_, _10039_, _07182_);
  and (_10041_, _08671_, _07911_);
  or (_10042_, _09450_, _07183_);
  or (_10043_, _10042_, _10041_);
  and (_10044_, _10043_, _06336_);
  and (_10045_, _10044_, _10040_);
  and (_10046_, _06372_, _05899_);
  and (_10047_, _08966_, _07911_);
  or (_10048_, _10047_, _09450_);
  and (_10049_, _10048_, _05968_);
  or (_10050_, _10049_, _10046_);
  or (_10051_, _10050_, _10045_);
  not (_10052_, _10046_);
  not (_10053_, \oc8051_golden_model_1.B [1]);
  nor (_10054_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_10055_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and (_10056_, _10055_, _10054_);
  and (_10057_, _10056_, _10053_);
  not (_10058_, \oc8051_golden_model_1.B [0]);
  and (_10059_, _10058_, \oc8051_golden_model_1.ACC [7]);
  nor (_10060_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_10061_, _10060_, _10059_);
  and (_10062_, _10061_, _10057_);
  and (_10063_, \oc8051_golden_model_1.B [0], _08506_);
  not (_10064_, _10063_);
  and (_10065_, _10060_, _10057_);
  and (_10066_, _10065_, _10064_);
  or (_10067_, _10066_, _08506_);
  not (_10068_, \oc8051_golden_model_1.ACC [6]);
  and (_10069_, \oc8051_golden_model_1.B [0], _10068_);
  nor (_10070_, _10069_, _08506_);
  nor (_10071_, _10070_, _10053_);
  not (_10072_, _10071_);
  and (_10073_, _10060_, _10056_);
  and (_10074_, _10073_, _10072_);
  nor (_10075_, _10074_, _10067_);
  nor (_10076_, _10075_, _10062_);
  and (_10077_, _10074_, \oc8051_golden_model_1.B [0]);
  nor (_10078_, _10077_, _10068_);
  and (_10079_, _10078_, _10053_);
  nor (_10080_, _10078_, _10053_);
  nor (_10081_, _10080_, _10079_);
  nor (_10082_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor (_10083_, _10082_, _09701_);
  nor (_10084_, _10083_, \oc8051_golden_model_1.ACC [4]);
  and (_10085_, \oc8051_golden_model_1.ACC [4], _10058_);
  nor (_10086_, _10085_, \oc8051_golden_model_1.ACC [5]);
  not (_10087_, \oc8051_golden_model_1.ACC [4]);
  and (_10088_, _10087_, \oc8051_golden_model_1.B [0]);
  nor (_10089_, _10088_, _10086_);
  nor (_10090_, _10089_, _10084_);
  not (_10091_, _10090_);
  and (_10092_, _10091_, _10081_);
  nor (_10093_, _10076_, \oc8051_golden_model_1.B [2]);
  nor (_10094_, _10093_, _10079_);
  not (_10095_, _10094_);
  nor (_10096_, _10095_, _10092_);
  not (_10097_, \oc8051_golden_model_1.B [3]);
  nor (_10098_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_10099_, _10098_, _10054_);
  and (_10100_, _10099_, _10097_);
  and (_10101_, \oc8051_golden_model_1.B [2], _08506_);
  not (_10102_, _10101_);
  and (_10103_, _10102_, _10100_);
  not (_10104_, _10103_);
  nor (_10105_, _10104_, _10096_);
  nor (_10106_, _10105_, _10076_);
  nor (_10107_, _10106_, _10062_);
  and (_10108_, _10099_, \oc8051_golden_model_1.ACC [7]);
  nor (_10109_, _10108_, _10100_);
  nor (_10110_, _10107_, \oc8051_golden_model_1.B [3]);
  not (_10111_, \oc8051_golden_model_1.B [2]);
  nor (_10112_, _10091_, _10081_);
  nor (_10113_, _10112_, _10092_);
  not (_10114_, _10113_);
  and (_10115_, _10114_, _10105_);
  nor (_10116_, _10105_, _10078_);
  nor (_10117_, _10116_, _10115_);
  and (_10118_, _10117_, _10111_);
  nor (_10119_, _10117_, _10111_);
  nor (_10120_, _10119_, _10118_);
  not (_10121_, _10120_);
  not (_10122_, \oc8051_golden_model_1.ACC [5]);
  nor (_10123_, _10105_, _10122_);
  and (_10124_, _10105_, _10083_);
  or (_10125_, _10124_, _10123_);
  and (_10126_, _10125_, _10053_);
  nor (_10127_, _10125_, _10053_);
  nor (_10128_, _10127_, _10088_);
  nor (_10129_, _10128_, _10126_);
  nor (_10130_, _10129_, _10121_);
  or (_10131_, _10130_, _10118_);
  nor (_10132_, _10131_, _10110_);
  nor (_10133_, _10132_, _10109_);
  nor (_10134_, _10133_, _10107_);
  nor (_10135_, _10134_, _10062_);
  not (_10136_, _10133_);
  and (_10137_, _10129_, _10121_);
  nor (_10138_, _10137_, _10130_);
  nor (_10139_, _10138_, _10136_);
  nor (_10140_, _10133_, _10117_);
  nor (_10141_, _10140_, _10139_);
  and (_10142_, _10141_, _10097_);
  nor (_10143_, _10141_, _10097_);
  nor (_10144_, _10143_, _10142_);
  not (_10145_, _10144_);
  nor (_10146_, _10133_, _10125_);
  nor (_10147_, _10127_, _10126_);
  and (_10148_, _10147_, _10088_);
  nor (_10149_, _10147_, _10088_);
  nor (_10150_, _10149_, _10148_);
  and (_10151_, _10150_, _10133_);
  or (_10152_, _10151_, _10146_);
  nor (_10153_, _10152_, \oc8051_golden_model_1.B [2]);
  and (_10154_, _10152_, \oc8051_golden_model_1.B [2]);
  nor (_10155_, _10088_, _10085_);
  and (_10156_, _10133_, _10155_);
  nor (_10157_, _10133_, \oc8051_golden_model_1.ACC [4]);
  nor (_10158_, _10157_, _10156_);
  and (_10159_, _10158_, _10053_);
  nor (_10160_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_10161_, _10160_, _09898_);
  nor (_10162_, _10161_, \oc8051_golden_model_1.ACC [2]);
  and (_10163_, _10058_, \oc8051_golden_model_1.ACC [2]);
  nor (_10164_, _10163_, \oc8051_golden_model_1.ACC [3]);
  not (_10165_, \oc8051_golden_model_1.ACC [2]);
  and (_10166_, \oc8051_golden_model_1.B [0], _10165_);
  nor (_10167_, _10166_, _10164_);
  nor (_10168_, _10167_, _10162_);
  not (_10169_, _10168_);
  nor (_10170_, _10158_, _10053_);
  nor (_10171_, _10170_, _10159_);
  and (_10172_, _10171_, _10169_);
  nor (_10173_, _10172_, _10159_);
  nor (_10174_, _10173_, _10154_);
  nor (_10175_, _10174_, _10153_);
  nor (_10176_, _10175_, _10145_);
  nor (_10177_, _10135_, \oc8051_golden_model_1.B [4]);
  nor (_10178_, _10177_, _10142_);
  not (_10179_, _10178_);
  nor (_10180_, _10179_, _10176_);
  not (_10181_, \oc8051_golden_model_1.B [5]);
  and (_10182_, _10098_, _10181_);
  and (_10183_, \oc8051_golden_model_1.B [4], _08506_);
  not (_10184_, _10183_);
  and (_10185_, _10184_, _10182_);
  not (_10186_, _10185_);
  nor (_10187_, _10186_, _10180_);
  nor (_10188_, _10187_, _10135_);
  nor (_10189_, _10188_, _10062_);
  not (_10190_, \oc8051_golden_model_1.B [4]);
  and (_10191_, _10175_, _10145_);
  nor (_10192_, _10191_, _10176_);
  not (_10193_, _10192_);
  and (_10194_, _10193_, _10187_);
  nor (_10195_, _10187_, _10141_);
  nor (_10196_, _10195_, _10194_);
  and (_10197_, _10196_, _10190_);
  nor (_10198_, _10196_, _10190_);
  nor (_10199_, _10198_, _10197_);
  not (_10200_, _10199_);
  nor (_10201_, _10187_, _10152_);
  nor (_10202_, _10154_, _10153_);
  and (_10203_, _10202_, _10173_);
  nor (_10204_, _10202_, _10173_);
  nor (_10205_, _10204_, _10203_);
  not (_10206_, _10205_);
  and (_10207_, _10206_, _10187_);
  nor (_10208_, _10207_, _10201_);
  nor (_10209_, _10208_, \oc8051_golden_model_1.B [3]);
  and (_10210_, _10208_, \oc8051_golden_model_1.B [3]);
  nor (_10211_, _10171_, _10169_);
  nor (_10212_, _10211_, _10172_);
  not (_10213_, _10212_);
  and (_10214_, _10213_, _10187_);
  nor (_10215_, _10187_, _10158_);
  nor (_10216_, _10215_, _10214_);
  and (_10217_, _10216_, _10111_);
  not (_10218_, \oc8051_golden_model_1.ACC [3]);
  nor (_10219_, _10187_, _10218_);
  and (_10220_, _10187_, _10161_);
  or (_10221_, _10220_, _10219_);
  and (_10222_, _10221_, _10053_);
  nor (_10223_, _10221_, _10053_);
  nor (_10224_, _10223_, _10166_);
  nor (_10225_, _10224_, _10222_);
  nor (_10226_, _10216_, _10111_);
  nor (_10227_, _10226_, _10217_);
  not (_10228_, _10227_);
  nor (_10229_, _10228_, _10225_);
  nor (_10230_, _10229_, _10217_);
  nor (_10231_, _10230_, _10210_);
  nor (_10232_, _10231_, _10209_);
  nor (_10233_, _10232_, _10200_);
  nor (_10234_, _10189_, \oc8051_golden_model_1.B [5]);
  nor (_10235_, _10234_, _10197_);
  not (_10236_, _10235_);
  nor (_10237_, _10236_, _10233_);
  not (_10238_, _10237_);
  not (_10239_, _10098_);
  and (_10240_, \oc8051_golden_model_1.B [5], _08506_);
  nor (_10241_, _10240_, _10239_);
  and (_10242_, _10241_, _10238_);
  nor (_10243_, _10242_, _10189_);
  nor (_10244_, _10243_, _10062_);
  not (_10245_, _10242_);
  and (_10246_, _10232_, _10200_);
  nor (_10247_, _10246_, _10233_);
  nor (_10248_, _10247_, _10245_);
  nor (_10249_, _10242_, _10196_);
  nor (_10250_, _10249_, _10248_);
  and (_10251_, _10250_, _10181_);
  nor (_10252_, _10250_, _10181_);
  nor (_10253_, _10252_, _10251_);
  not (_10254_, _10253_);
  nor (_10255_, _10210_, _10209_);
  nor (_10256_, _10255_, _10230_);
  and (_10257_, _10255_, _10230_);
  or (_10258_, _10257_, _10256_);
  nor (_10259_, _10258_, _10245_);
  and (_10260_, _10245_, _10208_);
  nor (_10261_, _10260_, _10259_);
  and (_10262_, _10261_, _10190_);
  nor (_10263_, _10261_, _10190_);
  and (_10264_, _10228_, _10225_);
  nor (_10265_, _10264_, _10229_);
  nor (_10266_, _10265_, _10245_);
  nor (_10267_, _10242_, _10216_);
  nor (_10268_, _10267_, _10266_);
  and (_10269_, _10268_, _10097_);
  nor (_10270_, _10223_, _10222_);
  nor (_10271_, _10270_, _10166_);
  and (_10272_, _10270_, _10166_);
  or (_10273_, _10272_, _10271_);
  nor (_10274_, _10273_, _10245_);
  nor (_10275_, _10242_, _10221_);
  nor (_10276_, _10275_, _10274_);
  and (_10277_, _10276_, _10111_);
  nor (_10278_, _10276_, _10111_);
  nor (_10279_, _10166_, _10163_);
  and (_10280_, _10242_, _10279_);
  nor (_10281_, _10242_, \oc8051_golden_model_1.ACC [2]);
  nor (_10282_, _10281_, _10280_);
  and (_10283_, _10282_, _10053_);
  and (_10284_, _05937_, \oc8051_golden_model_1.B [0]);
  not (_10285_, _10284_);
  nor (_10286_, _10282_, _10053_);
  nor (_10287_, _10286_, _10283_);
  and (_10288_, _10287_, _10285_);
  nor (_10289_, _10288_, _10283_);
  nor (_10290_, _10289_, _10278_);
  nor (_10291_, _10290_, _10277_);
  not (_10292_, _10291_);
  nor (_10293_, _10268_, _10097_);
  nor (_10294_, _10293_, _10269_);
  and (_10295_, _10294_, _10292_);
  nor (_10296_, _10295_, _10269_);
  nor (_10297_, _10296_, _10263_);
  nor (_10298_, _10297_, _10262_);
  nor (_10299_, _10298_, _10254_);
  nor (_10300_, _10244_, \oc8051_golden_model_1.B [6]);
  or (_10301_, _10300_, _10251_);
  or (_10302_, _10301_, _10299_);
  and (_10303_, \oc8051_golden_model_1.B [6], _08506_);
  nor (_10304_, _10303_, \oc8051_golden_model_1.B [7]);
  and (_10305_, _10304_, _10302_);
  nor (_10306_, _10305_, _10244_);
  or (_10307_, _10306_, _10062_);
  nor (_10308_, _10307_, \oc8051_golden_model_1.B [7]);
  nor (_10309_, _10308_, _10014_);
  not (_10310_, \oc8051_golden_model_1.B [6]);
  and (_10311_, _10298_, _10254_);
  nor (_10312_, _10311_, _10299_);
  not (_10313_, _10312_);
  and (_10314_, _10313_, _10305_);
  nor (_10315_, _10305_, _10250_);
  nor (_10316_, _10315_, _10314_);
  nor (_10317_, _10316_, _10310_);
  not (_10318_, _10317_);
  nor (_10319_, _10318_, _10309_);
  nor (_10320_, _10278_, _10277_);
  or (_10321_, _10320_, _10289_);
  nand (_10322_, _10320_, _10289_);
  and (_10323_, _10322_, _10321_);
  and (_10324_, _10323_, _10305_);
  nor (_10325_, _10305_, _10276_);
  nor (_10326_, _10325_, _10324_);
  and (_10327_, _10326_, _10097_);
  nor (_10328_, _10326_, _10097_);
  nor (_10329_, _10328_, _10327_);
  nor (_10330_, _10287_, _10285_);
  nor (_10331_, _10330_, _10288_);
  and (_10332_, _10331_, _10305_);
  not (_10333_, _10282_);
  nor (_10334_, _10305_, _10333_);
  nor (_10335_, _10334_, _10332_);
  and (_10336_, _10335_, \oc8051_golden_model_1.B [2]);
  nor (_10337_, _10335_, \oc8051_golden_model_1.B [2]);
  nor (_10338_, _10337_, _10336_);
  and (_10339_, _10338_, _10329_);
  nor (_10340_, _10305_, \oc8051_golden_model_1.ACC [1]);
  nor (_10341_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  or (_10342_, _10341_, _09975_);
  and (_10343_, _10305_, _10342_);
  nor (_10344_, _10343_, _10340_);
  and (_10345_, _10344_, _10053_);
  nor (_10346_, _10344_, _10053_);
  and (_10347_, _10058_, \oc8051_golden_model_1.ACC [0]);
  not (_10348_, _10347_);
  nor (_10349_, _10348_, _10346_);
  nor (_10350_, _10349_, _10345_);
  and (_10351_, _10350_, _10339_);
  not (_10352_, _10351_);
  and (_10353_, _10336_, _10329_);
  nor (_10354_, _10353_, _10328_);
  and (_10355_, _10354_, _10352_);
  nor (_10356_, _10294_, _10292_);
  nor (_10357_, _10356_, _10295_);
  and (_10358_, _10357_, _10305_);
  not (_10359_, _10268_);
  nor (_10360_, _10305_, _10359_);
  nor (_10361_, _10360_, _10358_);
  and (_10362_, _10361_, \oc8051_golden_model_1.B [4]);
  nor (_10363_, _10361_, \oc8051_golden_model_1.B [4]);
  nor (_10364_, _10363_, _10362_);
  nor (_10365_, _10263_, _10262_);
  nor (_10366_, _10365_, _10296_);
  and (_10367_, _10365_, _10296_);
  nor (_10368_, _10367_, _10366_);
  and (_10369_, _10368_, _10305_);
  nor (_10370_, _10305_, _10261_);
  or (_10371_, _10370_, _10369_);
  and (_10372_, _10371_, \oc8051_golden_model_1.B [5]);
  nor (_10373_, _10371_, \oc8051_golden_model_1.B [5]);
  nor (_10374_, _10373_, _10372_);
  and (_10375_, _10374_, _10364_);
  and (_10376_, _10316_, _10310_);
  nor (_10377_, _10376_, _10317_);
  not (_10378_, _10377_);
  nor (_10379_, _10378_, _10309_);
  and (_10380_, _10379_, _10375_);
  not (_10381_, _10380_);
  nor (_10382_, _10381_, _10355_);
  and (_10383_, _10244_, \oc8051_golden_model_1.B [7]);
  and (_10384_, _10374_, _10362_);
  nor (_10385_, _10384_, _10372_);
  not (_10386_, _10385_);
  and (_10387_, _10386_, _10379_);
  or (_10388_, _10387_, _10383_);
  or (_10389_, _10388_, _10382_);
  nor (_10390_, _10389_, _10319_);
  nor (_10391_, _10346_, _10345_);
  and (_10392_, \oc8051_golden_model_1.B [0], _05997_);
  not (_10393_, _10392_);
  and (_10394_, _10393_, _10391_);
  and (_10395_, _10394_, _10348_);
  and (_10396_, _10395_, _10339_);
  and (_10397_, _10396_, _10380_);
  nor (_10398_, _10397_, _10390_);
  or (_10399_, _10398_, _10062_);
  and (_10400_, _10399_, _10307_);
  or (_10401_, _10400_, _10052_);
  and (_10402_, _10401_, _10051_);
  and (_10403_, _10402_, _07198_);
  and (_10404_, _08770_, _07911_);
  or (_10405_, _10404_, _09450_);
  and (_10406_, _10405_, _06371_);
  or (_10407_, _10406_, _06367_);
  or (_10408_, _10407_, _10403_);
  and (_10409_, _08988_, _07911_);
  or (_10410_, _10409_, _09450_);
  or (_10411_, _10410_, _07218_);
  and (_10412_, _10411_, _07216_);
  and (_10413_, _10412_, _10408_);
  or (_10414_, _10413_, _09453_);
  and (_10415_, _10414_, _07213_);
  or (_10416_, _09450_, _08007_);
  and (_10417_, _10405_, _06366_);
  and (_10418_, _10417_, _10416_);
  or (_10419_, _10418_, _10415_);
  and (_10420_, _10419_, _07210_);
  and (_10421_, _09463_, _06541_);
  and (_10422_, _10421_, _10416_);
  or (_10423_, _10422_, _06383_);
  or (_10424_, _10423_, _10420_);
  and (_10425_, _08985_, _07911_);
  or (_10426_, _09450_, _07231_);
  or (_10427_, _10426_, _10425_);
  and (_10428_, _10427_, _07229_);
  and (_10429_, _10428_, _10424_);
  nor (_10430_, _08508_, _09454_);
  or (_10431_, _10430_, _09450_);
  and (_10432_, _10431_, _06528_);
  or (_10433_, _10432_, _06563_);
  or (_10434_, _10433_, _10429_);
  or (_10435_, _09460_, _07241_);
  and (_10436_, _10435_, _06571_);
  and (_10437_, _10436_, _10434_);
  and (_10438_, _09483_, _06199_);
  or (_10439_, _10438_, _06188_);
  or (_10440_, _10439_, _10437_);
  and (_10441_, _08503_, _07911_);
  or (_10442_, _09450_, _06189_);
  or (_10443_, _10442_, _10441_);
  and (_10444_, _10443_, _01452_);
  and (_10445_, _10444_, _10440_);
  or (_10446_, _10445_, _09449_);
  and (_41178_, _10446_, _43223_);
  nor (_10447_, _01452_, _08506_);
  and (_10448_, _05934_, _06259_);
  nand (_10449_, _10448_, _10068_);
  and (_10450_, _06372_, _06259_);
  not (_10451_, _10450_);
  and (_10452_, _06256_, _06380_);
  and (_10453_, _07325_, \oc8051_golden_model_1.PSW [7]);
  and (_10454_, _10453_, _09381_);
  and (_10455_, _10454_, _09380_);
  and (_10456_, _10455_, _09379_);
  and (_10457_, _10456_, _09378_);
  and (_10458_, _10457_, _09377_);
  and (_10459_, _10458_, _09376_);
  nor (_10460_, _10459_, _08562_);
  and (_10461_, _10459_, _08562_);
  nor (_10462_, _10461_, _10460_);
  nor (_10463_, _10462_, _08506_);
  and (_10464_, _10462_, _08506_);
  nor (_10465_, _10464_, _10463_);
  nor (_10466_, _10458_, _09376_);
  nor (_10467_, _10466_, _10459_);
  and (_10468_, _10467_, \oc8051_golden_model_1.ACC [6]);
  nor (_10469_, _10467_, _10068_);
  and (_10470_, _10467_, _10068_);
  nor (_10471_, _10470_, _10469_);
  not (_10472_, _10471_);
  nor (_10473_, _10457_, _09377_);
  nor (_10474_, _10473_, _10458_);
  and (_10475_, _10474_, \oc8051_golden_model_1.ACC [5]);
  nor (_10476_, _10474_, _10122_);
  and (_10477_, _10474_, _10122_);
  nor (_10478_, _10477_, _10476_);
  nor (_10479_, _10456_, _09378_);
  nor (_10480_, _10479_, _10457_);
  nand (_10481_, _10480_, \oc8051_golden_model_1.ACC [4]);
  nor (_10482_, _10480_, _10087_);
  and (_10483_, _10480_, _10087_);
  or (_10484_, _10483_, _10482_);
  nor (_10485_, _10455_, _09379_);
  nor (_10486_, _10485_, _10456_);
  and (_10487_, _10486_, \oc8051_golden_model_1.ACC [3]);
  nor (_10488_, _10486_, _10218_);
  and (_10489_, _10486_, _10218_);
  nor (_10490_, _10489_, _10488_);
  nor (_10491_, _10454_, _09380_);
  nor (_10492_, _10491_, _10455_);
  and (_10493_, _10492_, \oc8051_golden_model_1.ACC [2]);
  nor (_10494_, _10492_, _10165_);
  and (_10495_, _10492_, _10165_);
  nor (_10496_, _10495_, _10494_);
  nor (_10497_, _10453_, _09381_);
  nor (_10498_, _10497_, _10454_);
  and (_10499_, _10498_, \oc8051_golden_model_1.ACC [1]);
  and (_10500_, _10498_, _05937_);
  nor (_10501_, _10498_, _05937_);
  nor (_10502_, _10501_, _10500_);
  not (_10503_, _10502_);
  nor (_10504_, _07325_, \oc8051_golden_model_1.PSW [7]);
  nor (_10505_, _10504_, _10453_);
  and (_10506_, _10505_, \oc8051_golden_model_1.ACC [0]);
  and (_10507_, _10506_, _10503_);
  nor (_10508_, _10507_, _10499_);
  nor (_10509_, _10508_, _10496_);
  nor (_10510_, _10509_, _10493_);
  nor (_10511_, _10510_, _10490_);
  or (_10512_, _10511_, _10487_);
  nand (_10513_, _10512_, _10484_);
  and (_10514_, _10513_, _10481_);
  nor (_10515_, _10514_, _10478_);
  or (_10516_, _10515_, _10475_);
  and (_10517_, _10516_, _10472_);
  nor (_10518_, _10517_, _10468_);
  nor (_10519_, _10518_, _10465_);
  and (_10520_, _10518_, _10465_);
  nor (_10521_, _10520_, _10519_);
  and (_10522_, _07129_, _06380_);
  not (_10523_, _07492_);
  and (_10524_, _10523_, _06359_);
  nor (_10525_, _10524_, _05915_);
  nor (_10526_, _10525_, _10522_);
  or (_10527_, _10526_, _10521_);
  nor (_10528_, _08004_, _08506_);
  not (_10529_, _10528_);
  nor (_10530_, _07129_, _06805_);
  nor (_10531_, _10530_, _05918_);
  nand (_10532_, _10531_, _10529_);
  and (_10533_, _06372_, _05888_);
  not (_10534_, _10533_);
  or (_10535_, _08509_, _06532_);
  and (_10536_, _10535_, _10534_);
  nor (_10537_, _07914_, _08506_);
  not (_10538_, _07914_);
  nor (_10539_, _08004_, _10538_);
  or (_10540_, _10539_, _10537_);
  or (_10541_, _10540_, _07188_);
  and (_10542_, _06372_, _05969_);
  not (_10543_, _10542_);
  and (_10544_, _08351_, \oc8051_golden_model_1.PSW [7]);
  and (_10545_, _10544_, _08302_);
  and (_10546_, _10545_, _08397_);
  and (_10547_, _10546_, _08257_);
  and (_10548_, _10547_, _08497_);
  and (_10549_, _10548_, _08212_);
  and (_10550_, _10549_, _08109_);
  nor (_10551_, _10550_, _08006_);
  and (_10552_, _10550_, _08006_);
  nor (_10553_, _10552_, _10551_);
  and (_10554_, _10553_, \oc8051_golden_model_1.ACC [7]);
  nor (_10555_, _10553_, \oc8051_golden_model_1.ACC [7]);
  nor (_10556_, _10555_, _10554_);
  not (_10557_, _10556_);
  nor (_10558_, _10549_, _08109_);
  nor (_10559_, _10558_, _10550_);
  nor (_10560_, _10559_, _10068_);
  nor (_10561_, _10548_, _08212_);
  nor (_10562_, _10561_, _10549_);
  and (_10563_, _10562_, _10122_);
  nor (_10564_, _10562_, _10122_);
  nor (_10565_, _10547_, _08497_);
  nor (_10566_, _10565_, _10548_);
  nor (_10567_, _10566_, _10087_);
  nor (_10568_, _10567_, _10564_);
  nor (_10569_, _10568_, _10563_);
  nor (_10570_, _10564_, _10563_);
  not (_10571_, _10570_);
  and (_10572_, _10566_, _10087_);
  or (_10573_, _10572_, _10567_);
  or (_10574_, _10573_, _10571_);
  nor (_10575_, _10546_, _08257_);
  nor (_10576_, _10575_, _10547_);
  nor (_10577_, _10576_, _10218_);
  and (_10578_, _10576_, _10218_);
  nor (_10579_, _10578_, _10577_);
  nor (_10580_, _10545_, _08397_);
  nor (_10581_, _10580_, _10546_);
  nor (_10582_, _10581_, _10165_);
  and (_10583_, _10581_, _10165_);
  nor (_10584_, _10583_, _10582_);
  and (_10585_, _10584_, _10579_);
  nor (_10586_, _10544_, _08302_);
  nor (_10587_, _10586_, _10545_);
  nor (_10588_, _10587_, _05937_);
  and (_10589_, _10587_, _05937_);
  nor (_10590_, _08351_, \oc8051_golden_model_1.PSW [7]);
  nor (_10591_, _10590_, _10544_);
  and (_10592_, _10591_, _05997_);
  nor (_10593_, _10592_, _10589_);
  or (_10594_, _10593_, _10588_);
  nand (_10595_, _10594_, _10585_);
  and (_10596_, _10582_, _10579_);
  nor (_10597_, _10596_, _10577_);
  and (_10598_, _10597_, _10595_);
  nor (_10599_, _10598_, _10574_);
  nor (_10600_, _10599_, _10569_);
  and (_10601_, _10559_, _10068_);
  nor (_10602_, _10560_, _10601_);
  not (_10603_, _10602_);
  nor (_10604_, _10603_, _10600_);
  or (_10605_, _10604_, _10560_);
  and (_10606_, _10605_, _10557_);
  nor (_10607_, _10605_, _10557_);
  or (_10608_, _10607_, _10606_);
  and (_10609_, _10608_, _06510_);
  and (_10610_, _06256_, _05969_);
  not (_10611_, _10610_);
  and (_10612_, _09399_, \oc8051_golden_model_1.PSW [7]);
  nor (_10613_, _10612_, _09022_);
  and (_10614_, _10612_, _09022_);
  nor (_10615_, _10614_, _10613_);
  and (_10616_, _10615_, \oc8051_golden_model_1.ACC [7]);
  nor (_10617_, _10615_, \oc8051_golden_model_1.ACC [7]);
  nor (_10618_, _10617_, _10616_);
  not (_10619_, _10618_);
  and (_10620_, _09398_, \oc8051_golden_model_1.PSW [7]);
  nor (_10621_, _10620_, _09067_);
  nor (_10622_, _10621_, _10612_);
  nor (_10623_, _10622_, _10068_);
  and (_10624_, _09397_, \oc8051_golden_model_1.PSW [7]);
  nor (_10625_, _10624_, _09113_);
  nor (_10626_, _10625_, _10620_);
  and (_10627_, _10626_, _10122_);
  nor (_10628_, _10626_, _10122_);
  and (_10629_, _09396_, \oc8051_golden_model_1.PSW [7]);
  nor (_10630_, _10629_, _09159_);
  nor (_10631_, _10630_, _10624_);
  nor (_10632_, _10631_, _10087_);
  nor (_10633_, _10632_, _10628_);
  nor (_10634_, _10633_, _10627_);
  nor (_10635_, _10628_, _10627_);
  not (_10636_, _10635_);
  and (_10637_, _10631_, _10087_);
  or (_10638_, _10637_, _10632_);
  or (_10639_, _10638_, _10636_);
  and (_10640_, _09395_, \oc8051_golden_model_1.PSW [7]);
  nor (_10641_, _10640_, _09205_);
  nor (_10642_, _10641_, _10629_);
  nor (_10643_, _10642_, _10218_);
  and (_10644_, _10642_, _10218_);
  nor (_10645_, _10644_, _10643_);
  and (_10646_, _09394_, \oc8051_golden_model_1.PSW [7]);
  nor (_10648_, _10646_, _09251_);
  nor (_10649_, _10648_, _10640_);
  nor (_10650_, _10649_, _10165_);
  and (_10651_, _10649_, _10165_);
  nor (_10652_, _10651_, _10650_);
  and (_10653_, _10652_, _10645_);
  and (_10654_, _09342_, \oc8051_golden_model_1.PSW [7]);
  nor (_10655_, _10654_, _09297_);
  nor (_10656_, _10655_, _10646_);
  nor (_10657_, _10656_, _05937_);
  and (_10659_, _10656_, _05937_);
  nor (_10660_, _09342_, \oc8051_golden_model_1.PSW [7]);
  nor (_10661_, _10660_, _10654_);
  and (_10662_, _10661_, _05997_);
  nor (_10663_, _10662_, _10659_);
  or (_10664_, _10663_, _10657_);
  nand (_10665_, _10664_, _10653_);
  and (_10666_, _10650_, _10645_);
  nor (_10667_, _10666_, _10643_);
  and (_10668_, _10667_, _10665_);
  nor (_10670_, _10668_, _10639_);
  nor (_10671_, _10670_, _10634_);
  and (_10672_, _10622_, _10068_);
  nor (_10673_, _10623_, _10672_);
  not (_10674_, _10673_);
  nor (_10675_, _10674_, _10671_);
  or (_10676_, _10675_, _10623_);
  and (_10677_, _10676_, _10619_);
  nor (_10678_, _10676_, _10619_);
  or (_10679_, _10678_, _10677_);
  or (_10681_, _10679_, _10611_);
  nor (_10682_, _05952_, _05965_);
  nand (_10683_, _10682_, _08004_);
  and (_10684_, _08685_, _07914_);
  or (_10685_, _10684_, _10537_);
  and (_10686_, _10685_, _06251_);
  and (_10687_, _06372_, _06471_);
  not (_10688_, _10687_);
  or (_10689_, _10688_, _08671_);
  and (_10690_, _06471_, _06817_);
  nor (_10692_, _07053_, _06357_);
  nor (_10693_, _10692_, _05954_);
  nor (_10694_, _10693_, _10690_);
  nor (_10695_, _06811_, _06472_);
  and (_10696_, _07455_, _06471_);
  not (_10697_, _10696_);
  and (_10698_, _10697_, _10695_);
  and (_10699_, _06471_, _06348_);
  and (_10700_, _06361_, _06471_);
  nor (_10701_, _10700_, _10699_);
  and (_10703_, _10701_, _10698_);
  and (_10704_, _10703_, _10694_);
  nor (_10705_, _10704_, _08004_);
  or (_10706_, _06808_, \oc8051_golden_model_1.ACC [7]);
  nand (_10707_, _06808_, \oc8051_golden_model_1.ACC [7]);
  and (_10708_, _10707_, _10706_);
  and (_10709_, _10708_, _10704_);
  or (_10710_, _10709_, _10687_);
  or (_10711_, _10710_, _10705_);
  not (_10712_, _05955_);
  nor (_10714_, _06251_, _10712_);
  and (_10715_, _10714_, _10711_);
  and (_10716_, _10715_, _10689_);
  or (_10717_, _10716_, _10686_);
  and (_10718_, _06372_, _06250_);
  not (_10719_, _10718_);
  and (_10720_, _10719_, _10717_);
  nor (_10721_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor (_10722_, _10721_, _10218_);
  and (_10723_, _10722_, \oc8051_golden_model_1.ACC [4]);
  and (_10724_, _10723_, \oc8051_golden_model_1.ACC [5]);
  and (_10725_, _10724_, \oc8051_golden_model_1.ACC [6]);
  and (_10726_, _10725_, \oc8051_golden_model_1.ACC [7]);
  nor (_10727_, _10725_, \oc8051_golden_model_1.ACC [7]);
  nor (_10728_, _10727_, _10726_);
  nor (_10729_, _10723_, \oc8051_golden_model_1.ACC [5]);
  nor (_10730_, _10729_, _10724_);
  nor (_10731_, _10724_, \oc8051_golden_model_1.ACC [6]);
  nor (_10732_, _10731_, _10725_);
  nor (_10733_, _10732_, _10730_);
  not (_10734_, _10733_);
  and (_10735_, _10734_, _10728_);
  not (_10736_, _10735_);
  nor (_10737_, _10726_, \oc8051_golden_model_1.PSW [7]);
  and (_10738_, _10737_, _10736_);
  nor (_10739_, _10738_, _10733_);
  or (_10740_, _10739_, _10728_);
  and (_10741_, _10736_, _10718_);
  and (_10742_, _10741_, _10740_);
  or (_10743_, _10742_, _06475_);
  or (_10744_, _10743_, _10720_);
  nor (_10745_, _08545_, _08506_);
  and (_10746_, _08560_, _08545_);
  or (_10747_, _10746_, _10745_);
  or (_10748_, _10747_, _06476_);
  and (_10749_, _10748_, _07142_);
  and (_10750_, _10749_, _10744_);
  and (_10751_, _10540_, _06468_);
  or (_10752_, _10751_, _10682_);
  or (_10753_, _10752_, _10750_);
  and (_10754_, _10753_, _10683_);
  or (_10755_, _10754_, _07153_);
  or (_10756_, _08671_, _07353_);
  and (_10757_, _10756_, _06801_);
  and (_10758_, _10757_, _10755_);
  and (_10759_, _06372_, _06246_);
  nor (_10760_, _08006_, _06801_);
  or (_10761_, _10760_, _10759_);
  or (_10762_, _10761_, _10758_);
  nand (_10763_, _10759_, _10218_);
  and (_10764_, _10763_, _10762_);
  or (_10765_, _10764_, _06483_);
  and (_10766_, _08698_, _08545_);
  or (_10767_, _10766_, _10745_);
  or (_10768_, _10767_, _06484_);
  and (_10769_, _10768_, _07164_);
  and (_10770_, _10769_, _10765_);
  or (_10771_, _10745_, _08706_);
  and (_10772_, _10771_, _06461_);
  and (_10773_, _10772_, _10747_);
  or (_10774_, _10773_, _09487_);
  or (_10775_, _10774_, _10770_);
  nor (_10776_, _09994_, _09992_);
  nor (_10777_, _10776_, _09995_);
  or (_10778_, _10777_, _09494_);
  nand (_10779_, _05969_, _05657_);
  and (_10780_, _10779_, _10778_);
  and (_10781_, _10780_, _10775_);
  not (_10782_, _10465_);
  nor (_10783_, _10482_, _10476_);
  nor (_10784_, _10783_, _10477_);
  not (_10785_, _10478_);
  or (_10786_, _10484_, _10785_);
  and (_10787_, _10496_, _10490_);
  and (_10788_, _10505_, _05997_);
  nor (_10789_, _10788_, _10500_);
  or (_10790_, _10789_, _10501_);
  nand (_10791_, _10790_, _10787_);
  and (_10792_, _10494_, _10490_);
  nor (_10793_, _10792_, _10488_);
  and (_10794_, _10793_, _10791_);
  nor (_10795_, _10794_, _10786_);
  nor (_10796_, _10795_, _10784_);
  nor (_10797_, _10796_, _10472_);
  or (_10798_, _10797_, _10469_);
  and (_10799_, _10798_, _10782_);
  nor (_10800_, _10798_, _10782_);
  nor (_10801_, _10800_, _10799_);
  nor (_10802_, _10801_, _10779_);
  or (_10803_, _10802_, _10610_);
  or (_10804_, _10803_, _10781_);
  and (_10805_, _10804_, _06516_);
  and (_10806_, _10805_, _10681_);
  or (_10807_, _10806_, _10609_);
  and (_10808_, _10807_, _10543_);
  and (_10809_, _07921_, \oc8051_golden_model_1.PSW [7]);
  and (_10810_, _10809_, _07877_);
  and (_10811_, _10810_, _07869_);
  and (_10812_, _10811_, _07742_);
  nor (_10813_, _10812_, _07904_);
  and (_10814_, _10812_, _07904_);
  nor (_10815_, _10814_, _10813_);
  and (_10816_, _10815_, \oc8051_golden_model_1.ACC [7]);
  nor (_10817_, _10815_, \oc8051_golden_model_1.ACC [7]);
  nor (_10818_, _10817_, _10816_);
  not (_10819_, _10818_);
  nor (_10820_, _10811_, _07742_);
  nor (_10821_, _10820_, _10812_);
  nor (_10822_, _10821_, _10068_);
  and (_10823_, _10810_, _06244_);
  nor (_10824_, _10823_, _07862_);
  nor (_10825_, _10824_, _10811_);
  and (_10826_, _10825_, _10122_);
  nor (_10827_, _10825_, _10122_);
  nor (_10828_, _10810_, _06244_);
  nor (_10829_, _10828_, _10823_);
  nor (_10830_, _10829_, _10087_);
  nor (_10831_, _10830_, _10827_);
  nor (_10832_, _10831_, _10826_);
  nor (_10833_, _10827_, _10826_);
  not (_10834_, _10833_);
  and (_10835_, _10829_, _10087_);
  or (_10836_, _10835_, _10830_);
  or (_10837_, _10836_, _10834_);
  nor (_10838_, _08725_, _06328_);
  nor (_10839_, _10838_, _10810_);
  and (_10840_, _10839_, _10218_);
  nor (_10841_, _10839_, _10218_);
  nor (_10842_, _10841_, _10840_);
  nor (_10843_, _10809_, _06751_);
  nor (_10844_, _10843_, _08725_);
  and (_10845_, _10844_, _10165_);
  nor (_10846_, _10844_, _10165_);
  nor (_10847_, _10846_, _10845_);
  and (_10848_, _10847_, _10842_);
  and (_10849_, _06799_, \oc8051_golden_model_1.PSW [7]);
  nor (_10850_, _10849_, _06156_);
  nor (_10851_, _10850_, _10809_);
  and (_10852_, _10851_, _05937_);
  nor (_10853_, _10851_, _05937_);
  not (_10854_, \oc8051_golden_model_1.PSW [7]);
  and (_10855_, _06799_, _10854_);
  and (_10856_, _06802_, \oc8051_golden_model_1.PSW [7]);
  nor (_10857_, _10856_, _10855_);
  or (_10858_, _10857_, \oc8051_golden_model_1.ACC [0]);
  nor (_10859_, _10858_, _10853_);
  nor (_10860_, _10859_, _10852_);
  nand (_10861_, _10860_, _10848_);
  and (_10862_, _10846_, _10842_);
  nor (_10863_, _10862_, _10841_);
  and (_10864_, _10863_, _10861_);
  nor (_10865_, _10864_, _10837_);
  nor (_10866_, _10865_, _10832_);
  and (_10867_, _10821_, _10068_);
  nor (_10868_, _10822_, _10867_);
  not (_10869_, _10868_);
  nor (_10870_, _10869_, _10866_);
  or (_10871_, _10870_, _10822_);
  and (_10872_, _10871_, _10819_);
  nor (_10873_, _10871_, _10819_);
  or (_10874_, _10873_, _10872_);
  and (_10875_, _10874_, _10542_);
  or (_10876_, _10875_, _10808_);
  and (_10877_, _10876_, _05977_);
  and (_10878_, _06187_, _05976_);
  or (_10879_, _10878_, _10877_);
  and (_10880_, _10879_, _06242_);
  and (_10881_, _08726_, _08545_);
  or (_10882_, _10881_, _10745_);
  and (_10883_, _10882_, _06241_);
  or (_10884_, _10883_, _07187_);
  or (_10885_, _10884_, _10880_);
  and (_10886_, _10885_, _10541_);
  or (_10887_, _10886_, _07182_);
  and (_10888_, _08671_, _07914_);
  or (_10889_, _10537_, _07183_);
  or (_10890_, _10889_, _10888_);
  and (_10891_, _10890_, _06336_);
  and (_10892_, _10891_, _10887_);
  and (_10893_, _08966_, _07914_);
  or (_10894_, _10893_, _10537_);
  and (_10895_, _10894_, _05968_);
  or (_10896_, _10895_, _10046_);
  or (_10897_, _10896_, _10892_);
  or (_10898_, _10066_, _10052_);
  and (_10899_, _10898_, _05975_);
  and (_10900_, _10899_, _10897_);
  and (_10901_, _06187_, _05935_);
  or (_10902_, _10901_, _06371_);
  or (_10903_, _10902_, _10900_);
  and (_10904_, _06372_, _05894_);
  not (_10905_, _10904_);
  and (_10906_, _08770_, _07914_);
  or (_10907_, _10906_, _10537_);
  or (_10908_, _10907_, _07198_);
  and (_10909_, _10908_, _10905_);
  and (_10910_, _10909_, _10903_);
  and (_10911_, _10904_, _06187_);
  and (_10912_, _07492_, _05888_);
  or (_10913_, _10912_, _10911_);
  or (_10914_, _10913_, _10910_);
  and (_10915_, _08004_, _08506_);
  nor (_10916_, _10915_, _10528_);
  not (_10917_, _10912_);
  or (_10918_, _10917_, _10916_);
  nor (_10919_, _06359_, _06924_);
  not (_10920_, _10919_);
  and (_10921_, _10920_, _10918_);
  and (_10922_, _10921_, _10914_);
  and (_10923_, _10919_, _10916_);
  and (_10924_, _07129_, _05888_);
  or (_10925_, _10924_, _10923_);
  or (_10926_, _10925_, _10922_);
  not (_10927_, _10924_);
  or (_10928_, _10927_, _10916_);
  and (_10929_, _06256_, _05888_);
  not (_10930_, _10929_);
  and (_10931_, _10930_, _10928_);
  and (_10932_, _10931_, _10926_);
  nor (_10933_, _08671_, \oc8051_golden_model_1.ACC [7]);
  and (_10934_, _08671_, \oc8051_golden_model_1.ACC [7]);
  nor (_10935_, _10934_, _10933_);
  and (_10936_, _10929_, _10935_);
  or (_10937_, _10936_, _06531_);
  or (_10938_, _10937_, _10932_);
  and (_10939_, _10938_, _10536_);
  nor (_10940_, _06187_, \oc8051_golden_model_1.ACC [7]);
  and (_10941_, _06187_, \oc8051_golden_model_1.ACC [7]);
  nor (_10942_, _10941_, _10940_);
  and (_10943_, _10942_, _10533_);
  or (_10944_, _10943_, _06367_);
  or (_10945_, _10944_, _10939_);
  and (_10946_, _08988_, _07914_);
  or (_10947_, _10946_, _10537_);
  or (_10948_, _10947_, _07218_);
  and (_10949_, _10948_, _10945_);
  or (_10950_, _10949_, _06533_);
  nor (_10951_, _10537_, _07216_);
  nand (_10952_, _10523_, _10692_);
  and (_10953_, _10952_, _06365_);
  nor (_10954_, _10953_, _10951_);
  and (_10955_, _10954_, _10950_);
  and (_10956_, _10953_, _10528_);
  or (_10957_, _10956_, _10531_);
  or (_10958_, _10957_, _10955_);
  and (_10959_, _10958_, _10532_);
  and (_10960_, _06256_, _06365_);
  or (_10961_, _10960_, _10959_);
  not (_10962_, _10960_);
  or (_10963_, _10962_, _10934_);
  and (_10964_, _10963_, _06540_);
  and (_10965_, _10964_, _10961_);
  and (_10966_, _06372_, _06365_);
  nor (_10967_, _10966_, _06539_);
  not (_10968_, _10967_);
  or (_10969_, _10966_, _08507_);
  and (_10970_, _10969_, _10968_);
  or (_10971_, _10970_, _10965_);
  not (_10972_, _10966_);
  or (_10973_, _10972_, _10941_);
  and (_10974_, _10973_, _07213_);
  and (_10975_, _10974_, _10971_);
  nand (_10976_, _10907_, _06366_);
  nor (_10977_, _10976_, _08508_);
  or (_10978_, _10977_, _07032_);
  or (_10979_, _10978_, _10975_);
  and (_10980_, _06194_, _06382_);
  and (_10981_, _07053_, _06382_);
  nor (_10982_, _10981_, _10980_);
  nand (_10983_, _10915_, _07032_);
  and (_10984_, _10983_, _10982_);
  and (_10985_, _10984_, _10979_);
  and (_10986_, _06382_, _06817_);
  and (_10987_, _06361_, _06382_);
  or (_10988_, _10987_, _10986_);
  nor (_10989_, _10982_, _10915_);
  or (_10990_, _10989_, _10988_);
  or (_10991_, _10990_, _10985_);
  and (_10992_, _06382_, _06348_);
  not (_10993_, _10992_);
  nand (_10994_, _10988_, _10915_);
  and (_10995_, _10994_, _10993_);
  and (_10996_, _10995_, _10991_);
  nor (_10997_, _10915_, _10993_);
  and (_10998_, _06256_, _06382_);
  or (_10999_, _10998_, _10997_);
  or (_11000_, _10999_, _10996_);
  nand (_11001_, _10998_, _10933_);
  and (_11002_, _11001_, _06527_);
  and (_11003_, _11002_, _11000_);
  and (_11004_, _06372_, _06382_);
  nor (_11005_, _11004_, _06526_);
  not (_11006_, _11005_);
  not (_11007_, _11004_);
  nand (_11008_, _11007_, _08508_);
  and (_11009_, _11008_, _11006_);
  or (_11010_, _11009_, _11003_);
  nand (_11011_, _11004_, _10940_);
  and (_11012_, _11011_, _07231_);
  and (_11013_, _11012_, _11010_);
  not (_11014_, _10526_);
  and (_11015_, _08985_, _07914_);
  or (_11016_, _11015_, _10537_);
  and (_11017_, _11016_, _06383_);
  or (_11018_, _11017_, _11014_);
  or (_11019_, _11018_, _11013_);
  and (_11020_, _11019_, _10527_);
  or (_11021_, _11020_, _10452_);
  not (_11022_, _10452_);
  nand (_11023_, _10622_, \oc8051_golden_model_1.ACC [6]);
  and (_11024_, _10626_, \oc8051_golden_model_1.ACC [5]);
  nand (_11025_, _10631_, \oc8051_golden_model_1.ACC [4]);
  and (_11026_, _10642_, \oc8051_golden_model_1.ACC [3]);
  and (_11027_, _10649_, \oc8051_golden_model_1.ACC [2]);
  and (_11028_, _10656_, \oc8051_golden_model_1.ACC [1]);
  nor (_11029_, _10659_, _10657_);
  not (_11030_, _11029_);
  and (_11031_, _10661_, \oc8051_golden_model_1.ACC [0]);
  and (_11032_, _11031_, _11030_);
  nor (_11033_, _11032_, _11028_);
  nor (_11034_, _11033_, _10652_);
  nor (_11035_, _11034_, _11027_);
  nor (_11036_, _11035_, _10645_);
  or (_11037_, _11036_, _11026_);
  nand (_11038_, _11037_, _10638_);
  and (_11039_, _11038_, _11025_);
  nor (_11040_, _11039_, _10635_);
  or (_11041_, _11040_, _11024_);
  nand (_11042_, _11041_, _10674_);
  and (_11043_, _11042_, _11023_);
  nor (_11044_, _11043_, _10618_);
  and (_11045_, _11043_, _10618_);
  nor (_11046_, _11045_, _11044_);
  or (_11047_, _11046_, _11022_);
  and (_11048_, _11047_, _06538_);
  and (_11049_, _11048_, _11021_);
  and (_11050_, _06372_, _06380_);
  nor (_11051_, _11050_, _06537_);
  not (_11052_, _11051_);
  and (_11053_, _10559_, \oc8051_golden_model_1.ACC [6]);
  and (_11054_, _10562_, \oc8051_golden_model_1.ACC [5]);
  nand (_11055_, _10566_, \oc8051_golden_model_1.ACC [4]);
  and (_11056_, _10576_, \oc8051_golden_model_1.ACC [3]);
  and (_11057_, _10581_, \oc8051_golden_model_1.ACC [2]);
  and (_11058_, _10587_, \oc8051_golden_model_1.ACC [1]);
  nor (_11059_, _10589_, _10588_);
  not (_11060_, _11059_);
  and (_11061_, _10591_, \oc8051_golden_model_1.ACC [0]);
  and (_11062_, _11061_, _11060_);
  nor (_11063_, _11062_, _11058_);
  nor (_11064_, _11063_, _10584_);
  nor (_11065_, _11064_, _11057_);
  nor (_11066_, _11065_, _10579_);
  or (_11067_, _11066_, _11056_);
  nand (_11068_, _11067_, _10573_);
  and (_11069_, _11068_, _11055_);
  nor (_11070_, _11069_, _10570_);
  or (_11071_, _11070_, _11054_);
  and (_11072_, _11071_, _10603_);
  nor (_11073_, _11072_, _11053_);
  nor (_11074_, _11073_, _10556_);
  and (_11075_, _11073_, _10556_);
  nor (_11076_, _11075_, _11074_);
  or (_11077_, _11076_, _11050_);
  and (_11078_, _11077_, _11052_);
  or (_11079_, _11078_, _11049_);
  and (_11080_, _05934_, _06380_);
  not (_11081_, _11080_);
  not (_11082_, _11050_);
  nand (_11083_, _10821_, \oc8051_golden_model_1.ACC [6]);
  and (_11084_, _10825_, \oc8051_golden_model_1.ACC [5]);
  nand (_11085_, _10829_, \oc8051_golden_model_1.ACC [4]);
  and (_11086_, _10839_, \oc8051_golden_model_1.ACC [3]);
  and (_11087_, _10844_, \oc8051_golden_model_1.ACC [2]);
  and (_11088_, _10851_, \oc8051_golden_model_1.ACC [1]);
  nor (_11089_, _10853_, _10852_);
  not (_11090_, _11089_);
  nor (_11091_, _10857_, _05997_);
  and (_11092_, _11091_, _11090_);
  nor (_11093_, _11092_, _11088_);
  nor (_11094_, _11093_, _10847_);
  nor (_11095_, _11094_, _11087_);
  nor (_11096_, _11095_, _10842_);
  or (_11097_, _11096_, _11086_);
  nand (_11098_, _11097_, _10836_);
  and (_11099_, _11098_, _11085_);
  nor (_11100_, _11099_, _10833_);
  or (_11101_, _11100_, _11084_);
  nand (_11102_, _11101_, _10869_);
  and (_11103_, _11102_, _11083_);
  nor (_11104_, _11103_, _10818_);
  and (_11105_, _11103_, _10818_);
  nor (_11106_, _11105_, _11104_);
  or (_11107_, _11106_, _11082_);
  and (_11108_, _11107_, _11081_);
  and (_11109_, _11108_, _11079_);
  and (_11110_, _11080_, \oc8051_golden_model_1.ACC [6]);
  nor (_11111_, _10524_, _05923_);
  or (_11112_, _11111_, _11110_);
  or (_11113_, _11112_, _11109_);
  and (_11114_, _07129_, _06259_);
  not (_11115_, _11114_);
  not (_11116_, _11111_);
  nor (_11117_, _08106_, _10068_);
  and (_11118_, _08106_, _10068_);
  nor (_11119_, _11117_, _11118_);
  nor (_11120_, _08209_, _10122_);
  and (_11121_, _08209_, _10122_);
  nor (_11122_, _11121_, _11120_);
  nor (_11123_, _08494_, _10087_);
  nand (_11124_, _08494_, _10087_);
  not (_11125_, _11123_);
  and (_11126_, _11125_, _11124_);
  nor (_11127_, _07713_, _10218_);
  and (_11128_, _07713_, _10218_);
  nor (_11129_, _07578_, _10165_);
  and (_11130_, _07578_, _10165_);
  nor (_11131_, _11129_, _11130_);
  nor (_11132_, _07120_, _05937_);
  and (_11133_, _07120_, _05937_);
  nor (_11134_, _11132_, _11133_);
  and (_11135_, _07325_, \oc8051_golden_model_1.ACC [0]);
  and (_11136_, _11135_, _11134_);
  nor (_11137_, _11136_, _11132_);
  not (_11138_, _11137_);
  and (_11139_, _11138_, _11131_);
  nor (_11140_, _11139_, _11129_);
  nor (_11141_, _11140_, _11128_);
  or (_11142_, _11141_, _11127_);
  and (_11143_, _11142_, _11126_);
  nor (_11144_, _11143_, _11123_);
  not (_11145_, _11144_);
  and (_11146_, _11145_, _11122_);
  or (_11147_, _11146_, _11120_);
  and (_11148_, _11147_, _11119_);
  nor (_11149_, _11148_, _11117_);
  nor (_11150_, _11149_, _10916_);
  and (_11151_, _11149_, _10916_);
  or (_11152_, _11151_, _11150_);
  or (_11153_, _11152_, _11116_);
  and (_11154_, _11153_, _11115_);
  and (_11155_, _11154_, _11113_);
  and (_11156_, _06256_, _06259_);
  and (_11157_, _11152_, _11114_);
  or (_11158_, _11157_, _11156_);
  or (_11159_, _11158_, _11155_);
  not (_11160_, _11156_);
  and (_11161_, _09067_, \oc8051_golden_model_1.ACC [6]);
  nor (_11162_, _09067_, \oc8051_golden_model_1.ACC [6]);
  nor (_11163_, _11162_, _11161_);
  and (_11164_, _09113_, \oc8051_golden_model_1.ACC [5]);
  nor (_11165_, _09113_, \oc8051_golden_model_1.ACC [5]);
  or (_11166_, _11165_, _11164_);
  and (_11167_, _09159_, \oc8051_golden_model_1.ACC [4]);
  not (_11168_, _11167_);
  or (_11169_, _09159_, \oc8051_golden_model_1.ACC [4]);
  and (_11170_, _11169_, _11168_);
  and (_11171_, _09205_, \oc8051_golden_model_1.ACC [3]);
  nor (_11172_, _09205_, \oc8051_golden_model_1.ACC [3]);
  and (_11173_, _09251_, \oc8051_golden_model_1.ACC [2]);
  nor (_11174_, _09251_, \oc8051_golden_model_1.ACC [2]);
  nor (_11175_, _11174_, _11173_);
  and (_11176_, _09297_, \oc8051_golden_model_1.ACC [1]);
  nor (_11177_, _09297_, \oc8051_golden_model_1.ACC [1]);
  nor (_11178_, _11177_, _11176_);
  and (_11179_, _09342_, \oc8051_golden_model_1.ACC [0]);
  and (_11180_, _11179_, _11178_);
  nor (_11181_, _11180_, _11176_);
  not (_11182_, _11181_);
  and (_11183_, _11182_, _11175_);
  nor (_11184_, _11183_, _11173_);
  nor (_11185_, _11184_, _11172_);
  or (_11186_, _11185_, _11171_);
  nand (_11187_, _11186_, _11170_);
  and (_11188_, _11187_, _11168_);
  nor (_11189_, _11188_, _11166_);
  or (_11190_, _11189_, _11164_);
  and (_11191_, _11190_, _11163_);
  nor (_11192_, _11191_, _11161_);
  and (_11193_, _11192_, _10935_);
  nor (_11194_, _11192_, _10935_);
  or (_11195_, _11194_, _11193_);
  or (_11196_, _11195_, _11160_);
  and (_11197_, _11196_, _06295_);
  and (_11198_, _11197_, _11159_);
  nor (_11199_, _08108_, _10068_);
  not (_11200_, _11199_);
  and (_11201_, _08108_, _10068_);
  nor (_11202_, _11201_, _11199_);
  nor (_11203_, _08211_, _10122_);
  and (_11204_, _08211_, _10122_);
  nor (_11205_, _11204_, _11203_);
  nor (_11206_, _08496_, _10087_);
  not (_11207_, _11206_);
  and (_11208_, _08496_, _10087_);
  nor (_11209_, _11208_, _11206_);
  nor (_11210_, _08256_, _10218_);
  and (_11211_, _08256_, _10218_);
  nor (_11212_, _08396_, _10165_);
  and (_11213_, _08396_, _10165_);
  nor (_11214_, _11213_, _11212_);
  nor (_11215_, _08301_, _05937_);
  and (_11216_, _08301_, _05937_);
  nor (_11217_, _11216_, _11215_);
  and (_11218_, _08351_, \oc8051_golden_model_1.ACC [0]);
  and (_11219_, _11218_, _11217_);
  nor (_11220_, _11219_, _11215_);
  not (_11221_, _11220_);
  and (_11222_, _11221_, _11214_);
  nor (_11223_, _11222_, _11212_);
  nor (_11224_, _11223_, _11211_);
  or (_11225_, _11224_, _11210_);
  nand (_11226_, _11225_, _11209_);
  and (_11227_, _11226_, _11207_);
  not (_11228_, _11227_);
  and (_11229_, _11228_, _11205_);
  or (_11230_, _11229_, _11203_);
  nand (_11231_, _11230_, _11202_);
  and (_11232_, _11231_, _11200_);
  nor (_11233_, _11232_, _08509_);
  and (_11234_, _11232_, _08509_);
  or (_11235_, _11234_, _11233_);
  and (_11236_, _11235_, _06293_);
  or (_11237_, _11236_, _11198_);
  and (_11238_, _11237_, _10451_);
  nor (_11239_, _06326_, _10068_);
  and (_11240_, _06326_, _10068_);
  nor (_11241_, _11239_, _11240_);
  nand (_11242_, _06608_, _10122_);
  nor (_11243_, _06608_, _10122_);
  nor (_11244_, _06230_, _10087_);
  not (_11245_, _11244_);
  and (_11246_, _06230_, _10087_);
  nor (_11247_, _11244_, _11246_);
  nor (_11248_, _06292_, _10218_);
  and (_11249_, _06292_, _10218_);
  nor (_11250_, _06750_, _10165_);
  and (_11251_, _06750_, _10165_);
  nor (_11252_, _11250_, _11251_);
  nor (_11253_, _06155_, _05937_);
  and (_11254_, _06155_, _05937_);
  nor (_11255_, _11253_, _11254_);
  and (_11256_, _06799_, \oc8051_golden_model_1.ACC [0]);
  and (_11257_, _11256_, _11255_);
  nor (_11258_, _11257_, _11253_);
  not (_11259_, _11258_);
  and (_11260_, _11259_, _11252_);
  nor (_11261_, _11260_, _11250_);
  nor (_11262_, _11261_, _11249_);
  or (_11263_, _11262_, _11248_);
  nand (_11264_, _11263_, _11247_);
  and (_11265_, _11264_, _11245_);
  not (_11266_, _11265_);
  or (_11267_, _11266_, _11243_);
  and (_11268_, _11267_, _11242_);
  and (_11269_, _11268_, _11241_);
  nor (_11270_, _11269_, _11239_);
  nor (_11271_, _11270_, _10942_);
  and (_11272_, _11270_, _10942_);
  or (_11273_, _11272_, _11271_);
  and (_11274_, _11273_, _10450_);
  or (_11275_, _11274_, _10448_);
  or (_11276_, _11275_, _11238_);
  and (_11277_, _11276_, _10449_);
  or (_11278_, _11277_, _06563_);
  and (_11279_, _06372_, _05911_);
  not (_11280_, _11279_);
  or (_11281_, _10685_, _07241_);
  and (_11282_, _11281_, _11280_);
  and (_11283_, _11282_, _11278_);
  and (_11284_, _05934_, _05911_);
  and (_11285_, _10721_, _05997_);
  and (_11286_, _11285_, _10218_);
  and (_11287_, _11286_, _10087_);
  and (_11288_, _11287_, _10122_);
  and (_11289_, _11288_, _10068_);
  nor (_11290_, _11289_, _08506_);
  and (_11291_, _11289_, _08506_);
  or (_11292_, _11291_, _11290_);
  and (_11293_, _11292_, _11279_);
  or (_11294_, _11293_, _11284_);
  or (_11295_, _11294_, _11283_);
  nand (_11296_, _11284_, _10854_);
  and (_11297_, _11296_, _06571_);
  and (_11298_, _11297_, _11295_);
  and (_11299_, _10767_, _06199_);
  or (_11300_, _11299_, _06188_);
  or (_11301_, _11300_, _11298_);
  and (_11302_, _06372_, _05906_);
  not (_11303_, _11302_);
  and (_11304_, _08503_, _07914_);
  or (_11305_, _11304_, _10537_);
  or (_11306_, _11305_, _06189_);
  and (_11307_, _11306_, _11303_);
  and (_11308_, _11307_, _11301_);
  and (_11309_, _05934_, _05906_);
  and (_11310_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and (_11311_, _11310_, \oc8051_golden_model_1.ACC [2]);
  and (_11312_, _11311_, \oc8051_golden_model_1.ACC [3]);
  and (_11313_, _11312_, \oc8051_golden_model_1.ACC [4]);
  and (_11314_, _11313_, \oc8051_golden_model_1.ACC [5]);
  and (_11315_, _11314_, \oc8051_golden_model_1.ACC [6]);
  nor (_11316_, _11315_, _08506_);
  and (_11317_, _11315_, _08506_);
  or (_11318_, _11317_, _11316_);
  and (_11319_, _11318_, _11302_);
  or (_11320_, _11319_, _11309_);
  or (_11321_, _11320_, _11308_);
  nand (_11322_, _11309_, _05997_);
  and (_11323_, _11322_, _01452_);
  and (_11324_, _11323_, _11321_);
  or (_11325_, _11324_, _10447_);
  and (_41179_, _11325_, _43223_);
  not (_11326_, _07923_);
  and (_11327_, _11326_, \oc8051_golden_model_1.PCON [7]);
  and (_11328_, _08509_, _07923_);
  or (_11329_, _11328_, _11327_);
  and (_11330_, _11329_, _06533_);
  nor (_11331_, _08004_, _11326_);
  or (_11332_, _11331_, _11327_);
  or (_11333_, _11332_, _07188_);
  and (_11334_, _08685_, _07923_);
  or (_11335_, _11334_, _11327_);
  or (_11336_, _11335_, _06252_);
  and (_11337_, _07923_, \oc8051_golden_model_1.ACC [7]);
  or (_11338_, _11337_, _11327_);
  and (_11339_, _11338_, _07123_);
  and (_11340_, _07124_, \oc8051_golden_model_1.PCON [7]);
  or (_11341_, _11340_, _06251_);
  or (_11342_, _11341_, _11339_);
  and (_11343_, _11342_, _07142_);
  and (_11344_, _11343_, _11336_);
  and (_11345_, _11332_, _06468_);
  or (_11346_, _11345_, _11344_);
  and (_11347_, _11346_, _06801_);
  and (_11348_, _11338_, _06466_);
  or (_11349_, _11348_, _07187_);
  or (_11350_, _11349_, _11347_);
  and (_11351_, _11350_, _11333_);
  or (_11352_, _11351_, _07182_);
  and (_11353_, _08671_, _07923_);
  or (_11354_, _11327_, _07183_);
  or (_11355_, _11354_, _11353_);
  and (_11356_, _11355_, _06336_);
  and (_11357_, _11356_, _11352_);
  and (_11358_, _08966_, _07923_);
  or (_11359_, _11358_, _11327_);
  and (_11360_, _11359_, _05968_);
  or (_11361_, _11360_, _06371_);
  or (_11362_, _11361_, _11357_);
  and (_11363_, _08770_, _07923_);
  or (_11364_, _11363_, _11327_);
  or (_11365_, _11364_, _07198_);
  and (_11366_, _11365_, _11362_);
  or (_11367_, _11366_, _06367_);
  and (_11368_, _08988_, _07923_);
  or (_11369_, _11368_, _11327_);
  or (_11370_, _11369_, _07218_);
  and (_11371_, _11370_, _07216_);
  and (_11372_, _11371_, _11367_);
  or (_11373_, _11372_, _11330_);
  and (_11374_, _11373_, _07213_);
  or (_11375_, _11327_, _08007_);
  and (_11376_, _11364_, _06366_);
  and (_11377_, _11376_, _11375_);
  or (_11378_, _11377_, _11374_);
  and (_11379_, _11378_, _07210_);
  and (_11380_, _11338_, _06541_);
  and (_11381_, _11380_, _11375_);
  or (_11382_, _11381_, _06383_);
  or (_11383_, _11382_, _11379_);
  and (_11384_, _08985_, _07923_);
  or (_11385_, _11327_, _07231_);
  or (_11386_, _11385_, _11384_);
  and (_11387_, _11386_, _07229_);
  and (_11388_, _11387_, _11383_);
  nor (_11389_, _08508_, _11326_);
  or (_11390_, _11389_, _11327_);
  and (_11391_, _11390_, _06528_);
  or (_11392_, _11391_, _06563_);
  or (_11393_, _11392_, _11388_);
  or (_11394_, _11335_, _07241_);
  and (_11395_, _11394_, _06189_);
  and (_11396_, _11395_, _11393_);
  and (_11397_, _08503_, _07923_);
  or (_11398_, _11397_, _11327_);
  and (_11399_, _11398_, _06188_);
  or (_11400_, _11399_, _01456_);
  or (_11401_, _11400_, _11396_);
  or (_11402_, _01452_, \oc8051_golden_model_1.PCON [7]);
  and (_11403_, _11402_, _43223_);
  and (_41180_, _11403_, _11401_);
  not (_11404_, _07885_);
  and (_11405_, _11404_, \oc8051_golden_model_1.TMOD [7]);
  and (_11406_, _08509_, _07885_);
  or (_11407_, _11406_, _11405_);
  and (_11408_, _11407_, _06533_);
  and (_11409_, _08685_, _07885_);
  or (_11410_, _11409_, _11405_);
  or (_11411_, _11410_, _06252_);
  and (_11412_, _07885_, \oc8051_golden_model_1.ACC [7]);
  or (_11413_, _11412_, _11405_);
  and (_11414_, _11413_, _07123_);
  and (_11415_, _07124_, \oc8051_golden_model_1.TMOD [7]);
  or (_11416_, _11415_, _06251_);
  or (_11417_, _11416_, _11414_);
  and (_11418_, _11417_, _07142_);
  and (_11419_, _11418_, _11411_);
  nor (_11420_, _08004_, _11404_);
  or (_11421_, _11420_, _11405_);
  and (_11422_, _11421_, _06468_);
  or (_11423_, _11422_, _11419_);
  and (_11424_, _11423_, _06801_);
  and (_11425_, _11413_, _06466_);
  or (_11426_, _11425_, _07187_);
  or (_11427_, _11426_, _11424_);
  or (_11428_, _11421_, _07188_);
  and (_11429_, _11428_, _11427_);
  or (_11430_, _11429_, _07182_);
  and (_11431_, _08671_, _07885_);
  or (_11432_, _11405_, _07183_);
  or (_11433_, _11432_, _11431_);
  and (_11434_, _11433_, _06336_);
  and (_11435_, _11434_, _11430_);
  and (_11436_, _08966_, _07885_);
  or (_11437_, _11436_, _11405_);
  and (_11438_, _11437_, _05968_);
  or (_11439_, _11438_, _06371_);
  or (_11440_, _11439_, _11435_);
  and (_11441_, _08770_, _07885_);
  or (_11442_, _11441_, _11405_);
  or (_11443_, _11442_, _07198_);
  and (_11444_, _11443_, _11440_);
  or (_11445_, _11444_, _06367_);
  and (_11446_, _08988_, _07885_);
  or (_11447_, _11446_, _11405_);
  or (_11448_, _11447_, _07218_);
  and (_11449_, _11448_, _07216_);
  and (_11450_, _11449_, _11445_);
  or (_11451_, _11450_, _11408_);
  and (_11452_, _11451_, _07213_);
  or (_11453_, _11405_, _08007_);
  and (_11454_, _11442_, _06366_);
  and (_11455_, _11454_, _11453_);
  or (_11456_, _11455_, _11452_);
  and (_11457_, _11456_, _07210_);
  and (_11458_, _11413_, _06541_);
  and (_11459_, _11458_, _11453_);
  or (_11460_, _11459_, _06383_);
  or (_11461_, _11460_, _11457_);
  and (_11462_, _08985_, _07885_);
  or (_11463_, _11405_, _07231_);
  or (_11464_, _11463_, _11462_);
  and (_11465_, _11464_, _07229_);
  and (_11466_, _11465_, _11461_);
  nor (_11467_, _08508_, _11404_);
  or (_11468_, _11467_, _11405_);
  and (_11469_, _11468_, _06528_);
  or (_11470_, _11469_, _06563_);
  or (_11471_, _11470_, _11466_);
  or (_11472_, _11410_, _07241_);
  and (_11473_, _11472_, _06189_);
  and (_11474_, _11473_, _11471_);
  and (_11475_, _08503_, _07885_);
  or (_11476_, _11475_, _11405_);
  and (_11477_, _11476_, _06188_);
  or (_11478_, _11477_, _01456_);
  or (_11479_, _11478_, _11474_);
  or (_11480_, _01452_, \oc8051_golden_model_1.TMOD [7]);
  and (_11481_, _11480_, _43223_);
  and (_41181_, _11481_, _11479_);
  not (_11482_, \oc8051_golden_model_1.DPL [7]);
  nor (_11483_, _07932_, _11482_);
  and (_11484_, _08509_, _07932_);
  or (_11485_, _11484_, _11483_);
  and (_11486_, _11485_, _06533_);
  not (_11487_, _07932_);
  nor (_11488_, _08004_, _11487_);
  or (_11489_, _11488_, _11483_);
  or (_11490_, _11489_, _07188_);
  and (_11491_, _08685_, _07932_);
  or (_11492_, _11491_, _11483_);
  or (_11493_, _11492_, _06252_);
  and (_11494_, _07932_, \oc8051_golden_model_1.ACC [7]);
  or (_11495_, _11494_, _11483_);
  and (_11496_, _11495_, _07123_);
  nor (_11497_, _07123_, _11482_);
  or (_11498_, _11497_, _06251_);
  or (_11499_, _11498_, _11496_);
  and (_11500_, _11499_, _07142_);
  and (_11501_, _11500_, _11493_);
  and (_11502_, _11489_, _06468_);
  or (_11503_, _11502_, _06466_);
  or (_11504_, _11503_, _11501_);
  and (_11505_, _06490_, _05934_);
  not (_11506_, _11505_);
  or (_11507_, _11495_, _06801_);
  and (_11508_, _11507_, _11506_);
  and (_11509_, _11508_, _11504_);
  and (_11510_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_11511_, _11510_, \oc8051_golden_model_1.DPL [2]);
  and (_11512_, _11511_, \oc8051_golden_model_1.DPL [3]);
  and (_11513_, _11512_, \oc8051_golden_model_1.DPL [4]);
  and (_11514_, _11513_, \oc8051_golden_model_1.DPL [5]);
  and (_11515_, _11514_, \oc8051_golden_model_1.DPL [6]);
  nor (_11516_, _11515_, \oc8051_golden_model_1.DPL [7]);
  and (_11517_, _11515_, \oc8051_golden_model_1.DPL [7]);
  nor (_11518_, _11517_, _11516_);
  and (_11519_, _11518_, _11505_);
  or (_11520_, _11519_, _11509_);
  and (_11521_, _11520_, _06370_);
  nor (_11522_, _08769_, _06370_);
  or (_11523_, _11522_, _07187_);
  or (_11524_, _11523_, _11521_);
  and (_11525_, _11524_, _11490_);
  or (_11526_, _11525_, _07182_);
  and (_11527_, _08671_, _07932_);
  or (_11528_, _11483_, _07183_);
  or (_11529_, _11528_, _11527_);
  and (_11530_, _11529_, _06336_);
  and (_11531_, _11530_, _11526_);
  and (_11532_, _08966_, _07932_);
  or (_11533_, _11532_, _11483_);
  and (_11534_, _11533_, _05968_);
  or (_11535_, _11534_, _06371_);
  or (_11536_, _11535_, _11531_);
  and (_11537_, _08770_, _07932_);
  or (_11538_, _11537_, _11483_);
  or (_11539_, _11538_, _07198_);
  and (_11540_, _11539_, _11536_);
  or (_11541_, _11540_, _06367_);
  and (_11542_, _08988_, _07932_);
  or (_11543_, _11542_, _11483_);
  or (_11544_, _11543_, _07218_);
  and (_11545_, _11544_, _07216_);
  and (_11546_, _11545_, _11541_);
  or (_11547_, _11546_, _11486_);
  and (_11548_, _11547_, _07213_);
  or (_11549_, _11483_, _08007_);
  and (_11550_, _11538_, _06366_);
  and (_11551_, _11550_, _11549_);
  or (_11552_, _11551_, _11548_);
  and (_11553_, _11552_, _07210_);
  and (_11554_, _11495_, _06541_);
  and (_11555_, _11554_, _11549_);
  or (_11556_, _11555_, _06383_);
  or (_11557_, _11556_, _11553_);
  and (_11558_, _08985_, _07932_);
  or (_11559_, _11483_, _07231_);
  or (_11560_, _11559_, _11558_);
  and (_11561_, _11560_, _07229_);
  and (_11562_, _11561_, _11557_);
  nor (_11563_, _08508_, _11487_);
  or (_11564_, _11563_, _11483_);
  and (_11565_, _11564_, _06528_);
  or (_11566_, _11565_, _06563_);
  or (_11567_, _11566_, _11562_);
  or (_11568_, _11492_, _07241_);
  and (_11569_, _11568_, _06189_);
  and (_11570_, _11569_, _11567_);
  and (_11571_, _08503_, _07932_);
  or (_11572_, _11571_, _11483_);
  and (_11573_, _11572_, _06188_);
  or (_11574_, _11573_, _01456_);
  or (_11575_, _11574_, _11570_);
  or (_11576_, _01452_, \oc8051_golden_model_1.DPL [7]);
  and (_11577_, _11576_, _43223_);
  and (_41182_, _11577_, _11575_);
  not (_11578_, \oc8051_golden_model_1.DPH [7]);
  nor (_11579_, _07935_, _11578_);
  and (_11580_, _08509_, _08151_);
  or (_11581_, _11580_, _11579_);
  and (_11582_, _11581_, _06533_);
  not (_11583_, _08151_);
  nor (_11584_, _08004_, _11583_);
  or (_11585_, _11584_, _11579_);
  or (_11586_, _11585_, _07188_);
  and (_11587_, _08685_, _08151_);
  or (_11588_, _11587_, _11579_);
  or (_11589_, _11588_, _06252_);
  and (_11590_, _07935_, \oc8051_golden_model_1.ACC [7]);
  or (_11591_, _11590_, _11579_);
  and (_11592_, _11591_, _07123_);
  nor (_11593_, _07123_, _11578_);
  or (_11594_, _11593_, _06251_);
  or (_11595_, _11594_, _11592_);
  and (_11596_, _11595_, _07142_);
  and (_11597_, _11596_, _11589_);
  and (_11598_, _11585_, _06468_);
  or (_11599_, _11598_, _06466_);
  or (_11600_, _11599_, _11597_);
  or (_11601_, _11591_, _06801_);
  and (_11602_, _11601_, _11506_);
  and (_11603_, _11602_, _11600_);
  and (_11604_, _11517_, \oc8051_golden_model_1.DPH [0]);
  and (_11605_, _11604_, \oc8051_golden_model_1.DPH [1]);
  and (_11606_, _11605_, \oc8051_golden_model_1.DPH [2]);
  and (_11607_, _11606_, \oc8051_golden_model_1.DPH [3]);
  and (_11608_, _11607_, \oc8051_golden_model_1.DPH [4]);
  and (_11609_, _11608_, \oc8051_golden_model_1.DPH [5]);
  and (_11610_, _11609_, \oc8051_golden_model_1.DPH [6]);
  nand (_11611_, _11610_, \oc8051_golden_model_1.DPH [7]);
  or (_11612_, _11610_, \oc8051_golden_model_1.DPH [7]);
  and (_11613_, _11612_, _11611_);
  and (_11614_, _11613_, _11505_);
  or (_11615_, _11614_, _11603_);
  and (_11616_, _11615_, _06370_);
  and (_11617_, _06369_, _06187_);
  or (_11618_, _11617_, _07187_);
  or (_11619_, _11618_, _11616_);
  and (_11620_, _11619_, _11586_);
  or (_11621_, _11620_, _07182_);
  or (_11622_, _11579_, _07183_);
  and (_11623_, _08671_, _07935_);
  or (_11624_, _11623_, _11622_);
  and (_11625_, _11624_, _06336_);
  and (_11626_, _11625_, _11621_);
  and (_11627_, _08966_, _07935_);
  or (_11628_, _11627_, _11579_);
  and (_11629_, _11628_, _05968_);
  or (_11630_, _11629_, _06371_);
  or (_11631_, _11630_, _11626_);
  and (_11632_, _08770_, _07935_);
  or (_11633_, _11632_, _11579_);
  or (_11634_, _11633_, _07198_);
  and (_11635_, _11634_, _11631_);
  or (_11636_, _11635_, _06367_);
  and (_11637_, _08988_, _07935_);
  or (_11638_, _11637_, _11579_);
  or (_11639_, _11638_, _07218_);
  and (_11640_, _11639_, _07216_);
  and (_11641_, _11640_, _11636_);
  or (_11642_, _11641_, _11582_);
  and (_11643_, _11642_, _07213_);
  or (_11644_, _11579_, _08007_);
  and (_11645_, _11633_, _06366_);
  and (_11646_, _11645_, _11644_);
  or (_11647_, _11646_, _11643_);
  and (_11648_, _11647_, _07210_);
  and (_11649_, _11591_, _06541_);
  and (_11650_, _11649_, _11644_);
  or (_11651_, _11650_, _06383_);
  or (_11652_, _11651_, _11648_);
  and (_11653_, _08985_, _08151_);
  or (_11654_, _11579_, _07231_);
  or (_11655_, _11654_, _11653_);
  and (_11656_, _11655_, _07229_);
  and (_11657_, _11656_, _11652_);
  nor (_11658_, _08508_, _11583_);
  or (_11659_, _11658_, _11579_);
  and (_11660_, _11659_, _06528_);
  or (_11661_, _11660_, _06563_);
  or (_11662_, _11661_, _11657_);
  or (_11663_, _11588_, _07241_);
  and (_11664_, _11663_, _06189_);
  and (_11665_, _11664_, _11662_);
  and (_11666_, _08503_, _08151_);
  or (_11667_, _11666_, _11579_);
  and (_11668_, _11667_, _06188_);
  or (_11669_, _11668_, _01456_);
  or (_11670_, _11669_, _11665_);
  or (_11671_, _01452_, \oc8051_golden_model_1.DPH [7]);
  and (_11672_, _11671_, _43223_);
  and (_41185_, _11672_, _11670_);
  not (_11673_, _07940_);
  and (_11674_, _11673_, \oc8051_golden_model_1.TL1 [7]);
  and (_11675_, _08509_, _07940_);
  or (_11676_, _11675_, _11674_);
  and (_11677_, _11676_, _06533_);
  nor (_11678_, _08004_, _11673_);
  or (_11679_, _11678_, _11674_);
  or (_11680_, _11679_, _07188_);
  and (_11681_, _08685_, _07940_);
  or (_11682_, _11681_, _11674_);
  or (_11683_, _11682_, _06252_);
  and (_11684_, _07940_, \oc8051_golden_model_1.ACC [7]);
  or (_11685_, _11684_, _11674_);
  and (_11686_, _11685_, _07123_);
  and (_11687_, _07124_, \oc8051_golden_model_1.TL1 [7]);
  or (_11688_, _11687_, _06251_);
  or (_11689_, _11688_, _11686_);
  and (_11690_, _11689_, _07142_);
  and (_11691_, _11690_, _11683_);
  and (_11692_, _11679_, _06468_);
  or (_11693_, _11692_, _11691_);
  and (_11694_, _11693_, _06801_);
  and (_11695_, _11685_, _06466_);
  or (_11696_, _11695_, _07187_);
  or (_11697_, _11696_, _11694_);
  and (_11698_, _11697_, _11680_);
  or (_11699_, _11698_, _07182_);
  and (_11700_, _08671_, _07940_);
  or (_11701_, _11674_, _07183_);
  or (_11702_, _11701_, _11700_);
  and (_11703_, _11702_, _06336_);
  and (_11704_, _11703_, _11699_);
  and (_11705_, _08966_, _07940_);
  or (_11706_, _11705_, _11674_);
  and (_11707_, _11706_, _05968_);
  or (_11708_, _11707_, _06371_);
  or (_11709_, _11708_, _11704_);
  and (_11710_, _08770_, _07940_);
  or (_11711_, _11710_, _11674_);
  or (_11712_, _11711_, _07198_);
  and (_11713_, _11712_, _11709_);
  or (_11714_, _11713_, _06367_);
  and (_11715_, _08988_, _07940_);
  or (_11716_, _11715_, _11674_);
  or (_11717_, _11716_, _07218_);
  and (_11718_, _11717_, _07216_);
  and (_11719_, _11718_, _11714_);
  or (_11720_, _11719_, _11677_);
  and (_11721_, _11720_, _07213_);
  or (_11722_, _11674_, _08007_);
  and (_11723_, _11711_, _06366_);
  and (_11724_, _11723_, _11722_);
  or (_11725_, _11724_, _11721_);
  and (_11726_, _11725_, _07210_);
  and (_11727_, _11685_, _06541_);
  and (_11728_, _11727_, _11722_);
  or (_11729_, _11728_, _06383_);
  or (_11730_, _11729_, _11726_);
  and (_11731_, _08985_, _07940_);
  or (_11732_, _11674_, _07231_);
  or (_11733_, _11732_, _11731_);
  and (_11734_, _11733_, _07229_);
  and (_11735_, _11734_, _11730_);
  nor (_11736_, _08508_, _11673_);
  or (_11737_, _11736_, _11674_);
  and (_11738_, _11737_, _06528_);
  or (_11739_, _11738_, _06563_);
  or (_11740_, _11739_, _11735_);
  or (_11741_, _11682_, _07241_);
  and (_11742_, _11741_, _06189_);
  and (_11743_, _11742_, _11740_);
  and (_11744_, _08503_, _07940_);
  or (_11745_, _11744_, _11674_);
  and (_11746_, _11745_, _06188_);
  or (_11747_, _11746_, _01456_);
  or (_11748_, _11747_, _11743_);
  or (_11749_, _01452_, \oc8051_golden_model_1.TL1 [7]);
  and (_11750_, _11749_, _43223_);
  and (_41186_, _11750_, _11748_);
  not (_11751_, _07893_);
  and (_11752_, _11751_, \oc8051_golden_model_1.TL0 [7]);
  and (_11753_, _08509_, _08139_);
  or (_11754_, _11753_, _11752_);
  and (_11755_, _11754_, _06533_);
  and (_11756_, _08685_, _08139_);
  or (_11757_, _11756_, _11752_);
  or (_11758_, _11757_, _06252_);
  and (_11759_, _07893_, \oc8051_golden_model_1.ACC [7]);
  or (_11760_, _11759_, _11752_);
  and (_11761_, _11760_, _07123_);
  and (_11762_, _07124_, \oc8051_golden_model_1.TL0 [7]);
  or (_11763_, _11762_, _06251_);
  or (_11764_, _11763_, _11761_);
  and (_11765_, _11764_, _07142_);
  and (_11766_, _11765_, _11758_);
  not (_11767_, _08139_);
  nor (_11768_, _08004_, _11767_);
  or (_11769_, _11768_, _11752_);
  and (_11770_, _11769_, _06468_);
  or (_11771_, _11770_, _11766_);
  and (_11772_, _11771_, _06801_);
  and (_11773_, _11760_, _06466_);
  or (_11774_, _11773_, _07187_);
  or (_11775_, _11774_, _11772_);
  or (_11776_, _11769_, _07188_);
  and (_11777_, _11776_, _11775_);
  or (_11778_, _11777_, _07182_);
  or (_11779_, _11752_, _07183_);
  and (_11780_, _08671_, _07893_);
  or (_11781_, _11780_, _11779_);
  and (_11782_, _11781_, _06336_);
  and (_11783_, _11782_, _11778_);
  and (_11784_, _08966_, _07893_);
  or (_11785_, _11784_, _11752_);
  and (_11786_, _11785_, _05968_);
  or (_11787_, _11786_, _06371_);
  or (_11788_, _11787_, _11783_);
  and (_11789_, _08770_, _07893_);
  or (_11790_, _11789_, _11752_);
  or (_11791_, _11790_, _07198_);
  and (_11792_, _11791_, _11788_);
  or (_11793_, _11792_, _06367_);
  and (_11794_, _08988_, _07893_);
  or (_11795_, _11794_, _11752_);
  or (_11796_, _11795_, _07218_);
  and (_11797_, _11796_, _07216_);
  and (_11798_, _11797_, _11793_);
  or (_11799_, _11798_, _11755_);
  and (_11800_, _11799_, _07213_);
  or (_11801_, _11752_, _08007_);
  and (_11802_, _11790_, _06366_);
  and (_11803_, _11802_, _11801_);
  or (_11804_, _11803_, _11800_);
  and (_11805_, _11804_, _07210_);
  and (_11806_, _11760_, _06541_);
  and (_11807_, _11806_, _11801_);
  or (_11808_, _11807_, _06383_);
  or (_11809_, _11808_, _11805_);
  and (_11810_, _08985_, _08139_);
  or (_11811_, _11752_, _07231_);
  or (_11812_, _11811_, _11810_);
  and (_11813_, _11812_, _07229_);
  and (_11814_, _11813_, _11809_);
  nor (_11815_, _08508_, _11767_);
  or (_11816_, _11815_, _11752_);
  and (_11817_, _11816_, _06528_);
  or (_11818_, _11817_, _06563_);
  or (_11819_, _11818_, _11814_);
  or (_11820_, _11757_, _07241_);
  and (_11821_, _11820_, _06189_);
  and (_11822_, _11821_, _11819_);
  and (_11823_, _08503_, _08139_);
  or (_11824_, _11823_, _11752_);
  and (_11825_, _11824_, _06188_);
  or (_11826_, _11825_, _01456_);
  or (_11827_, _11826_, _11822_);
  or (_11828_, _01452_, \oc8051_golden_model_1.TL0 [7]);
  and (_11829_, _11828_, _43223_);
  and (_41187_, _11829_, _11827_);
  and (_11830_, _01456_, \oc8051_golden_model_1.TCON [7]);
  not (_11831_, _07897_);
  and (_11832_, _11831_, \oc8051_golden_model_1.TCON [7]);
  and (_11833_, _08509_, _07897_);
  or (_11834_, _11833_, _11832_);
  and (_11835_, _11834_, _06533_);
  nor (_11836_, _08004_, _11831_);
  or (_11837_, _11836_, _11832_);
  or (_11838_, _11837_, _07188_);
  or (_11839_, _11837_, _07142_);
  and (_11840_, _08685_, _07897_);
  or (_11841_, _11840_, _11832_);
  or (_11842_, _11841_, _06252_);
  and (_11843_, _07897_, \oc8051_golden_model_1.ACC [7]);
  or (_11844_, _11843_, _11832_);
  and (_11845_, _11844_, _07123_);
  and (_11846_, _07124_, \oc8051_golden_model_1.TCON [7]);
  or (_11847_, _11846_, _06251_);
  or (_11848_, _11847_, _11845_);
  and (_11849_, _11848_, _06476_);
  and (_11850_, _11849_, _11842_);
  not (_11851_, _08528_);
  and (_11852_, _11851_, \oc8051_golden_model_1.TCON [7]);
  and (_11853_, _08560_, _08528_);
  or (_11854_, _11853_, _11852_);
  and (_11855_, _11854_, _06475_);
  or (_11856_, _11855_, _06468_);
  or (_11857_, _11856_, _11850_);
  and (_11858_, _11857_, _11839_);
  or (_11859_, _11858_, _06466_);
  or (_11860_, _11844_, _06801_);
  and (_11861_, _11860_, _06484_);
  and (_11862_, _11861_, _11859_);
  and (_11863_, _08698_, _08528_);
  or (_11864_, _11863_, _11852_);
  and (_11865_, _11864_, _06483_);
  or (_11866_, _11865_, _11862_);
  and (_11867_, _11866_, _07164_);
  and (_11868_, _08707_, _08528_);
  or (_11869_, _11868_, _11852_);
  and (_11870_, _11869_, _06461_);
  or (_11871_, _11870_, _11867_);
  and (_11872_, _11871_, _06242_);
  and (_11873_, _08726_, _08528_);
  or (_11874_, _11873_, _11852_);
  and (_11875_, _11874_, _06241_);
  or (_11876_, _11875_, _07187_);
  or (_11877_, _11876_, _11872_);
  and (_11878_, _11877_, _11838_);
  or (_11879_, _11878_, _07182_);
  and (_11880_, _08671_, _07897_);
  or (_11881_, _11832_, _07183_);
  or (_11882_, _11881_, _11880_);
  and (_11883_, _11882_, _06336_);
  and (_11884_, _11883_, _11879_);
  and (_11885_, _08966_, _07897_);
  or (_11886_, _11885_, _11832_);
  and (_11887_, _11886_, _05968_);
  or (_11888_, _11887_, _06371_);
  or (_11889_, _11888_, _11884_);
  and (_11890_, _08770_, _07897_);
  or (_11891_, _11890_, _11832_);
  or (_11892_, _11891_, _07198_);
  and (_11893_, _11892_, _11889_);
  or (_11894_, _11893_, _06367_);
  and (_11895_, _08988_, _07897_);
  or (_11896_, _11895_, _11832_);
  or (_11897_, _11896_, _07218_);
  and (_11898_, _11897_, _07216_);
  and (_11899_, _11898_, _11894_);
  or (_11900_, _11899_, _11835_);
  and (_11901_, _11900_, _07213_);
  or (_11902_, _11832_, _08007_);
  and (_11903_, _11891_, _06366_);
  and (_11904_, _11903_, _11902_);
  or (_11905_, _11904_, _11901_);
  and (_11906_, _11905_, _07210_);
  and (_11907_, _11844_, _06541_);
  and (_11908_, _11907_, _11902_);
  or (_11909_, _11908_, _06383_);
  or (_11910_, _11909_, _11906_);
  and (_11911_, _08985_, _07897_);
  or (_11912_, _11832_, _07231_);
  or (_11913_, _11912_, _11911_);
  and (_11914_, _11913_, _07229_);
  and (_11915_, _11914_, _11910_);
  nor (_11916_, _08508_, _11831_);
  or (_11917_, _11916_, _11832_);
  and (_11918_, _11917_, _06528_);
  or (_11919_, _11918_, _06563_);
  or (_11920_, _11919_, _11915_);
  or (_11921_, _11841_, _07241_);
  and (_11922_, _11921_, _06571_);
  and (_11923_, _11922_, _11920_);
  and (_11924_, _11864_, _06199_);
  or (_11925_, _11924_, _06188_);
  or (_11926_, _11925_, _11923_);
  and (_11927_, _08503_, _07897_);
  or (_11928_, _11832_, _06189_);
  or (_11929_, _11928_, _11927_);
  and (_11930_, _11929_, _01452_);
  and (_11931_, _11930_, _11926_);
  or (_11932_, _11931_, _11830_);
  and (_41188_, _11932_, _43223_);
  not (_11933_, _07879_);
  and (_11934_, _11933_, \oc8051_golden_model_1.TH1 [7]);
  and (_11935_, _08509_, _07879_);
  or (_11936_, _11935_, _11934_);
  and (_11937_, _11936_, _06533_);
  and (_11938_, _08685_, _07879_);
  or (_11939_, _11938_, _11934_);
  or (_11940_, _11939_, _06252_);
  and (_11941_, _07879_, \oc8051_golden_model_1.ACC [7]);
  or (_11942_, _11941_, _11934_);
  and (_11943_, _11942_, _07123_);
  and (_11944_, _07124_, \oc8051_golden_model_1.TH1 [7]);
  or (_11945_, _11944_, _06251_);
  or (_11946_, _11945_, _11943_);
  and (_11947_, _11946_, _07142_);
  and (_11948_, _11947_, _11940_);
  nor (_11949_, _08004_, _11933_);
  or (_11950_, _11949_, _11934_);
  and (_11951_, _11950_, _06468_);
  or (_11952_, _11951_, _11948_);
  and (_11953_, _11952_, _06801_);
  and (_11954_, _11942_, _06466_);
  or (_11955_, _11954_, _07187_);
  or (_11956_, _11955_, _11953_);
  or (_11957_, _11950_, _07188_);
  and (_11958_, _11957_, _11956_);
  or (_11959_, _11958_, _07182_);
  and (_11960_, _08671_, _07879_);
  or (_11961_, _11934_, _07183_);
  or (_11962_, _11961_, _11960_);
  and (_11963_, _11962_, _06336_);
  and (_11964_, _11963_, _11959_);
  and (_11965_, _08966_, _07879_);
  or (_11966_, _11965_, _11934_);
  and (_11967_, _11966_, _05968_);
  or (_11968_, _11967_, _06371_);
  or (_11969_, _11968_, _11964_);
  and (_11970_, _08770_, _07879_);
  or (_11971_, _11970_, _11934_);
  or (_11972_, _11971_, _07198_);
  and (_11973_, _11972_, _11969_);
  or (_11974_, _11973_, _06367_);
  and (_11975_, _08988_, _07879_);
  or (_11976_, _11975_, _11934_);
  or (_11977_, _11976_, _07218_);
  and (_11978_, _11977_, _07216_);
  and (_11979_, _11978_, _11974_);
  or (_11980_, _11979_, _11937_);
  and (_11981_, _11980_, _07213_);
  or (_11982_, _11934_, _08007_);
  and (_11983_, _11971_, _06366_);
  and (_11984_, _11983_, _11982_);
  or (_11985_, _11984_, _11981_);
  and (_11986_, _11985_, _07210_);
  and (_11987_, _11942_, _06541_);
  and (_11988_, _11987_, _11982_);
  or (_11989_, _11988_, _06383_);
  or (_11990_, _11989_, _11986_);
  and (_11991_, _08985_, _07879_);
  or (_11992_, _11934_, _07231_);
  or (_11993_, _11992_, _11991_);
  and (_11994_, _11993_, _07229_);
  and (_11995_, _11994_, _11990_);
  nor (_11996_, _08508_, _11933_);
  or (_11997_, _11996_, _11934_);
  and (_11998_, _11997_, _06528_);
  or (_11999_, _11998_, _06563_);
  or (_12000_, _11999_, _11995_);
  or (_12001_, _11939_, _07241_);
  and (_12002_, _12001_, _06189_);
  and (_12003_, _12002_, _12000_);
  and (_12004_, _08503_, _07879_);
  or (_12005_, _12004_, _11934_);
  and (_12006_, _12005_, _06188_);
  or (_12007_, _12006_, _01456_);
  or (_12008_, _12007_, _12003_);
  or (_12009_, _01452_, \oc8051_golden_model_1.TH1 [7]);
  and (_12010_, _12009_, _43223_);
  and (_41189_, _12010_, _12008_);
  not (_12011_, _07889_);
  and (_12012_, _12011_, \oc8051_golden_model_1.TH0 [7]);
  and (_12013_, _08509_, _07889_);
  or (_12014_, _12013_, _12012_);
  and (_12015_, _12014_, _06533_);
  nor (_12016_, _08004_, _12011_);
  or (_12017_, _12016_, _12012_);
  or (_12018_, _12017_, _07188_);
  and (_12019_, _08685_, _07889_);
  or (_12020_, _12019_, _12012_);
  or (_12021_, _12020_, _06252_);
  and (_12022_, _07889_, \oc8051_golden_model_1.ACC [7]);
  or (_12023_, _12022_, _12012_);
  and (_12024_, _12023_, _07123_);
  and (_12025_, _07124_, \oc8051_golden_model_1.TH0 [7]);
  or (_12026_, _12025_, _06251_);
  or (_12027_, _12026_, _12024_);
  and (_12028_, _12027_, _07142_);
  and (_12029_, _12028_, _12021_);
  and (_12030_, _12017_, _06468_);
  or (_12031_, _12030_, _12029_);
  and (_12032_, _12031_, _06801_);
  and (_12033_, _12023_, _06466_);
  or (_12034_, _12033_, _07187_);
  or (_12035_, _12034_, _12032_);
  and (_12036_, _12035_, _12018_);
  or (_12037_, _12036_, _07182_);
  and (_12038_, _08671_, _07889_);
  or (_12039_, _12012_, _07183_);
  or (_12040_, _12039_, _12038_);
  and (_12041_, _12040_, _06336_);
  and (_12042_, _12041_, _12037_);
  and (_12043_, _08966_, _07889_);
  or (_12044_, _12043_, _12012_);
  and (_12045_, _12044_, _05968_);
  or (_12046_, _12045_, _06371_);
  or (_12047_, _12046_, _12042_);
  and (_12048_, _08770_, _07889_);
  or (_12049_, _12048_, _12012_);
  or (_12050_, _12049_, _07198_);
  and (_12051_, _12050_, _12047_);
  or (_12052_, _12051_, _06367_);
  and (_12053_, _08988_, _07889_);
  or (_12054_, _12053_, _12012_);
  or (_12055_, _12054_, _07218_);
  and (_12056_, _12055_, _07216_);
  and (_12057_, _12056_, _12052_);
  or (_12058_, _12057_, _12015_);
  and (_12059_, _12058_, _07213_);
  or (_12060_, _12012_, _08007_);
  and (_12061_, _12049_, _06366_);
  and (_12062_, _12061_, _12060_);
  or (_12063_, _12062_, _12059_);
  and (_12064_, _12063_, _07210_);
  and (_12065_, _12023_, _06541_);
  and (_12066_, _12065_, _12060_);
  or (_12067_, _12066_, _06383_);
  or (_12068_, _12067_, _12064_);
  and (_12069_, _08985_, _07889_);
  or (_12070_, _12012_, _07231_);
  or (_12071_, _12070_, _12069_);
  and (_12072_, _12071_, _07229_);
  and (_12073_, _12072_, _12068_);
  nor (_12074_, _08508_, _12011_);
  or (_12075_, _12074_, _12012_);
  and (_12076_, _12075_, _06528_);
  or (_12077_, _12076_, _06563_);
  or (_12078_, _12077_, _12073_);
  or (_12079_, _12020_, _07241_);
  and (_12080_, _12079_, _06189_);
  and (_12081_, _12080_, _12078_);
  and (_12082_, _08503_, _07889_);
  or (_12083_, _12082_, _12012_);
  and (_12084_, _12083_, _06188_);
  or (_12085_, _12084_, _01456_);
  or (_12086_, _12085_, _12081_);
  or (_12087_, _01452_, \oc8051_golden_model_1.TH0 [7]);
  and (_12088_, _12087_, _43223_);
  and (_41191_, _12088_, _12086_);
  not (_12089_, _05924_);
  not (_12090_, \oc8051_golden_model_1.PC [15]);
  and (_12091_, _08514_, _05571_);
  and (_12092_, _12091_, \oc8051_golden_model_1.PC [7]);
  and (_12093_, _12092_, \oc8051_golden_model_1.PC [8]);
  and (_12094_, _12093_, \oc8051_golden_model_1.PC [9]);
  and (_12095_, _12094_, \oc8051_golden_model_1.PC [10]);
  and (_12096_, _12095_, \oc8051_golden_model_1.PC [11]);
  and (_12097_, _12096_, \oc8051_golden_model_1.PC [12]);
  and (_12098_, _12097_, \oc8051_golden_model_1.PC [13]);
  nand (_12099_, _12098_, \oc8051_golden_model_1.PC [14]);
  nand (_12100_, _12099_, _12090_);
  or (_12101_, _12099_, _12090_);
  and (_12102_, _12101_, _12100_);
  or (_12103_, _05923_, _05965_);
  not (_12104_, _12103_);
  nor (_12105_, _12104_, _11156_);
  or (_12106_, _12105_, _12102_);
  nor (_12107_, _09432_, \oc8051_golden_model_1.PC [14]);
  nor (_12108_, _12107_, _09433_);
  and (_12109_, _12108_, _06187_);
  nor (_12110_, _12108_, _06187_);
  nor (_12111_, _12110_, _12109_);
  nor (_12112_, _09431_, \oc8051_golden_model_1.PC [13]);
  nor (_12113_, _12112_, _09432_);
  and (_12114_, _12113_, _06187_);
  nor (_12115_, _12113_, _06187_);
  nor (_12116_, _09430_, \oc8051_golden_model_1.PC [12]);
  nor (_12117_, _12116_, _09431_);
  and (_12118_, _12117_, _06187_);
  not (_12119_, \oc8051_golden_model_1.PC [11]);
  nor (_12120_, _09429_, _12119_);
  and (_12121_, _09429_, _12119_);
  or (_12122_, _12121_, _12120_);
  and (_12123_, _12122_, _06187_);
  nor (_12124_, _12122_, _06187_);
  nor (_12125_, _12124_, _12123_);
  nor (_12126_, _09436_, \oc8051_golden_model_1.PC [10]);
  nor (_12127_, _12126_, _09429_);
  and (_12128_, _12127_, _06187_);
  nor (_12129_, _12127_, _06187_);
  nor (_12130_, _12129_, _12128_);
  and (_12131_, _12130_, _12125_);
  nor (_12132_, _09435_, \oc8051_golden_model_1.PC [9]);
  nor (_12133_, _12132_, _09436_);
  and (_12134_, _12133_, _06187_);
  nor (_12135_, _12133_, _06187_);
  nor (_12136_, _12135_, _12134_);
  and (_12137_, _08518_, _06187_);
  nor (_12138_, _08518_, _06187_);
  and (_12139_, _08513_, _06073_);
  nor (_12140_, _12139_, \oc8051_golden_model_1.PC [6]);
  nor (_12141_, _12140_, _08515_);
  not (_12142_, _12141_);
  nor (_12143_, _12142_, _06326_);
  and (_12144_, _12142_, _06326_);
  nor (_12145_, _12144_, _12143_);
  and (_12146_, _06073_, \oc8051_golden_model_1.PC [4]);
  nor (_12147_, _12146_, \oc8051_golden_model_1.PC [5]);
  nor (_12148_, _12147_, _12139_);
  not (_12149_, _12148_);
  nor (_12150_, _12149_, _06608_);
  and (_12151_, _12149_, _06608_);
  nor (_12152_, _06073_, \oc8051_golden_model_1.PC [4]);
  nor (_12153_, _12152_, _12146_);
  not (_12154_, _12153_);
  nor (_12155_, _12154_, _06230_);
  nor (_12156_, _06292_, _06095_);
  and (_12157_, _06292_, _06095_);
  nor (_12158_, _06750_, _06019_);
  nor (_12159_, _06155_, \oc8051_golden_model_1.PC [1]);
  and (_12160_, _06799_, \oc8051_golden_model_1.PC [0]);
  and (_12161_, _06155_, \oc8051_golden_model_1.PC [1]);
  nor (_12162_, _12161_, _12159_);
  and (_12163_, _12162_, _12160_);
  nor (_12164_, _12163_, _12159_);
  and (_12165_, _06750_, _06019_);
  nor (_12166_, _12165_, _12158_);
  not (_12167_, _12166_);
  nor (_12168_, _12167_, _12164_);
  nor (_12169_, _12168_, _12158_);
  nor (_12170_, _12169_, _12157_);
  nor (_12171_, _12170_, _12156_);
  and (_12172_, _12154_, _06230_);
  nor (_12173_, _12172_, _12155_);
  not (_12174_, _12173_);
  nor (_12175_, _12174_, _12171_);
  nor (_12176_, _12175_, _12155_);
  nor (_12177_, _12176_, _12151_);
  nor (_12178_, _12177_, _12150_);
  not (_12179_, _12178_);
  and (_12180_, _12179_, _12145_);
  nor (_12181_, _12180_, _12143_);
  nor (_12182_, _12181_, _12138_);
  or (_12183_, _12182_, _12137_);
  nor (_12184_, _08516_, \oc8051_golden_model_1.PC [8]);
  nor (_12185_, _12184_, _09435_);
  and (_12186_, _12185_, _06187_);
  nor (_12187_, _12185_, _06187_);
  nor (_12188_, _12187_, _12186_);
  and (_12189_, _12188_, _12183_);
  and (_12190_, _12189_, _12136_);
  and (_12191_, _12190_, _12131_);
  nor (_12192_, _12186_, _12134_);
  not (_12193_, _12192_);
  and (_12194_, _12193_, _12131_);
  or (_12195_, _12194_, _12128_);
  or (_12196_, _12195_, _12191_);
  nor (_12197_, _12196_, _12123_);
  nor (_12198_, _12117_, _06187_);
  nor (_12199_, _12198_, _12118_);
  not (_12200_, _12199_);
  nor (_12201_, _12200_, _12197_);
  nor (_12202_, _12201_, _12118_);
  nor (_12203_, _12202_, _12115_);
  nor (_12204_, _12203_, _12114_);
  not (_12205_, _12204_);
  and (_12206_, _12205_, _12111_);
  nor (_12207_, _12206_, _12109_);
  nor (_12208_, _09443_, _06187_);
  and (_12209_, _09443_, _06187_);
  nor (_12210_, _12209_, _12208_);
  and (_12211_, _12210_, _12207_);
  nor (_12212_, _12210_, _12207_);
  or (_12213_, _12212_, _12211_);
  or (_12214_, _12213_, _10854_);
  and (_12215_, _06382_, _06198_);
  or (_12216_, _09443_, \oc8051_golden_model_1.PSW [7]);
  and (_12217_, _12216_, _12215_);
  and (_12218_, _12217_, _12214_);
  and (_12219_, _06365_, _06348_);
  not (_12220_, _12219_);
  or (_12221_, _06361_, _06358_);
  and (_12222_, _12221_, _06365_);
  and (_12223_, _06365_, _06192_);
  nor (_12224_, _12223_, _12222_);
  and (_12225_, _12224_, _12220_);
  and (_12226_, _12225_, _10962_);
  or (_12227_, _12226_, _12102_);
  nor (_12228_, _10533_, _06531_);
  not (_12229_, _12228_);
  nor (_12230_, _10929_, _10924_);
  nor (_12231_, _10919_, _10912_);
  and (_12232_, _12231_, _12230_);
  or (_12233_, _12232_, _12102_);
  or (_12234_, _09443_, _08972_);
  and (_12235_, _09427_, _05968_);
  not (_12236_, _10779_);
  nor (_12237_, _12236_, _10610_);
  or (_12238_, _12237_, _12102_);
  and (_12239_, _05967_, _06490_);
  not (_12240_, _12239_);
  nor (_12241_, _11505_, _09487_);
  and (_12242_, _12241_, _12240_);
  not (_12243_, _12242_);
  and (_12244_, _12243_, _12102_);
  and (_12245_, _06337_, _05934_);
  not (_12246_, _12245_);
  nor (_12247_, _09416_, \oc8051_golden_model_1.PC [14]);
  nor (_12248_, _12247_, _09417_);
  and (_12249_, _12248_, _08770_);
  nor (_12250_, _12248_, _08770_);
  nor (_12251_, _12250_, _12249_);
  nor (_12252_, _09415_, \oc8051_golden_model_1.PC [13]);
  nor (_12253_, _12252_, _09416_);
  nor (_12254_, _12253_, _08770_);
  and (_12255_, _12253_, _08770_);
  not (_12256_, _12255_);
  nor (_12257_, _09414_, \oc8051_golden_model_1.PC [12]);
  nor (_12258_, _12257_, _09415_);
  not (_12259_, _12258_);
  nor (_12260_, _12259_, _08769_);
  nor (_12261_, _09413_, _12119_);
  and (_12262_, _09413_, _12119_);
  or (_12263_, _12262_, _12261_);
  not (_12264_, _12263_);
  nor (_12265_, _12264_, _08769_);
  and (_12266_, _12264_, _08769_);
  nor (_12267_, _09420_, \oc8051_golden_model_1.PC [10]);
  nor (_12268_, _12267_, _09413_);
  not (_12269_, _12268_);
  nor (_12270_, _12269_, _08769_);
  and (_12271_, _12269_, _08769_);
  nor (_12272_, _12271_, _12270_);
  nor (_12273_, _09419_, \oc8051_golden_model_1.PC [9]);
  nor (_12274_, _12273_, _09420_);
  not (_12275_, _12274_);
  nor (_12276_, _12275_, _08769_);
  and (_12277_, _12275_, _08769_);
  nor (_12278_, _09361_, \oc8051_golden_model_1.PC [8]);
  nor (_12279_, _12278_, _09419_);
  not (_12280_, _12279_);
  nor (_12281_, _12280_, _08769_);
  not (_12282_, _09363_);
  nor (_12283_, _08769_, _12282_);
  and (_12284_, _08769_, _12282_);
  and (_12285_, _09359_, _08513_);
  nor (_12286_, _12285_, \oc8051_golden_model_1.PC [6]);
  nor (_12287_, _12286_, _09360_);
  not (_12288_, _12287_);
  nor (_12289_, _12288_, _08802_);
  and (_12290_, _12288_, _08802_);
  nor (_12291_, _12290_, _12289_);
  and (_12292_, _09359_, \oc8051_golden_model_1.PC [4]);
  nor (_12293_, _12292_, \oc8051_golden_model_1.PC [5]);
  nor (_12294_, _12293_, _12285_);
  not (_12295_, _12294_);
  nor (_12296_, _12295_, _08867_);
  and (_12297_, _12295_, _08867_);
  nor (_12298_, _09359_, \oc8051_golden_model_1.PC [4]);
  nor (_12299_, _12298_, _12292_);
  not (_12300_, _12299_);
  nor (_12301_, _12300_, _08834_);
  nor (_12302_, _09358_, \oc8051_golden_model_1.PC [3]);
  nor (_12303_, _12302_, _09359_);
  not (_12304_, _12303_);
  nor (_12305_, _12304_, _06458_);
  and (_12306_, _12304_, _06458_);
  and (_12307_, _05592_, _05552_);
  nor (_12308_, _12307_, _09358_);
  not (_12309_, _12308_);
  nor (_12310_, _12309_, _06651_);
  nor (_12311_, _07018_, _05978_);
  nor (_12312_, _06912_, \oc8051_golden_model_1.PC [0]);
  and (_12313_, _07018_, _05978_);
  nor (_12314_, _12313_, _12311_);
  and (_12315_, _12314_, _12312_);
  nor (_12316_, _12315_, _12311_);
  and (_12317_, _12309_, _06651_);
  nor (_12318_, _12317_, _12310_);
  not (_12319_, _12318_);
  nor (_12320_, _12319_, _12316_);
  nor (_12321_, _12320_, _12310_);
  nor (_12322_, _12321_, _12306_);
  nor (_12323_, _12322_, _12305_);
  and (_12324_, _12300_, _08834_);
  nor (_12325_, _12324_, _12301_);
  not (_12326_, _12325_);
  nor (_12327_, _12326_, _12323_);
  nor (_12328_, _12327_, _12301_);
  nor (_12329_, _12328_, _12297_);
  nor (_12330_, _12329_, _12296_);
  not (_12331_, _12330_);
  and (_12332_, _12331_, _12291_);
  nor (_12333_, _12332_, _12289_);
  nor (_12334_, _12333_, _12284_);
  or (_12335_, _12334_, _12283_);
  and (_12336_, _12280_, _08769_);
  nor (_12337_, _12336_, _12281_);
  and (_12338_, _12337_, _12335_);
  nor (_12339_, _12338_, _12281_);
  nor (_12340_, _12339_, _12277_);
  nor (_12341_, _12340_, _12276_);
  not (_12342_, _12341_);
  and (_12343_, _12342_, _12272_);
  nor (_12344_, _12343_, _12270_);
  nor (_12345_, _12344_, _12266_);
  or (_12346_, _12345_, _12265_);
  and (_12347_, _12259_, _08769_);
  nor (_12348_, _12347_, _12260_);
  and (_12349_, _12348_, _12346_);
  nor (_12350_, _12349_, _12260_);
  and (_12351_, _12350_, _12256_);
  or (_12352_, _12351_, _12254_);
  not (_12353_, _12352_);
  and (_12354_, _12353_, _12251_);
  nor (_12355_, _12354_, _12249_);
  not (_12356_, _09427_);
  and (_12357_, _12356_, _08769_);
  nor (_12358_, _12356_, _08769_);
  nor (_12359_, _12358_, _12357_);
  and (_12360_, _12359_, _12355_);
  nor (_12361_, _12359_, _12355_);
  or (_12362_, _12361_, _12360_);
  or (_12363_, _08671_, _07904_);
  and (_12364_, _12363_, _08718_);
  or (_12365_, _09067_, _06326_);
  nand (_12366_, _09067_, _06326_);
  and (_12367_, _12366_, _12365_);
  and (_12368_, _12367_, _12364_);
  nand (_12369_, _09113_, _06608_);
  or (_12370_, _09113_, _06608_);
  and (_12371_, _12370_, _12369_);
  nand (_12372_, _09159_, _06230_);
  or (_12373_, _09159_, _06230_);
  and (_12374_, _12373_, _12372_);
  and (_12375_, _12374_, _12371_);
  and (_12376_, _12375_, _12368_);
  or (_12377_, _09205_, _06292_);
  nand (_12378_, _09205_, _06292_);
  and (_12379_, _12378_, _12377_);
  or (_12380_, _09251_, _06750_);
  nand (_12381_, _09251_, _06750_);
  and (_12382_, _12381_, _12380_);
  and (_12383_, _12382_, _12379_);
  nand (_12384_, _09342_, _06802_);
  or (_12385_, _09297_, _06155_);
  nand (_12386_, _09297_, _06155_);
  and (_12387_, _12386_, _12385_);
  and (_12388_, _12387_, _12384_);
  and (_12389_, _12388_, _12383_);
  or (_12390_, _09342_, _06802_);
  and (_12391_, _12390_, _12389_);
  and (_12392_, _12391_, _12376_);
  or (_12393_, _12392_, _12362_);
  nand (_12394_, _12392_, _12356_);
  and (_12395_, _12394_, _06344_);
  and (_12396_, _12395_, _12393_);
  and (_12397_, _09443_, _06466_);
  and (_12398_, _08351_, _08301_);
  and (_12399_, _08679_, _12398_);
  and (_12400_, _08108_, _08006_);
  and (_12401_, _12400_, _08676_);
  and (_12402_, _12401_, _12399_);
  or (_12403_, _12402_, _12362_);
  nand (_12404_, _12401_, _12399_);
  or (_12405_, _12404_, _09427_);
  and (_12406_, _12405_, _12403_);
  or (_12407_, _12406_, _06252_);
  and (_12408_, _08106_, _08004_);
  and (_12409_, _12408_, _08563_);
  and (_12410_, _07120_, _07325_);
  and (_12411_, _12410_, _08564_);
  and (_12412_, _12411_, _12409_);
  and (_12413_, _12412_, _09443_);
  nand (_12414_, _12411_, _12409_);
  and (_12415_, _12414_, _12213_);
  or (_12416_, _12415_, _12413_);
  or (_12417_, _12416_, _08573_);
  not (_12418_, _06808_);
  nor (_12419_, _07480_, _07441_);
  and (_12420_, _12419_, _12418_);
  or (_12421_, _12420_, _12102_);
  nor (_12422_, _07123_, \oc8051_golden_model_1.PC [15]);
  nand (_12423_, _12422_, _12420_);
  and (_12424_, _12423_, _12421_);
  or (_12425_, _12424_, _06705_);
  nor (_12426_, _10687_, _10712_);
  and (_12427_, _12426_, _10704_);
  nor (_12428_, _07123_, _06705_);
  or (_12429_, _12428_, _09443_);
  and (_12430_, _12429_, _12427_);
  and (_12431_, _12430_, _12425_);
  not (_12432_, _12427_);
  and (_12433_, _12432_, _12102_);
  or (_12434_, _12433_, _08572_);
  or (_12435_, _12434_, _12431_);
  and (_12436_, _12435_, _07338_);
  and (_12437_, _12436_, _12417_);
  and (_12438_, _12102_, _07134_);
  or (_12439_, _12438_, _06251_);
  or (_12440_, _12439_, _12437_);
  and (_12441_, _12440_, _12407_);
  and (_12442_, _06250_, _05934_);
  nor (_12443_, _12442_, _10718_);
  not (_12444_, _12443_);
  or (_12445_, _12444_, _12441_);
  nor (_12446_, _06468_, _07474_);
  and (_12447_, _12446_, _06476_);
  or (_12448_, _12443_, _12102_);
  and (_12449_, _12448_, _12447_);
  and (_12450_, _12449_, _12445_);
  nor (_12451_, _10682_, _07153_);
  not (_12452_, _12451_);
  not (_12453_, _12447_);
  and (_12454_, _12453_, _09443_);
  or (_12455_, _12454_, _12452_);
  or (_12456_, _12455_, _12450_);
  or (_12457_, _12451_, _12102_);
  and (_12458_, _12457_, _06801_);
  and (_12459_, _12458_, _12456_);
  or (_12460_, _12459_, _12397_);
  and (_12461_, _06246_, _05934_);
  nor (_12462_, _12461_, _10759_);
  and (_12463_, _12462_, _12460_);
  not (_12464_, _12462_);
  and (_12465_, _12464_, _12102_);
  not (_12466_, _05953_);
  nor (_12467_, _06247_, _12466_);
  and (_12468_, _12467_, _06484_);
  not (_12469_, _12468_);
  or (_12470_, _12469_, _12465_);
  or (_12471_, _12470_, _12463_);
  or (_12472_, _12468_, _09443_);
  and (_12473_, _12472_, _12471_);
  not (_12474_, _06360_);
  and (_12475_, _07129_, _06337_);
  and (_12476_, _07492_, _06337_);
  nor (_12477_, _12476_, _12475_);
  and (_12478_, _12477_, _12474_);
  not (_12479_, _12478_);
  or (_12480_, _12479_, _12473_);
  not (_12481_, _08005_);
  and (_12482_, _08004_, _06187_);
  nor (_12483_, _12482_, _12481_);
  nor (_12484_, _08106_, _07742_);
  and (_12485_, _08106_, _07742_);
  nor (_12486_, _12485_, _12484_);
  and (_12487_, _12486_, _12483_);
  or (_12488_, _08209_, _07862_);
  and (_12489_, _08209_, _07862_);
  not (_12490_, _12489_);
  and (_12491_, _12490_, _12488_);
  and (_12492_, _08494_, _06244_);
  nor (_12493_, _08494_, _06244_);
  nor (_12494_, _12493_, _12492_);
  and (_12495_, _12494_, _12491_);
  and (_12496_, _12495_, _12487_);
  and (_12497_, _07713_, _06328_);
  and (_12498_, _07578_, _06751_);
  nor (_12499_, _12498_, _12497_);
  or (_12500_, _07713_, _06328_);
  or (_12501_, _07578_, _06751_);
  and (_12502_, _12501_, _12500_);
  and (_12503_, _12502_, _12499_);
  or (_12504_, _07120_, _06156_);
  and (_12505_, _07120_, _06156_);
  not (_12506_, _12505_);
  and (_12507_, _12506_, _12504_);
  nand (_12508_, _07325_, _06802_);
  or (_12509_, _07325_, _06802_);
  and (_12510_, _12509_, _12508_);
  and (_12511_, _12510_, _12507_);
  and (_12512_, _12511_, _12503_);
  and (_12513_, _12512_, _12496_);
  or (_12514_, _12513_, _12362_);
  nand (_12515_, _12513_, _12356_);
  and (_12516_, _12515_, _12514_);
  or (_12517_, _12516_, _12478_);
  and (_12518_, _12517_, _06345_);
  and (_12519_, _12518_, _12480_);
  or (_12520_, _12519_, _06338_);
  or (_12521_, _12520_, _12396_);
  not (_12522_, _06373_);
  nor (_12523_, _11210_, _11211_);
  nor (_12524_, _12523_, _11214_);
  not (_12525_, _11217_);
  nor (_12526_, _08351_, \oc8051_golden_model_1.ACC [0]);
  or (_12527_, _12526_, _11218_);
  and (_12528_, _12527_, _12525_);
  and (_12529_, _12528_, _12524_);
  nor (_12530_, _11205_, _11209_);
  nor (_12531_, _11202_, _08509_);
  and (_12532_, _12531_, _12530_);
  and (_12533_, _12532_, _12529_);
  not (_12534_, _12533_);
  and (_12535_, _12534_, _12362_);
  not (_12536_, _06338_);
  and (_12537_, _12533_, _09427_);
  or (_12538_, _12537_, _12536_);
  or (_12539_, _12538_, _12535_);
  and (_12540_, _12539_, _12522_);
  and (_12541_, _12540_, _12521_);
  nor (_12542_, _11248_, _11249_);
  nor (_12543_, _12542_, _11252_);
  and (_12544_, _06802_, _05997_);
  nor (_12545_, _12544_, _11256_);
  nor (_12546_, _12545_, _11255_);
  and (_12547_, _12546_, _12543_);
  nor (_12548_, _06608_, \oc8051_golden_model_1.ACC [5]);
  and (_12549_, _06608_, \oc8051_golden_model_1.ACC [5]);
  nor (_12550_, _12549_, _12548_);
  not (_12551_, _12550_);
  nor (_12552_, _12551_, _11247_);
  nor (_12553_, _11241_, _10942_);
  and (_12554_, _12553_, _12552_);
  and (_12555_, _12554_, _12547_);
  or (_12556_, _12555_, _12362_);
  nand (_12557_, _12555_, _12356_);
  and (_12558_, _12557_, _06373_);
  and (_12559_, _12558_, _12556_);
  or (_12560_, _12559_, _12541_);
  and (_12561_, _12560_, _12246_);
  nand (_12562_, _12245_, _12102_);
  and (_12563_, _06664_, _06490_);
  not (_12564_, _12563_);
  not (_12565_, _07169_);
  nor (_12566_, _07174_, _06460_);
  and (_12567_, _12566_, _12565_);
  and (_12568_, _12567_, _12564_);
  not (_12569_, _07170_);
  nor (_12570_, _06461_, _07471_);
  and (_12571_, _12570_, _12569_);
  and (_12572_, _12571_, _07445_);
  and (_12573_, _12572_, _12568_);
  nand (_12574_, _12573_, _12562_);
  or (_12575_, _12574_, _12561_);
  or (_12576_, _12573_, _09443_);
  and (_12577_, _12576_, _12242_);
  and (_12578_, _12577_, _12575_);
  or (_12579_, _12578_, _12244_);
  and (_12580_, _06506_, _05958_);
  and (_12581_, _12580_, _12579_);
  not (_12582_, _12237_);
  not (_12583_, _12580_);
  and (_12584_, _12583_, _09443_);
  or (_12585_, _12584_, _12582_);
  or (_12586_, _12585_, _12581_);
  and (_12587_, _12586_, _12238_);
  nor (_12588_, _10542_, _06510_);
  not (_12589_, _12588_);
  or (_12590_, _12589_, _12587_);
  or (_12591_, _12588_, _09443_);
  and (_12592_, _12591_, _05977_);
  and (_12593_, _12592_, _12590_);
  and (_12594_, _12102_, _05976_);
  nor (_12595_, _06241_, _05970_);
  not (_12596_, _12595_);
  or (_12597_, _12596_, _12594_);
  or (_12598_, _12597_, _12593_);
  or (_12599_, _12595_, _09443_);
  and (_12600_, _12599_, _06370_);
  and (_12601_, _12600_, _12598_);
  and (_12602_, _09427_, _06369_);
  nor (_12603_, _07187_, _07182_);
  not (_12604_, _12603_);
  or (_12605_, _12604_, _12602_);
  or (_12606_, _12605_, _12601_);
  or (_12607_, _12603_, _09443_);
  and (_12608_, _12607_, _06336_);
  and (_12609_, _12608_, _12606_);
  or (_12610_, _12609_, _12235_);
  nor (_12611_, _10046_, _05935_);
  and (_12612_, _12611_, _12610_);
  nor (_12613_, _06332_, _05900_);
  not (_12614_, _12613_);
  not (_12615_, _12611_);
  and (_12616_, _12615_, _12102_);
  or (_12617_, _12616_, _12614_);
  or (_12618_, _12617_, _12612_);
  and (_12619_, _05899_, _06198_);
  not (_12620_, _12619_);
  or (_12621_, _12613_, _09443_);
  and (_12622_, _12621_, _12620_);
  and (_12623_, _12622_, _12618_);
  and (_12624_, _12619_, _12213_);
  or (_12625_, _12624_, _08973_);
  or (_12626_, _12625_, _12623_);
  and (_12627_, _12626_, _12234_);
  or (_12628_, _12627_, _06371_);
  or (_12629_, _09427_, _07198_);
  and (_12630_, _12629_, _10905_);
  and (_12631_, _12630_, _12628_);
  and (_12632_, _10904_, _09443_);
  or (_12633_, _12632_, _12631_);
  and (_12634_, _05934_, _05894_);
  not (_12635_, _12634_);
  and (_12636_, _12635_, _12633_);
  not (_12637_, \oc8051_golden_model_1.DPH [0]);
  and (_12638_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_12639_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_12640_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12641_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12642_, _12641_, _12640_);
  and (_12643_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12644_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12645_, _12644_, _12643_);
  not (_12646_, _12645_);
  and (_12647_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12648_, _06084_, _06080_);
  nor (_12649_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12650_, _12649_, _12647_);
  not (_12651_, _12650_);
  nor (_12652_, _12651_, _12648_);
  nor (_12653_, _12652_, _12647_);
  nor (_12654_, _12653_, _12646_);
  nor (_12655_, _12654_, _12643_);
  not (_12656_, _12655_);
  and (_12657_, _12656_, _12642_);
  nor (_12658_, _12657_, _12640_);
  nor (_12659_, _12658_, _12639_);
  nor (_12660_, _12659_, _12638_);
  nor (_12661_, _12660_, _12637_);
  and (_12662_, _12661_, \oc8051_golden_model_1.DPH [1]);
  and (_12663_, _12662_, \oc8051_golden_model_1.DPH [2]);
  and (_12665_, _12663_, \oc8051_golden_model_1.DPH [3]);
  and (_12666_, _12665_, \oc8051_golden_model_1.DPH [4]);
  and (_12667_, _12666_, \oc8051_golden_model_1.DPH [5]);
  and (_12668_, _12667_, \oc8051_golden_model_1.DPH [6]);
  nand (_12669_, _12668_, \oc8051_golden_model_1.DPH [7]);
  or (_12670_, _12668_, \oc8051_golden_model_1.DPH [7]);
  and (_12671_, _12670_, _12634_);
  and (_12672_, _12671_, _12669_);
  nor (_12673_, _06331_, _05895_);
  not (_12674_, _12673_);
  or (_12675_, _12674_, _12672_);
  or (_12676_, _12675_, _12636_);
  and (_12677_, _05894_, _06198_);
  not (_12678_, _12677_);
  or (_12679_, _12673_, _09443_);
  and (_12680_, _12679_, _12678_);
  and (_12681_, _12680_, _12676_);
  not (_12682_, _12232_);
  or (_12683_, _12213_, _11291_);
  not (_12684_, _11291_);
  or (_12686_, _12684_, _09443_);
  and (_12687_, _12686_, _12677_);
  and (_12688_, _12687_, _12683_);
  or (_12689_, _12688_, _12682_);
  or (_12690_, _12689_, _12681_);
  and (_12691_, _12690_, _12233_);
  or (_12692_, _12691_, _12229_);
  or (_12693_, _12228_, _09443_);
  and (_12694_, _12693_, _07218_);
  and (_12695_, _12694_, _12692_);
  and (_12696_, _09427_, _06367_);
  nor (_12697_, _06533_, _05889_);
  not (_12698_, _12697_);
  or (_12699_, _12698_, _12696_);
  or (_12700_, _12699_, _12695_);
  and (_12701_, _05888_, _06198_);
  not (_12702_, _12701_);
  or (_12703_, _12697_, _09443_);
  and (_12704_, _12703_, _12702_);
  and (_12705_, _12704_, _12700_);
  or (_12706_, _12213_, _12684_);
  or (_12707_, _11291_, _09443_);
  and (_12708_, _12707_, _12701_);
  and (_12709_, _12708_, _12706_);
  not (_12710_, _12226_);
  or (_12711_, _12710_, _12709_);
  or (_12712_, _12711_, _12705_);
  and (_12713_, _12712_, _12227_);
  or (_12714_, _12713_, _10968_);
  or (_12715_, _10967_, _09443_);
  and (_12716_, _12715_, _07213_);
  and (_12717_, _12716_, _12714_);
  and (_12718_, _09427_, _06366_);
  nor (_12719_, _06541_, _07209_);
  not (_12720_, _12719_);
  or (_12721_, _12720_, _12718_);
  or (_12722_, _12721_, _12717_);
  and (_12723_, _06365_, _06198_);
  not (_12724_, _12723_);
  or (_12725_, _12719_, _09443_);
  and (_12726_, _12725_, _12724_);
  and (_12727_, _12726_, _12722_);
  or (_12728_, _12213_, \oc8051_golden_model_1.PSW [7]);
  or (_12729_, _09443_, _10854_);
  and (_12730_, _12729_, _12723_);
  and (_12731_, _12730_, _12728_);
  or (_12732_, _12731_, _12727_);
  nor (_12733_, _07020_, _06654_);
  nor (_12734_, _07440_, _05921_);
  not (_12735_, _12734_);
  and (_12736_, _12735_, _12733_);
  and (_12737_, _12736_, _12732_);
  not (_12738_, _12736_);
  and (_12739_, _12738_, _12102_);
  or (_12740_, _12739_, _11006_);
  or (_12741_, _12740_, _12737_);
  or (_12742_, _11005_, _09443_);
  and (_12743_, _12742_, _07231_);
  and (_12744_, _12743_, _12741_);
  and (_12745_, _09427_, _06383_);
  not (_12746_, _05922_);
  nor (_12747_, _06528_, _12746_);
  not (_12748_, _12747_);
  or (_12749_, _12748_, _12745_);
  or (_12750_, _12749_, _12744_);
  not (_12751_, _12215_);
  or (_12752_, _12747_, _09443_);
  and (_12753_, _12752_, _12751_);
  and (_12754_, _12753_, _12750_);
  or (_12755_, _12754_, _12218_);
  and (_12756_, _10526_, _11022_);
  and (_12757_, _12756_, _12755_);
  not (_12758_, _12756_);
  and (_12759_, _12758_, _12102_);
  or (_12760_, _12759_, _11052_);
  or (_12761_, _12760_, _12757_);
  or (_12762_, _11051_, _09443_);
  and (_12763_, _12762_, _11081_);
  and (_12764_, _12763_, _12761_);
  and (_12765_, _12102_, _11080_);
  or (_12766_, _12765_, _06547_);
  or (_12767_, _12766_, _12764_);
  nand (_12768_, _08004_, _06547_);
  and (_12769_, _12768_, _12767_);
  or (_12770_, _12769_, _07228_);
  or (_12771_, _09443_, _05916_);
  and (_12772_, _12771_, _06946_);
  and (_12773_, _12772_, _12770_);
  not (_12774_, _12105_);
  not (_12775_, _07931_);
  and (_12776_, _08539_, \oc8051_golden_model_1.P3 [2]);
  and (_12777_, _08537_, \oc8051_golden_model_1.IE [2]);
  nor (_12778_, _12777_, _12776_);
  and (_12779_, _08533_, \oc8051_golden_model_1.SCON [2]);
  and (_12780_, _08535_, \oc8051_golden_model_1.P2 [2]);
  nor (_12781_, _12780_, _12779_);
  and (_12782_, _12781_, _12778_);
  and (_12783_, _08541_, \oc8051_golden_model_1.IP [2]);
  and (_12784_, _08543_, \oc8051_golden_model_1.PSW [2]);
  and (_12785_, _08545_, \oc8051_golden_model_1.ACC [2]);
  and (_12786_, _08547_, \oc8051_golden_model_1.B [2]);
  or (_12787_, _12786_, _12785_);
  or (_12788_, _12787_, _12784_);
  nor (_12789_, _12788_, _12783_);
  and (_12790_, _08528_, \oc8051_golden_model_1.TCON [2]);
  and (_12791_, _07920_, \oc8051_golden_model_1.P0 [2]);
  and (_12792_, _08531_, \oc8051_golden_model_1.P1 [2]);
  or (_12793_, _12792_, _12791_);
  nor (_12794_, _12793_, _12790_);
  and (_12795_, _12794_, _12789_);
  and (_12796_, _12795_, _12782_);
  and (_12797_, _12796_, _08395_);
  nor (_12798_, _12797_, _12775_);
  not (_12799_, _08134_);
  and (_12800_, _07920_, \oc8051_golden_model_1.P0 [1]);
  and (_12801_, _08528_, \oc8051_golden_model_1.TCON [1]);
  and (_12802_, _08531_, \oc8051_golden_model_1.P1 [1]);
  and (_12803_, _08533_, \oc8051_golden_model_1.SCON [1]);
  and (_12804_, _08535_, \oc8051_golden_model_1.P2 [1]);
  and (_12805_, _08537_, \oc8051_golden_model_1.IE [1]);
  and (_12806_, _08539_, \oc8051_golden_model_1.P3 [1]);
  and (_12807_, _08541_, \oc8051_golden_model_1.IP [1]);
  and (_12808_, _08543_, \oc8051_golden_model_1.PSW [1]);
  and (_12809_, _08545_, \oc8051_golden_model_1.ACC [1]);
  and (_12810_, _08547_, \oc8051_golden_model_1.B [1]);
  or (_12811_, _12810_, _12809_);
  or (_12812_, _12811_, _12808_);
  or (_12813_, _12812_, _12807_);
  or (_12814_, _12813_, _12806_);
  or (_12815_, _12814_, _12805_);
  or (_12816_, _12815_, _12804_);
  or (_12817_, _12816_, _12803_);
  or (_12818_, _12817_, _12802_);
  or (_12819_, _12818_, _12801_);
  nor (_12820_, _12819_, _12800_);
  and (_12821_, _12820_, _08300_);
  nor (_12822_, _12821_, _12799_);
  nor (_12823_, _12822_, _12798_);
  and (_12824_, _08533_, \oc8051_golden_model_1.SCON [4]);
  and (_12825_, _08539_, \oc8051_golden_model_1.P3 [4]);
  and (_12826_, _08537_, \oc8051_golden_model_1.IE [4]);
  or (_12827_, _12826_, _12825_);
  nor (_12828_, _12827_, _12824_);
  and (_12829_, _08528_, \oc8051_golden_model_1.TCON [4]);
  and (_12830_, _07920_, \oc8051_golden_model_1.P0 [4]);
  and (_12831_, _08531_, \oc8051_golden_model_1.P1 [4]);
  or (_12832_, _12831_, _12830_);
  nor (_12833_, _12832_, _12829_);
  and (_12834_, _08541_, \oc8051_golden_model_1.IP [4]);
  and (_12835_, _08547_, \oc8051_golden_model_1.B [4]);
  and (_12836_, _08545_, \oc8051_golden_model_1.ACC [4]);
  or (_12837_, _12836_, _12835_);
  nor (_12838_, _12837_, _12834_);
  and (_12839_, _08543_, \oc8051_golden_model_1.PSW [4]);
  and (_12840_, _08535_, \oc8051_golden_model_1.P2 [4]);
  nor (_12841_, _12840_, _12839_);
  and (_12842_, _12841_, _12838_);
  and (_12843_, _12842_, _12833_);
  and (_12844_, _12843_, _12828_);
  and (_12845_, _12844_, _08495_);
  and (_12846_, _07860_, _06751_);
  not (_12847_, _12846_);
  nor (_12848_, _12847_, _12845_);
  nor (_12849_, _12848_, _08705_);
  and (_12850_, _12849_, _12823_);
  and (_12851_, _07860_, _06750_);
  not (_12852_, _12851_);
  and (_12853_, _07920_, \oc8051_golden_model_1.P0 [0]);
  and (_12854_, _08528_, \oc8051_golden_model_1.TCON [0]);
  and (_12855_, _08531_, \oc8051_golden_model_1.P1 [0]);
  and (_12856_, _08533_, \oc8051_golden_model_1.SCON [0]);
  and (_12857_, _08535_, \oc8051_golden_model_1.P2 [0]);
  and (_12858_, _08537_, \oc8051_golden_model_1.IE [0]);
  and (_12859_, _08539_, \oc8051_golden_model_1.P3 [0]);
  and (_12860_, _08543_, \oc8051_golden_model_1.PSW [0]);
  and (_12861_, _08541_, \oc8051_golden_model_1.IP [0]);
  and (_12862_, _08547_, \oc8051_golden_model_1.B [0]);
  and (_12863_, _08545_, \oc8051_golden_model_1.ACC [0]);
  or (_12864_, _12863_, _12862_);
  or (_12865_, _12864_, _12861_);
  or (_12866_, _12865_, _12860_);
  or (_12867_, _12866_, _12859_);
  or (_12868_, _12867_, _12858_);
  or (_12869_, _12868_, _12857_);
  or (_12870_, _12869_, _12856_);
  or (_12871_, _12870_, _12855_);
  or (_12872_, _12871_, _12854_);
  nor (_12873_, _12872_, _12853_);
  not (_12874_, _12873_);
  nor (_12875_, _12874_, _08350_);
  nor (_12876_, _12875_, _12852_);
  and (_12877_, _08535_, \oc8051_golden_model_1.P2 [6]);
  and (_12878_, _08539_, \oc8051_golden_model_1.P3 [6]);
  and (_12879_, _08537_, \oc8051_golden_model_1.IE [6]);
  or (_12880_, _12879_, _12878_);
  nor (_12881_, _12880_, _12877_);
  and (_12882_, _08528_, \oc8051_golden_model_1.TCON [6]);
  and (_12883_, _08531_, \oc8051_golden_model_1.P1 [6]);
  and (_12884_, _07920_, \oc8051_golden_model_1.P0 [6]);
  or (_12885_, _12884_, _12883_);
  nor (_12886_, _12885_, _12882_);
  and (_12887_, _08541_, \oc8051_golden_model_1.IP [6]);
  and (_12888_, _08545_, \oc8051_golden_model_1.ACC [6]);
  and (_12889_, _08547_, \oc8051_golden_model_1.B [6]);
  or (_12890_, _12889_, _12888_);
  nor (_12891_, _12890_, _12887_);
  and (_12892_, _08533_, \oc8051_golden_model_1.SCON [6]);
  and (_12893_, _08543_, \oc8051_golden_model_1.PSW [6]);
  nor (_12894_, _12893_, _12892_);
  and (_12895_, _12894_, _12891_);
  and (_12896_, _12895_, _12886_);
  and (_12897_, _12896_, _12881_);
  and (_12898_, _12897_, _08107_);
  and (_12899_, _07891_, _06751_);
  not (_12900_, _12899_);
  nor (_12901_, _12900_, _12898_);
  nor (_12902_, _12901_, _12876_);
  not (_12903_, _08150_);
  and (_12904_, _07920_, \oc8051_golden_model_1.P0 [3]);
  and (_12905_, _08528_, \oc8051_golden_model_1.TCON [3]);
  and (_12906_, _08531_, \oc8051_golden_model_1.P1 [3]);
  and (_12907_, _08533_, \oc8051_golden_model_1.SCON [3]);
  and (_12908_, _08535_, \oc8051_golden_model_1.P2 [3]);
  and (_12909_, _08537_, \oc8051_golden_model_1.IE [3]);
  and (_12910_, _08539_, \oc8051_golden_model_1.P3 [3]);
  and (_12911_, _08541_, \oc8051_golden_model_1.IP [3]);
  and (_12912_, _08543_, \oc8051_golden_model_1.PSW [3]);
  and (_12913_, _08545_, \oc8051_golden_model_1.ACC [3]);
  and (_12914_, _08547_, \oc8051_golden_model_1.B [3]);
  or (_12915_, _12914_, _12913_);
  or (_12916_, _12915_, _12912_);
  or (_12917_, _12916_, _12911_);
  or (_12918_, _12917_, _12910_);
  or (_12919_, _12918_, _12909_);
  or (_12920_, _12919_, _12908_);
  or (_12921_, _12920_, _12907_);
  or (_12922_, _12921_, _12906_);
  or (_12923_, _12922_, _12905_);
  nor (_12924_, _12923_, _12904_);
  and (_12925_, _12924_, _08255_);
  nor (_12926_, _12925_, _12903_);
  and (_12927_, _08539_, \oc8051_golden_model_1.P3 [5]);
  and (_12928_, _08537_, \oc8051_golden_model_1.IE [5]);
  nor (_12929_, _12928_, _12927_);
  and (_12930_, _08533_, \oc8051_golden_model_1.SCON [5]);
  and (_12931_, _08535_, \oc8051_golden_model_1.P2 [5]);
  nor (_12932_, _12931_, _12930_);
  and (_12933_, _12932_, _12929_);
  and (_12934_, _08543_, \oc8051_golden_model_1.PSW [5]);
  and (_12935_, _08541_, \oc8051_golden_model_1.IP [5]);
  and (_12936_, _08545_, \oc8051_golden_model_1.ACC [5]);
  and (_12937_, _08547_, \oc8051_golden_model_1.B [5]);
  or (_12938_, _12937_, _12936_);
  or (_12939_, _12938_, _12935_);
  nor (_12940_, _12939_, _12934_);
  and (_12941_, _08528_, \oc8051_golden_model_1.TCON [5]);
  and (_12942_, _07920_, \oc8051_golden_model_1.P0 [5]);
  and (_12943_, _08531_, \oc8051_golden_model_1.P1 [5]);
  or (_12944_, _12943_, _12942_);
  nor (_12945_, _12944_, _12941_);
  and (_12946_, _12945_, _12940_);
  and (_12947_, _12946_, _12933_);
  and (_12948_, _12947_, _08210_);
  and (_12949_, _07851_, _06751_);
  not (_12950_, _12949_);
  nor (_12951_, _12950_, _12948_);
  nor (_12952_, _12951_, _12926_);
  and (_12953_, _12952_, _12902_);
  and (_12954_, _12953_, _12850_);
  not (_12955_, _12954_);
  or (_12956_, _12362_, _12955_);
  or (_12957_, _09427_, _12954_);
  and (_12958_, _12957_, _06381_);
  and (_12959_, _12958_, _12956_);
  or (_12960_, _12959_, _12774_);
  or (_12961_, _12960_, _12773_);
  and (_12962_, _12961_, _12106_);
  nor (_12963_, _10450_, _06293_);
  not (_12964_, _12963_);
  or (_12965_, _12964_, _12962_);
  not (_12966_, _10448_);
  or (_12967_, _12963_, _09443_);
  and (_12968_, _12967_, _12966_);
  and (_12969_, _12968_, _12965_);
  and (_12970_, _12102_, _10448_);
  or (_12971_, _12970_, _06260_);
  or (_12972_, _12971_, _12969_);
  nand (_12973_, _08004_, _06260_);
  and (_12974_, _12973_, _12972_);
  or (_12975_, _12974_, _12089_);
  or (_12976_, _09443_, _05924_);
  and (_12977_, _12976_, _06564_);
  and (_12978_, _12977_, _12975_);
  or (_12979_, _12362_, _12954_);
  nand (_12980_, _12356_, _12954_);
  and (_12981_, _12980_, _12979_);
  and (_12982_, _12981_, _06377_);
  and (_12983_, _09012_, _07463_);
  and (_12984_, _12983_, _07403_);
  not (_12985_, _12984_);
  or (_12986_, _12985_, _12982_);
  or (_12987_, _12986_, _12978_);
  or (_12988_, _12984_, _12102_);
  and (_12989_, _12988_, _07241_);
  and (_12990_, _12989_, _12987_);
  nor (_12991_, _11284_, _11279_);
  not (_12992_, _12991_);
  and (_12993_, _09443_, _06563_);
  or (_12994_, _12993_, _12992_);
  or (_12995_, _12994_, _12990_);
  or (_12996_, _12102_, _12991_);
  and (_12997_, _12996_, _08505_);
  and (_12998_, _12997_, _12995_);
  and (_12999_, _06378_, _06187_);
  or (_13000_, _12999_, _05912_);
  or (_13001_, _13000_, _12998_);
  or (_13002_, _09443_, _05913_);
  and (_13003_, _13002_, _06571_);
  and (_13004_, _13003_, _13001_);
  and (_13005_, _12981_, _06199_);
  and (_13006_, _09371_, _07414_);
  not (_13007_, _13006_);
  or (_13008_, _13007_, _13005_);
  or (_13009_, _13008_, _13004_);
  or (_13010_, _13006_, _12102_);
  and (_13011_, _13010_, _06189_);
  and (_13012_, _13011_, _13009_);
  nor (_13013_, _11309_, _11302_);
  not (_13014_, _13013_);
  and (_13015_, _09443_, _06188_);
  or (_13016_, _13015_, _13014_);
  or (_13017_, _13016_, _13012_);
  not (_13018_, _06342_);
  or (_13019_, _12102_, _13013_);
  and (_13020_, _13019_, _13018_);
  and (_13021_, _13020_, _13017_);
  and (_13022_, _06342_, _06187_);
  or (_13023_, _13022_, _05907_);
  or (_13024_, _13023_, _13021_);
  and (_13025_, _06198_, _05906_);
  not (_13026_, _13025_);
  or (_13027_, _09443_, _05908_);
  and (_13028_, _13027_, _13026_);
  and (_13029_, _13028_, _13024_);
  and (_13030_, _13025_, _12102_);
  or (_13031_, _13030_, _13029_);
  or (_13032_, _13031_, _01456_);
  or (_13033_, _01452_, \oc8051_golden_model_1.PC [15]);
  and (_13034_, _13033_, _43223_);
  and (_41192_, _13034_, _13032_);
  not (_13035_, _07881_);
  and (_13036_, _13035_, \oc8051_golden_model_1.P2 [7]);
  and (_13037_, _08509_, _07881_);
  or (_13038_, _13037_, _13036_);
  and (_13039_, _13038_, _06533_);
  nor (_13040_, _08004_, _13035_);
  or (_13041_, _13040_, _13036_);
  or (_13042_, _13041_, _07188_);
  not (_13043_, _08535_);
  and (_13044_, _13043_, \oc8051_golden_model_1.P2 [7]);
  and (_13045_, _08698_, _08535_);
  or (_13046_, _13045_, _13044_);
  and (_13047_, _13046_, _06483_);
  or (_13048_, _13041_, _07142_);
  and (_13049_, _08685_, _07881_);
  or (_13050_, _13049_, _13036_);
  or (_13051_, _13050_, _06252_);
  and (_13052_, _07881_, \oc8051_golden_model_1.ACC [7]);
  or (_13053_, _13052_, _13036_);
  and (_13054_, _13053_, _07123_);
  and (_13055_, _07124_, \oc8051_golden_model_1.P2 [7]);
  or (_13056_, _13055_, _06251_);
  or (_13057_, _13056_, _13054_);
  and (_13058_, _13057_, _06476_);
  and (_13059_, _13058_, _13051_);
  and (_13060_, _08560_, _08535_);
  or (_13061_, _13060_, _13044_);
  and (_13062_, _13061_, _06475_);
  or (_13063_, _13062_, _06468_);
  or (_13064_, _13063_, _13059_);
  and (_13065_, _13064_, _13048_);
  or (_13066_, _13065_, _06466_);
  or (_13067_, _13053_, _06801_);
  and (_13068_, _13067_, _06484_);
  and (_13069_, _13068_, _13066_);
  or (_13070_, _13069_, _13047_);
  and (_13071_, _13070_, _07164_);
  or (_13072_, _13044_, _08706_);
  and (_13073_, _13072_, _06461_);
  and (_13074_, _13073_, _13061_);
  or (_13075_, _13074_, _13071_);
  and (_13076_, _13075_, _06242_);
  and (_13077_, _08726_, _08535_);
  or (_13078_, _13077_, _13044_);
  and (_13079_, _13078_, _06241_);
  or (_13080_, _13079_, _07187_);
  or (_13081_, _13080_, _13076_);
  and (_13082_, _13081_, _13042_);
  or (_13083_, _13082_, _07182_);
  and (_13084_, _08671_, _07881_);
  or (_13085_, _13036_, _07183_);
  or (_13086_, _13085_, _13084_);
  and (_13087_, _13086_, _06336_);
  and (_13088_, _13087_, _13083_);
  and (_13089_, _08966_, _07881_);
  or (_13090_, _13089_, _13036_);
  and (_13091_, _13090_, _05968_);
  or (_13092_, _13091_, _06371_);
  or (_13093_, _13092_, _13088_);
  and (_13094_, _08770_, _07881_);
  or (_13095_, _13094_, _13036_);
  or (_13096_, _13095_, _07198_);
  and (_13097_, _13096_, _13093_);
  or (_13098_, _13097_, _06367_);
  and (_13099_, _08988_, _07881_);
  or (_13100_, _13099_, _13036_);
  or (_13101_, _13100_, _07218_);
  and (_13102_, _13101_, _07216_);
  and (_13103_, _13102_, _13098_);
  or (_13104_, _13103_, _13039_);
  and (_13105_, _13104_, _07213_);
  or (_13106_, _13036_, _08007_);
  and (_13107_, _13095_, _06366_);
  and (_13108_, _13107_, _13106_);
  or (_13109_, _13108_, _13105_);
  and (_13110_, _13109_, _07210_);
  and (_13111_, _13053_, _06541_);
  and (_13112_, _13111_, _13106_);
  or (_13113_, _13112_, _06383_);
  or (_13114_, _13113_, _13110_);
  and (_13115_, _08985_, _07881_);
  or (_13116_, _13036_, _07231_);
  or (_13117_, _13116_, _13115_);
  and (_13118_, _13117_, _07229_);
  and (_13119_, _13118_, _13114_);
  nor (_13120_, _08508_, _13035_);
  or (_13121_, _13120_, _13036_);
  and (_13122_, _13121_, _06528_);
  or (_13123_, _13122_, _06563_);
  or (_13124_, _13123_, _13119_);
  or (_13125_, _13050_, _07241_);
  and (_13126_, _13125_, _06571_);
  and (_13127_, _13126_, _13124_);
  and (_13128_, _13046_, _06199_);
  or (_13129_, _13128_, _06188_);
  or (_13130_, _13129_, _13127_);
  and (_13131_, _08503_, _07881_);
  or (_13132_, _13036_, _06189_);
  or (_13133_, _13132_, _13131_);
  and (_13134_, _13133_, _01452_);
  and (_13135_, _13134_, _13130_);
  nor (_13136_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_13137_, _13136_, _00000_);
  or (_41193_, _13137_, _13135_);
  not (_13138_, _07871_);
  and (_13139_, _13138_, \oc8051_golden_model_1.P3 [7]);
  and (_13140_, _08509_, _07871_);
  or (_13141_, _13140_, _13139_);
  and (_13142_, _13141_, _06533_);
  nor (_13143_, _08004_, _13138_);
  or (_13144_, _13143_, _13139_);
  or (_13145_, _13144_, _07188_);
  not (_13146_, _08539_);
  and (_13147_, _13146_, \oc8051_golden_model_1.P3 [7]);
  and (_13148_, _08698_, _08539_);
  or (_13149_, _13148_, _13147_);
  and (_13150_, _13149_, _06483_);
  or (_13151_, _13144_, _07142_);
  and (_13152_, _08685_, _07871_);
  or (_13153_, _13152_, _13139_);
  or (_13154_, _13153_, _06252_);
  and (_13155_, _07871_, \oc8051_golden_model_1.ACC [7]);
  or (_13156_, _13155_, _13139_);
  and (_13157_, _13156_, _07123_);
  and (_13158_, _07124_, \oc8051_golden_model_1.P3 [7]);
  or (_13159_, _13158_, _06251_);
  or (_13160_, _13159_, _13157_);
  and (_13161_, _13160_, _06476_);
  and (_13162_, _13161_, _13154_);
  and (_13163_, _08560_, _08539_);
  or (_13164_, _13163_, _13147_);
  and (_13165_, _13164_, _06475_);
  or (_13166_, _13165_, _06468_);
  or (_13167_, _13166_, _13162_);
  and (_13168_, _13167_, _13151_);
  or (_13169_, _13168_, _06466_);
  or (_13170_, _13156_, _06801_);
  and (_13171_, _13170_, _06484_);
  and (_13172_, _13171_, _13169_);
  or (_13173_, _13172_, _13150_);
  and (_13174_, _13173_, _07164_);
  and (_13175_, _08707_, _08539_);
  or (_13176_, _13175_, _13147_);
  and (_13177_, _13176_, _06461_);
  or (_13178_, _13177_, _13174_);
  and (_13179_, _13178_, _06242_);
  and (_13180_, _08726_, _08539_);
  or (_13181_, _13180_, _13147_);
  and (_13182_, _13181_, _06241_);
  or (_13183_, _13182_, _07187_);
  or (_13184_, _13183_, _13179_);
  and (_13185_, _13184_, _13145_);
  or (_13186_, _13185_, _07182_);
  and (_13187_, _08671_, _07871_);
  or (_13188_, _13139_, _07183_);
  or (_13189_, _13188_, _13187_);
  and (_13190_, _13189_, _06336_);
  and (_13191_, _13190_, _13186_);
  and (_13192_, _08966_, _07871_);
  or (_13193_, _13192_, _13139_);
  and (_13194_, _13193_, _05968_);
  or (_13195_, _13194_, _06371_);
  or (_13196_, _13195_, _13191_);
  and (_13197_, _08770_, _07871_);
  or (_13198_, _13197_, _13139_);
  or (_13199_, _13198_, _07198_);
  and (_13200_, _13199_, _13196_);
  or (_13201_, _13200_, _06367_);
  and (_13202_, _08988_, _07871_);
  or (_13203_, _13202_, _13139_);
  or (_13204_, _13203_, _07218_);
  and (_13205_, _13204_, _07216_);
  and (_13206_, _13205_, _13201_);
  or (_13207_, _13206_, _13142_);
  and (_13208_, _13207_, _07213_);
  or (_13209_, _13139_, _08007_);
  and (_13210_, _13198_, _06366_);
  and (_13211_, _13210_, _13209_);
  or (_13212_, _13211_, _13208_);
  and (_13213_, _13212_, _07210_);
  and (_13214_, _13156_, _06541_);
  and (_13215_, _13214_, _13209_);
  or (_13216_, _13215_, _06383_);
  or (_13217_, _13216_, _13213_);
  and (_13218_, _08985_, _07871_);
  or (_13219_, _13139_, _07231_);
  or (_13220_, _13219_, _13218_);
  and (_13221_, _13220_, _07229_);
  and (_13222_, _13221_, _13217_);
  nor (_13223_, _08508_, _13138_);
  or (_13224_, _13223_, _13139_);
  and (_13225_, _13224_, _06528_);
  or (_13226_, _13225_, _06563_);
  or (_13227_, _13226_, _13222_);
  or (_13228_, _13153_, _07241_);
  and (_13229_, _13228_, _06571_);
  and (_13230_, _13229_, _13227_);
  and (_13231_, _13149_, _06199_);
  or (_13232_, _13231_, _06188_);
  or (_13233_, _13232_, _13230_);
  and (_13234_, _08503_, _07871_);
  or (_13235_, _13139_, _06189_);
  or (_13236_, _13235_, _13234_);
  and (_13237_, _13236_, _01452_);
  and (_13238_, _13237_, _13233_);
  nor (_13239_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_13240_, _13239_, _00000_);
  or (_41194_, _13240_, _13238_);
  not (_13241_, _07899_);
  and (_13242_, _13241_, \oc8051_golden_model_1.P0 [7]);
  and (_13243_, _08509_, _07899_);
  or (_13244_, _13243_, _13242_);
  and (_13245_, _13244_, _06533_);
  nor (_13246_, _08004_, _13241_);
  or (_13247_, _13246_, _13242_);
  or (_13248_, _13247_, _07188_);
  or (_13249_, _13247_, _07142_);
  and (_13250_, _08685_, _07899_);
  or (_13251_, _13250_, _13242_);
  or (_13252_, _13251_, _06252_);
  and (_13253_, _07899_, \oc8051_golden_model_1.ACC [7]);
  or (_13254_, _13253_, _13242_);
  and (_13255_, _13254_, _07123_);
  and (_13256_, _07124_, \oc8051_golden_model_1.P0 [7]);
  or (_13257_, _13256_, _06251_);
  or (_13258_, _13257_, _13255_);
  and (_13259_, _13258_, _06476_);
  and (_13260_, _13259_, _13252_);
  not (_13261_, _07920_);
  and (_13262_, _13261_, \oc8051_golden_model_1.P0 [7]);
  and (_13263_, _08560_, _07920_);
  or (_13264_, _13263_, _13262_);
  and (_13265_, _13264_, _06475_);
  or (_13266_, _13265_, _06468_);
  or (_13267_, _13266_, _13260_);
  and (_13268_, _13267_, _13249_);
  or (_13269_, _13268_, _06466_);
  or (_13270_, _13254_, _06801_);
  and (_13271_, _13270_, _06484_);
  and (_13272_, _13271_, _13269_);
  and (_13273_, _08698_, _07920_);
  or (_13274_, _13273_, _13262_);
  and (_13275_, _13274_, _06483_);
  or (_13276_, _13275_, _13272_);
  and (_13277_, _13276_, _07164_);
  and (_13278_, _08707_, _07920_);
  or (_13279_, _13278_, _13262_);
  and (_13280_, _13279_, _06461_);
  or (_13281_, _13280_, _13277_);
  and (_13282_, _13281_, _06242_);
  and (_13283_, _08726_, _07920_);
  or (_13284_, _13283_, _13262_);
  and (_13285_, _13284_, _06241_);
  or (_13286_, _13285_, _07187_);
  or (_13287_, _13286_, _13282_);
  and (_13288_, _13287_, _13248_);
  or (_13289_, _13288_, _07182_);
  and (_13290_, _08671_, _07899_);
  or (_13291_, _13242_, _07183_);
  or (_13292_, _13291_, _13290_);
  and (_13293_, _13292_, _06336_);
  and (_13294_, _13293_, _13289_);
  and (_13295_, _08966_, _07899_);
  or (_13296_, _13295_, _13242_);
  and (_13297_, _13296_, _05968_);
  or (_13298_, _13297_, _06371_);
  or (_13299_, _13298_, _13294_);
  and (_13300_, _08770_, _07899_);
  or (_13301_, _13300_, _13242_);
  or (_13302_, _13301_, _07198_);
  and (_13303_, _13302_, _13299_);
  or (_13304_, _13303_, _06367_);
  and (_13305_, _08988_, _07899_);
  or (_13306_, _13305_, _13242_);
  or (_13307_, _13306_, _07218_);
  and (_13308_, _13307_, _07216_);
  and (_13309_, _13308_, _13304_);
  or (_13310_, _13309_, _13245_);
  and (_13311_, _13310_, _07213_);
  or (_13312_, _13242_, _08007_);
  and (_13313_, _13301_, _06366_);
  and (_13314_, _13313_, _13312_);
  or (_13315_, _13314_, _13311_);
  and (_13316_, _13315_, _07210_);
  and (_13317_, _13254_, _06541_);
  and (_13318_, _13317_, _13312_);
  or (_13319_, _13318_, _06383_);
  or (_13320_, _13319_, _13316_);
  and (_13321_, _08985_, _07899_);
  or (_13322_, _13242_, _07231_);
  or (_13323_, _13322_, _13321_);
  and (_13324_, _13323_, _07229_);
  and (_13325_, _13324_, _13320_);
  nor (_13326_, _08508_, _13241_);
  or (_13327_, _13326_, _13242_);
  and (_13328_, _13327_, _06528_);
  or (_13329_, _13328_, _06563_);
  or (_13330_, _13329_, _13325_);
  or (_13331_, _13251_, _07241_);
  and (_13332_, _13331_, _06571_);
  and (_13333_, _13332_, _13330_);
  and (_13334_, _13274_, _06199_);
  or (_13335_, _13334_, _06188_);
  or (_13336_, _13335_, _13333_);
  and (_13337_, _08503_, _07899_);
  or (_13338_, _13242_, _06189_);
  or (_13339_, _13338_, _13337_);
  and (_13340_, _13339_, _01452_);
  and (_13341_, _13340_, _13336_);
  nor (_13342_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_13343_, _13342_, _00000_);
  or (_41195_, _13343_, _13341_);
  nor (_13344_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_13345_, _13344_, _00000_);
  not (_13346_, _07945_);
  and (_13347_, _13346_, \oc8051_golden_model_1.P1 [7]);
  and (_13348_, _08509_, _07945_);
  or (_13349_, _13348_, _13347_);
  and (_13350_, _13349_, _06533_);
  nor (_13351_, _08004_, _13346_);
  or (_13352_, _13351_, _13347_);
  or (_13353_, _13352_, _07188_);
  or (_13354_, _13352_, _07142_);
  and (_13355_, _08685_, _07945_);
  or (_13356_, _13355_, _13347_);
  or (_13357_, _13356_, _06252_);
  and (_13358_, _07945_, \oc8051_golden_model_1.ACC [7]);
  or (_13359_, _13358_, _13347_);
  and (_13360_, _13359_, _07123_);
  and (_13361_, _07124_, \oc8051_golden_model_1.P1 [7]);
  or (_13362_, _13361_, _06251_);
  or (_13363_, _13362_, _13360_);
  and (_13364_, _13363_, _06476_);
  and (_13365_, _13364_, _13357_);
  not (_13366_, _08531_);
  and (_13367_, _13366_, \oc8051_golden_model_1.P1 [7]);
  and (_13368_, _08560_, _08531_);
  or (_13369_, _13368_, _13367_);
  and (_13370_, _13369_, _06475_);
  or (_13371_, _13370_, _06468_);
  or (_13372_, _13371_, _13365_);
  and (_13373_, _13372_, _13354_);
  or (_13374_, _13373_, _06466_);
  or (_13375_, _13359_, _06801_);
  and (_13376_, _13375_, _06484_);
  and (_13377_, _13376_, _13374_);
  and (_13378_, _08698_, _08531_);
  or (_13379_, _13378_, _13367_);
  and (_13380_, _13379_, _06483_);
  or (_13381_, _13380_, _13377_);
  and (_13382_, _13381_, _07164_);
  or (_13383_, _13367_, _08706_);
  and (_13384_, _13383_, _06461_);
  and (_13385_, _13384_, _13369_);
  or (_13386_, _13385_, _13382_);
  and (_13387_, _13386_, _06242_);
  and (_13388_, _08726_, _08531_);
  or (_13389_, _13388_, _13367_);
  and (_13390_, _13389_, _06241_);
  or (_13391_, _13390_, _07187_);
  or (_13392_, _13391_, _13387_);
  and (_13393_, _13392_, _13353_);
  or (_13394_, _13393_, _07182_);
  and (_13395_, _08671_, _07945_);
  or (_13396_, _13347_, _07183_);
  or (_13397_, _13396_, _13395_);
  and (_13398_, _13397_, _06336_);
  and (_13399_, _13398_, _13394_);
  and (_13400_, _08966_, _07945_);
  or (_13401_, _13400_, _13347_);
  and (_13402_, _13401_, _05968_);
  or (_13403_, _13402_, _06371_);
  or (_13404_, _13403_, _13399_);
  and (_13405_, _08770_, _07945_);
  or (_13406_, _13405_, _13347_);
  or (_13407_, _13406_, _07198_);
  and (_13408_, _13407_, _13404_);
  or (_13409_, _13408_, _06367_);
  and (_13410_, _08988_, _07945_);
  or (_13411_, _13410_, _13347_);
  or (_13412_, _13411_, _07218_);
  and (_13413_, _13412_, _07216_);
  and (_13414_, _13413_, _13409_);
  or (_13415_, _13414_, _13350_);
  and (_13416_, _13415_, _07213_);
  or (_13417_, _13347_, _08007_);
  and (_13418_, _13406_, _06366_);
  and (_13419_, _13418_, _13417_);
  or (_13420_, _13419_, _13416_);
  and (_13421_, _13420_, _07210_);
  and (_13422_, _13359_, _06541_);
  and (_13423_, _13422_, _13417_);
  or (_13424_, _13423_, _06383_);
  or (_13425_, _13424_, _13421_);
  and (_13426_, _08985_, _07945_);
  or (_13427_, _13347_, _07231_);
  or (_13428_, _13427_, _13426_);
  and (_13429_, _13428_, _07229_);
  and (_13430_, _13429_, _13425_);
  nor (_13431_, _08508_, _13346_);
  or (_13432_, _13431_, _13347_);
  and (_13433_, _13432_, _06528_);
  or (_13434_, _13433_, _06563_);
  or (_13435_, _13434_, _13430_);
  or (_13436_, _13356_, _07241_);
  and (_13437_, _13436_, _06571_);
  and (_13438_, _13437_, _13435_);
  and (_13439_, _13379_, _06199_);
  or (_13440_, _13439_, _06188_);
  or (_13441_, _13440_, _13438_);
  and (_13442_, _08503_, _07945_);
  or (_13443_, _13347_, _06189_);
  or (_13444_, _13443_, _13442_);
  and (_13445_, _13444_, _01452_);
  and (_13446_, _13445_, _13441_);
  or (_41197_, _13446_, _13345_);
  and (_13447_, _01456_, \oc8051_golden_model_1.IP [7]);
  not (_13448_, _07918_);
  and (_13449_, _13448_, \oc8051_golden_model_1.IP [7]);
  and (_13450_, _08509_, _07918_);
  or (_13451_, _13450_, _13449_);
  and (_13452_, _13451_, _06533_);
  nor (_13453_, _08004_, _13448_);
  or (_13454_, _13453_, _13449_);
  or (_13455_, _13454_, _07188_);
  or (_13456_, _13454_, _07142_);
  and (_13457_, _08685_, _07918_);
  or (_13458_, _13457_, _13449_);
  or (_13459_, _13458_, _06252_);
  and (_13460_, _07918_, \oc8051_golden_model_1.ACC [7]);
  or (_13461_, _13460_, _13449_);
  and (_13462_, _13461_, _07123_);
  and (_13463_, _07124_, \oc8051_golden_model_1.IP [7]);
  or (_13464_, _13463_, _06251_);
  or (_13465_, _13464_, _13462_);
  and (_13466_, _13465_, _06476_);
  and (_13467_, _13466_, _13459_);
  not (_13468_, _08541_);
  and (_13469_, _13468_, \oc8051_golden_model_1.IP [7]);
  and (_13470_, _08560_, _08541_);
  or (_13471_, _13470_, _13469_);
  and (_13472_, _13471_, _06475_);
  or (_13473_, _13472_, _06468_);
  or (_13474_, _13473_, _13467_);
  and (_13475_, _13474_, _13456_);
  or (_13476_, _13475_, _06466_);
  or (_13477_, _13461_, _06801_);
  and (_13478_, _13477_, _06484_);
  and (_13479_, _13478_, _13476_);
  and (_13480_, _08698_, _08541_);
  or (_13481_, _13480_, _13469_);
  and (_13482_, _13481_, _06483_);
  or (_13483_, _13482_, _13479_);
  and (_13484_, _13483_, _07164_);
  and (_13485_, _08707_, _08541_);
  or (_13486_, _13485_, _13469_);
  and (_13487_, _13486_, _06461_);
  or (_13488_, _13487_, _13484_);
  and (_13489_, _13488_, _06242_);
  and (_13490_, _08726_, _08541_);
  or (_13491_, _13490_, _13469_);
  and (_13492_, _13491_, _06241_);
  or (_13493_, _13492_, _07187_);
  or (_13494_, _13493_, _13489_);
  and (_13495_, _13494_, _13455_);
  or (_13496_, _13495_, _07182_);
  and (_13497_, _08671_, _07918_);
  or (_13498_, _13449_, _07183_);
  or (_13499_, _13498_, _13497_);
  and (_13500_, _13499_, _06336_);
  and (_13501_, _13500_, _13496_);
  and (_13502_, _08966_, _07918_);
  or (_13503_, _13502_, _13449_);
  and (_13504_, _13503_, _05968_);
  or (_13505_, _13504_, _06371_);
  or (_13506_, _13505_, _13501_);
  and (_13507_, _08770_, _07918_);
  or (_13508_, _13507_, _13449_);
  or (_13509_, _13508_, _07198_);
  and (_13510_, _13509_, _13506_);
  or (_13511_, _13510_, _06367_);
  and (_13512_, _08988_, _07918_);
  or (_13513_, _13512_, _13449_);
  or (_13514_, _13513_, _07218_);
  and (_13515_, _13514_, _07216_);
  and (_13516_, _13515_, _13511_);
  or (_13517_, _13516_, _13452_);
  and (_13518_, _13517_, _07213_);
  or (_13519_, _13449_, _08007_);
  and (_13520_, _13508_, _06366_);
  and (_13521_, _13520_, _13519_);
  or (_13522_, _13521_, _13518_);
  and (_13523_, _13522_, _07210_);
  and (_13524_, _13461_, _06541_);
  and (_13525_, _13524_, _13519_);
  or (_13526_, _13525_, _06383_);
  or (_13527_, _13526_, _13523_);
  and (_13528_, _08985_, _07918_);
  or (_13529_, _13449_, _07231_);
  or (_13530_, _13529_, _13528_);
  and (_13531_, _13530_, _07229_);
  and (_13532_, _13531_, _13527_);
  nor (_13533_, _08508_, _13448_);
  or (_13534_, _13533_, _13449_);
  and (_13535_, _13534_, _06528_);
  or (_13536_, _13535_, _06563_);
  or (_13537_, _13536_, _13532_);
  or (_13538_, _13458_, _07241_);
  and (_13539_, _13538_, _06571_);
  and (_13540_, _13539_, _13537_);
  and (_13541_, _13481_, _06199_);
  or (_13542_, _13541_, _06188_);
  or (_13543_, _13542_, _13540_);
  and (_13544_, _08503_, _07918_);
  or (_13545_, _13449_, _06189_);
  or (_13546_, _13545_, _13544_);
  and (_13547_, _13546_, _01452_);
  and (_13548_, _13547_, _13543_);
  or (_13549_, _13548_, _13447_);
  and (_41198_, _13549_, _43223_);
  and (_13550_, _01456_, \oc8051_golden_model_1.IE [7]);
  not (_13551_, _07865_);
  and (_13552_, _13551_, \oc8051_golden_model_1.IE [7]);
  and (_13553_, _08509_, _07865_);
  or (_13554_, _13553_, _13552_);
  and (_13555_, _13554_, _06533_);
  nor (_13556_, _08004_, _13551_);
  or (_13557_, _13556_, _13552_);
  or (_13558_, _13557_, _07188_);
  or (_13559_, _13557_, _07142_);
  and (_13560_, _08685_, _07865_);
  or (_13561_, _13560_, _13552_);
  or (_13562_, _13561_, _06252_);
  and (_13563_, _07865_, \oc8051_golden_model_1.ACC [7]);
  or (_13564_, _13563_, _13552_);
  and (_13565_, _13564_, _07123_);
  and (_13566_, _07124_, \oc8051_golden_model_1.IE [7]);
  or (_13567_, _13566_, _06251_);
  or (_13568_, _13567_, _13565_);
  and (_13569_, _13568_, _06476_);
  and (_13570_, _13569_, _13562_);
  not (_13571_, _08537_);
  and (_13572_, _13571_, \oc8051_golden_model_1.IE [7]);
  and (_13573_, _08560_, _08537_);
  or (_13574_, _13573_, _13572_);
  and (_13575_, _13574_, _06475_);
  or (_13576_, _13575_, _06468_);
  or (_13577_, _13576_, _13570_);
  and (_13578_, _13577_, _13559_);
  or (_13579_, _13578_, _06466_);
  or (_13580_, _13564_, _06801_);
  and (_13581_, _13580_, _06484_);
  and (_13582_, _13581_, _13579_);
  and (_13583_, _08698_, _08537_);
  or (_13584_, _13583_, _13572_);
  and (_13585_, _13584_, _06483_);
  or (_13586_, _13585_, _13582_);
  and (_13587_, _13586_, _07164_);
  and (_13588_, _08707_, _08537_);
  or (_13589_, _13588_, _13572_);
  and (_13590_, _13589_, _06461_);
  or (_13591_, _13590_, _13587_);
  and (_13592_, _13591_, _06242_);
  and (_13593_, _08726_, _08537_);
  or (_13594_, _13593_, _13572_);
  and (_13595_, _13594_, _06241_);
  or (_13596_, _13595_, _07187_);
  or (_13597_, _13596_, _13592_);
  and (_13598_, _13597_, _13558_);
  or (_13599_, _13598_, _07182_);
  and (_13601_, _08671_, _07865_);
  or (_13602_, _13552_, _07183_);
  or (_13603_, _13602_, _13601_);
  and (_13604_, _13603_, _06336_);
  and (_13605_, _13604_, _13599_);
  and (_13606_, _08966_, _07865_);
  or (_13607_, _13606_, _13552_);
  and (_13608_, _13607_, _05968_);
  or (_13609_, _13608_, _06371_);
  or (_13610_, _13609_, _13605_);
  and (_13612_, _08770_, _07865_);
  or (_13613_, _13612_, _13552_);
  or (_13614_, _13613_, _07198_);
  and (_13615_, _13614_, _13610_);
  or (_13616_, _13615_, _06367_);
  and (_13617_, _08988_, _07865_);
  or (_13618_, _13617_, _13552_);
  or (_13619_, _13618_, _07218_);
  and (_13620_, _13619_, _07216_);
  and (_13621_, _13620_, _13616_);
  or (_13623_, _13621_, _13555_);
  and (_13624_, _13623_, _07213_);
  or (_13625_, _13552_, _08007_);
  and (_13626_, _13613_, _06366_);
  and (_13627_, _13626_, _13625_);
  or (_13628_, _13627_, _13624_);
  and (_13629_, _13628_, _07210_);
  and (_13630_, _13564_, _06541_);
  and (_13631_, _13630_, _13625_);
  or (_13632_, _13631_, _06383_);
  or (_13634_, _13632_, _13629_);
  and (_13635_, _08985_, _07865_);
  or (_13636_, _13552_, _07231_);
  or (_13637_, _13636_, _13635_);
  and (_13638_, _13637_, _07229_);
  and (_13639_, _13638_, _13634_);
  nor (_13640_, _08508_, _13551_);
  or (_13641_, _13640_, _13552_);
  and (_13642_, _13641_, _06528_);
  or (_13643_, _13642_, _06563_);
  or (_13645_, _13643_, _13639_);
  or (_13646_, _13561_, _07241_);
  and (_13647_, _13646_, _06571_);
  and (_13648_, _13647_, _13645_);
  and (_13649_, _13584_, _06199_);
  or (_13650_, _13649_, _06188_);
  or (_13651_, _13650_, _13648_);
  and (_13652_, _08503_, _07865_);
  or (_13653_, _13552_, _06189_);
  or (_13654_, _13653_, _13652_);
  and (_13656_, _13654_, _01452_);
  and (_13657_, _13656_, _13651_);
  or (_13658_, _13657_, _13550_);
  and (_41199_, _13658_, _43223_);
  and (_13659_, _01456_, \oc8051_golden_model_1.SCON [7]);
  not (_13660_, _07943_);
  and (_13661_, _13660_, \oc8051_golden_model_1.SCON [7]);
  and (_13662_, _08509_, _07943_);
  or (_13663_, _13662_, _13661_);
  and (_13664_, _13663_, _06533_);
  nor (_13666_, _08004_, _13660_);
  or (_13667_, _13666_, _13661_);
  or (_13668_, _13667_, _07188_);
  or (_13669_, _13667_, _07142_);
  and (_13670_, _08685_, _07943_);
  or (_13671_, _13670_, _13661_);
  or (_13672_, _13671_, _06252_);
  and (_13673_, _07943_, \oc8051_golden_model_1.ACC [7]);
  or (_13674_, _13673_, _13661_);
  and (_13675_, _13674_, _07123_);
  and (_13677_, _07124_, \oc8051_golden_model_1.SCON [7]);
  or (_13678_, _13677_, _06251_);
  or (_13679_, _13678_, _13675_);
  and (_13680_, _13679_, _06476_);
  and (_13681_, _13680_, _13672_);
  not (_13682_, _08533_);
  and (_13683_, _13682_, \oc8051_golden_model_1.SCON [7]);
  and (_13684_, _08560_, _08533_);
  or (_13685_, _13684_, _13683_);
  and (_13686_, _13685_, _06475_);
  or (_13688_, _13686_, _06468_);
  or (_13689_, _13688_, _13681_);
  and (_13690_, _13689_, _13669_);
  or (_13691_, _13690_, _06466_);
  or (_13692_, _13674_, _06801_);
  and (_13693_, _13692_, _06484_);
  and (_13694_, _13693_, _13691_);
  and (_13695_, _08698_, _08533_);
  or (_13696_, _13695_, _13683_);
  and (_13697_, _13696_, _06483_);
  or (_13699_, _13697_, _13694_);
  and (_13700_, _13699_, _07164_);
  and (_13701_, _08707_, _08533_);
  or (_13702_, _13701_, _13683_);
  and (_13703_, _13702_, _06461_);
  or (_13704_, _13703_, _13700_);
  and (_13705_, _13704_, _06242_);
  and (_13706_, _08726_, _08533_);
  or (_13707_, _13706_, _13683_);
  and (_13708_, _13707_, _06241_);
  or (_13710_, _13708_, _07187_);
  or (_13711_, _13710_, _13705_);
  and (_13712_, _13711_, _13668_);
  or (_13713_, _13712_, _07182_);
  and (_13714_, _08671_, _07943_);
  or (_13715_, _13661_, _07183_);
  or (_13716_, _13715_, _13714_);
  and (_13717_, _13716_, _06336_);
  and (_13718_, _13717_, _13713_);
  and (_13719_, _08966_, _07943_);
  or (_13721_, _13719_, _13661_);
  and (_13722_, _13721_, _05968_);
  or (_13723_, _13722_, _06371_);
  or (_13724_, _13723_, _13718_);
  and (_13725_, _08770_, _07943_);
  or (_13726_, _13725_, _13661_);
  or (_13727_, _13726_, _07198_);
  and (_13728_, _13727_, _13724_);
  or (_13729_, _13728_, _06367_);
  and (_13730_, _08988_, _07943_);
  or (_13732_, _13730_, _13661_);
  or (_13733_, _13732_, _07218_);
  and (_13734_, _13733_, _07216_);
  and (_13735_, _13734_, _13729_);
  or (_13736_, _13735_, _13664_);
  and (_13737_, _13736_, _07213_);
  or (_13738_, _13661_, _08007_);
  and (_13739_, _13726_, _06366_);
  and (_13740_, _13739_, _13738_);
  or (_13741_, _13740_, _13737_);
  and (_13743_, _13741_, _07210_);
  and (_13744_, _13674_, _06541_);
  and (_13745_, _13744_, _13738_);
  or (_13746_, _13745_, _06383_);
  or (_13747_, _13746_, _13743_);
  and (_13748_, _08985_, _07943_);
  or (_13749_, _13661_, _07231_);
  or (_13750_, _13749_, _13748_);
  and (_13751_, _13750_, _07229_);
  and (_13752_, _13751_, _13747_);
  nor (_13753_, _08508_, _13660_);
  or (_13754_, _13753_, _13661_);
  and (_13755_, _13754_, _06528_);
  or (_13756_, _13755_, _06563_);
  or (_13757_, _13756_, _13752_);
  or (_13758_, _13671_, _07241_);
  and (_13759_, _13758_, _06571_);
  and (_13760_, _13759_, _13757_);
  and (_13761_, _13696_, _06199_);
  or (_13762_, _13761_, _06188_);
  or (_13763_, _13762_, _13760_);
  and (_13764_, _08503_, _07943_);
  or (_13765_, _13661_, _06189_);
  or (_13766_, _13765_, _13764_);
  and (_13767_, _13766_, _01452_);
  and (_13768_, _13767_, _13763_);
  or (_13769_, _13768_, _13659_);
  and (_41200_, _13769_, _43223_);
  not (_13770_, \oc8051_golden_model_1.SP [7]);
  nor (_13771_, _07928_, _13770_);
  and (_13772_, _08509_, _08135_);
  or (_13773_, _13772_, _13771_);
  and (_13774_, _13773_, _06533_);
  not (_13775_, _08135_);
  nor (_13776_, _08004_, _13775_);
  or (_13777_, _13771_, _07182_);
  or (_13778_, _13777_, _13776_);
  and (_13779_, _13778_, _12604_);
  and (_13780_, _08685_, _08135_);
  or (_13781_, _13780_, _13771_);
  or (_13782_, _13781_, _06252_);
  nor (_13783_, _07123_, _13770_);
  and (_13784_, _07928_, \oc8051_golden_model_1.ACC [7]);
  or (_13785_, _13784_, _13771_);
  and (_13786_, _13785_, _07123_);
  or (_13787_, _13786_, _13783_);
  and (_13788_, _13787_, _07272_);
  and (_13789_, _07719_, \oc8051_golden_model_1.SP [4]);
  and (_13790_, _13789_, \oc8051_golden_model_1.SP [5]);
  and (_13791_, _13790_, \oc8051_golden_model_1.SP [6]);
  or (_13792_, _13791_, \oc8051_golden_model_1.SP [7]);
  nand (_13793_, _13791_, \oc8051_golden_model_1.SP [7]);
  and (_13794_, _13793_, _13792_);
  and (_13795_, _13794_, _06705_);
  or (_13796_, _13795_, _06251_);
  or (_13797_, _13796_, _13788_);
  and (_13798_, _13797_, _05950_);
  and (_13799_, _13798_, _13782_);
  and (_13800_, _13794_, _07474_);
  or (_13801_, _13800_, _06468_);
  or (_13802_, _13801_, _13799_);
  not (_13803_, \oc8051_golden_model_1.SP [6]);
  not (_13804_, \oc8051_golden_model_1.SP [5]);
  not (_13805_, \oc8051_golden_model_1.SP [4]);
  and (_13806_, _08592_, _13805_);
  and (_13807_, _13806_, _13804_);
  and (_13808_, _13807_, _13803_);
  and (_13809_, _13808_, _06235_);
  nor (_13810_, _13809_, _13770_);
  and (_13811_, _13809_, _13770_);
  nor (_13812_, _13811_, _13810_);
  nand (_13813_, _13812_, _06468_);
  and (_13814_, _13813_, _13802_);
  or (_13815_, _13814_, _06466_);
  or (_13816_, _13785_, _06801_);
  and (_13817_, _13816_, _07523_);
  and (_13818_, _13817_, _13815_);
  and (_13819_, _13790_, \oc8051_golden_model_1.SP [0]);
  and (_13820_, _13819_, \oc8051_golden_model_1.SP [6]);
  nor (_13821_, _13820_, _13770_);
  and (_13822_, _13820_, _13770_);
  or (_13823_, _13822_, _13821_);
  and (_13824_, _13823_, _06247_);
  or (_13825_, _13824_, _07472_);
  or (_13826_, _13825_, _13818_);
  or (_13827_, _13794_, _07473_);
  and (_13828_, _13827_, _07188_);
  and (_13829_, _13828_, _13826_);
  or (_13830_, _13829_, _13779_);
  or (_13831_, _13771_, _07183_);
  and (_13832_, _08671_, _07928_);
  or (_13833_, _13832_, _13831_);
  and (_13834_, _13833_, _06336_);
  and (_13835_, _13834_, _13830_);
  and (_13836_, _08966_, _08135_);
  or (_13837_, _13836_, _13771_);
  and (_13838_, _13837_, _05968_);
  or (_13839_, _13838_, _06371_);
  or (_13840_, _13839_, _13835_);
  and (_13841_, _08770_, _07928_);
  or (_13842_, _13841_, _13771_);
  or (_13843_, _13842_, _07198_);
  and (_13844_, _13843_, _13840_);
  or (_13845_, _13844_, _05895_);
  not (_13846_, _05895_);
  or (_13847_, _13794_, _13846_);
  and (_13848_, _13847_, _13845_);
  or (_13849_, _13848_, _06367_);
  and (_13850_, _08988_, _07928_);
  or (_13851_, _13850_, _13771_);
  or (_13852_, _13851_, _07218_);
  and (_13853_, _13852_, _07216_);
  and (_13854_, _13853_, _13849_);
  or (_13855_, _13854_, _13774_);
  and (_13856_, _13855_, _07213_);
  or (_13857_, _13771_, _08007_);
  and (_13858_, _13842_, _06366_);
  and (_13859_, _13858_, _13857_);
  or (_13860_, _13859_, _13856_);
  and (_13861_, _13860_, _12719_);
  and (_13862_, _13785_, _06541_);
  and (_13863_, _13862_, _13857_);
  and (_13864_, _13794_, _07209_);
  or (_13865_, _13864_, _06383_);
  or (_13866_, _13865_, _13863_);
  or (_13867_, _13866_, _13861_);
  and (_13868_, _08985_, _07928_);
  or (_13869_, _13868_, _13771_);
  or (_13870_, _13869_, _07231_);
  and (_13871_, _13870_, _13867_);
  or (_13872_, _13871_, _06528_);
  not (_13873_, _06547_);
  nor (_13874_, _08508_, _13775_);
  or (_13875_, _13771_, _07229_);
  or (_13876_, _13875_, _13874_);
  and (_13877_, _13876_, _13873_);
  and (_13878_, _13877_, _13872_);
  or (_13879_, _13808_, \oc8051_golden_model_1.SP [7]);
  nand (_13880_, _13808_, \oc8051_golden_model_1.SP [7]);
  and (_13881_, _13880_, _13879_);
  and (_13882_, _13881_, _06547_);
  or (_13883_, _13882_, _07228_);
  or (_13884_, _13883_, _13878_);
  or (_13885_, _13794_, _05916_);
  and (_13886_, _13885_, _13884_);
  or (_13887_, _13886_, _06260_);
  or (_13888_, _13881_, _06261_);
  and (_13889_, _13888_, _07241_);
  and (_13890_, _13889_, _13887_);
  and (_13891_, _13781_, _06563_);
  or (_13892_, _13891_, _07812_);
  or (_13893_, _13892_, _13890_);
  or (_13894_, _13794_, _07250_);
  and (_13895_, _13894_, _06189_);
  and (_13896_, _13895_, _13893_);
  and (_13897_, _08503_, _08135_);
  or (_13898_, _13897_, _13771_);
  and (_13899_, _13898_, _06188_);
  or (_13900_, _13899_, _01456_);
  or (_13901_, _13900_, _13896_);
  or (_13902_, _01452_, \oc8051_golden_model_1.SP [7]);
  and (_13903_, _13902_, _43223_);
  and (_41201_, _13903_, _13901_);
  not (_13904_, _07857_);
  and (_13905_, _13904_, \oc8051_golden_model_1.SBUF [7]);
  and (_13906_, _08509_, _07857_);
  or (_13907_, _13906_, _13905_);
  and (_13908_, _13907_, _06533_);
  nor (_13909_, _08004_, _13904_);
  or (_13910_, _13909_, _13905_);
  or (_13911_, _13910_, _07188_);
  and (_13912_, _08685_, _07857_);
  or (_13913_, _13912_, _13905_);
  or (_13914_, _13913_, _06252_);
  and (_13915_, _07857_, \oc8051_golden_model_1.ACC [7]);
  or (_13916_, _13915_, _13905_);
  and (_13917_, _13916_, _07123_);
  and (_13918_, _07124_, \oc8051_golden_model_1.SBUF [7]);
  or (_13919_, _13918_, _06251_);
  or (_13920_, _13919_, _13917_);
  and (_13921_, _13920_, _07142_);
  and (_13922_, _13921_, _13914_);
  and (_13923_, _13910_, _06468_);
  or (_13924_, _13923_, _13922_);
  and (_13925_, _13924_, _06801_);
  and (_13926_, _13916_, _06466_);
  or (_13927_, _13926_, _07187_);
  or (_13928_, _13927_, _13925_);
  and (_13929_, _13928_, _13911_);
  or (_13930_, _13929_, _07182_);
  and (_13931_, _08671_, _07857_);
  or (_13932_, _13905_, _07183_);
  or (_13933_, _13932_, _13931_);
  and (_13934_, _13933_, _06336_);
  and (_13935_, _13934_, _13930_);
  and (_13936_, _08966_, _07857_);
  or (_13937_, _13936_, _13905_);
  and (_13938_, _13937_, _05968_);
  or (_13939_, _13938_, _06371_);
  or (_13940_, _13939_, _13935_);
  and (_13941_, _08770_, _07857_);
  or (_13942_, _13941_, _13905_);
  or (_13943_, _13942_, _07198_);
  and (_13944_, _13943_, _13940_);
  or (_13945_, _13944_, _06367_);
  and (_13946_, _08988_, _07857_);
  or (_13947_, _13946_, _13905_);
  or (_13948_, _13947_, _07218_);
  and (_13949_, _13948_, _07216_);
  and (_13950_, _13949_, _13945_);
  or (_13951_, _13950_, _13908_);
  and (_13952_, _13951_, _07213_);
  or (_13953_, _13905_, _08007_);
  and (_13954_, _13942_, _06366_);
  and (_13955_, _13954_, _13953_);
  or (_13956_, _13955_, _13952_);
  and (_13957_, _13956_, _07210_);
  and (_13958_, _13916_, _06541_);
  and (_13959_, _13958_, _13953_);
  or (_13960_, _13959_, _06383_);
  or (_13961_, _13960_, _13957_);
  and (_13962_, _08985_, _07857_);
  or (_13963_, _13905_, _07231_);
  or (_13964_, _13963_, _13962_);
  and (_13965_, _13964_, _07229_);
  and (_13966_, _13965_, _13961_);
  nor (_13967_, _08508_, _13904_);
  or (_13968_, _13967_, _13905_);
  and (_13969_, _13968_, _06528_);
  or (_13970_, _13969_, _06563_);
  or (_13971_, _13970_, _13966_);
  or (_13972_, _13913_, _07241_);
  and (_13973_, _13972_, _06189_);
  and (_13974_, _13973_, _13971_);
  and (_13975_, _08503_, _07857_);
  or (_13976_, _13975_, _13905_);
  and (_13977_, _13976_, _06188_);
  or (_13978_, _13977_, _01456_);
  or (_13979_, _13978_, _13974_);
  or (_13980_, _01452_, \oc8051_golden_model_1.SBUF [7]);
  and (_13981_, _13980_, _43223_);
  and (_41202_, _13981_, _13979_);
  nor (_13982_, _01452_, _10854_);
  nor (_13983_, _08543_, _10854_);
  and (_13984_, _08698_, _08543_);
  or (_13985_, _13984_, _13983_);
  or (_13986_, _13985_, _06571_);
  nor (_13987_, _07907_, _10854_);
  and (_13988_, _08509_, _07907_);
  or (_13989_, _13988_, _13987_);
  and (_13990_, _13989_, _06533_);
  and (_13991_, _08966_, _07907_);
  or (_13992_, _13991_, _13987_);
  and (_13993_, _13992_, _05968_);
  not (_13994_, _07907_);
  nor (_13995_, _08004_, _13994_);
  or (_13996_, _13995_, _13987_);
  or (_13997_, _13996_, _07188_);
  and (_13998_, _10550_, _08007_);
  and (_13999_, _10560_, _10556_);
  nor (_14000_, _13999_, _10554_);
  nand (_14001_, _10602_, _10556_);
  or (_14002_, _14001_, _10600_);
  and (_14003_, _14002_, _14000_);
  or (_14004_, _14003_, _13998_);
  and (_14005_, _14004_, _06510_);
  not (_14006_, _06504_);
  not (_14007_, _06505_);
  nor (_14008_, _12954_, _14007_);
  and (_14009_, _08560_, _08543_);
  or (_14010_, _14009_, _13983_);
  or (_14011_, _13983_, _08706_);
  and (_14012_, _14011_, _06461_);
  and (_14013_, _14012_, _14010_);
  and (_14014_, _08685_, _07907_);
  or (_14015_, _14014_, _13987_);
  or (_14016_, _14015_, _06252_);
  and (_14017_, _07907_, \oc8051_golden_model_1.ACC [7]);
  or (_14018_, _14017_, _13987_);
  and (_14019_, _14018_, _07123_);
  nor (_14020_, _07123_, _10854_);
  or (_14021_, _14020_, _06251_);
  or (_14022_, _14021_, _14019_);
  and (_14023_, _14022_, _10719_);
  and (_14024_, _14023_, _14016_);
  nor (_14025_, _10738_, _10719_);
  or (_14026_, _12442_, _06475_);
  or (_14027_, _14026_, _14025_);
  or (_14028_, _14027_, _14024_);
  or (_14029_, _14010_, _06476_);
  and (_14030_, _14029_, _07142_);
  and (_14031_, _14030_, _14028_);
  and (_14032_, _13996_, _06468_);
  or (_14033_, _14032_, _06466_);
  or (_14034_, _14033_, _14031_);
  or (_14035_, _14018_, _06801_);
  nor (_14036_, _12461_, _06483_);
  and (_14037_, _14036_, _14035_);
  and (_14038_, _14037_, _14034_);
  and (_14039_, _13985_, _06483_);
  or (_14040_, _14039_, _12479_);
  or (_14041_, _14040_, _14038_);
  not (_14042_, _12513_);
  and (_14043_, _12508_, _12504_);
  or (_14044_, _12505_, _14043_);
  and (_14045_, _14044_, _12503_);
  and (_14046_, _12500_, _12498_);
  or (_14047_, _14046_, _12497_);
  or (_14048_, _14047_, _14045_);
  and (_14049_, _14048_, _12496_);
  or (_14050_, _12492_, _12489_);
  and (_14051_, _12487_, _14050_);
  and (_14052_, _14051_, _12488_);
  and (_14053_, _12485_, _08005_);
  or (_14054_, _14053_, _12482_);
  or (_14055_, _14054_, _14052_);
  or (_14056_, _14055_, _14049_);
  and (_14057_, _14056_, _14042_);
  or (_14058_, _14057_, _12478_);
  and (_14059_, _14058_, _06345_);
  and (_14060_, _14059_, _14041_);
  not (_14061_, _12385_);
  and (_14062_, _14061_, _12383_);
  not (_14063_, _12380_);
  nand (_14064_, _12378_, _14063_);
  nand (_14065_, _14064_, _12377_);
  or (_14066_, _14065_, _12389_);
  or (_14067_, _14066_, _14062_);
  and (_14068_, _14067_, _12376_);
  nand (_14069_, _12373_, _12370_);
  and (_14070_, _12368_, _14069_);
  and (_14071_, _14070_, _12369_);
  nand (_14072_, _12363_, _12365_);
  and (_14073_, _14072_, _08718_);
  or (_14074_, _14073_, _14071_);
  or (_14075_, _14074_, _14068_);
  nor (_14076_, _12392_, _06345_);
  and (_14077_, _14076_, _14075_);
  or (_14078_, _14077_, _14060_);
  and (_14079_, _14078_, _12536_);
  nand (_14080_, _08211_, \oc8051_golden_model_1.ACC [5]);
  nor (_14081_, _08211_, \oc8051_golden_model_1.ACC [5]);
  nor (_14082_, _08496_, \oc8051_golden_model_1.ACC [4]);
  or (_14083_, _14082_, _14081_);
  and (_14084_, _14083_, _14080_);
  and (_14085_, _14084_, _12531_);
  nor (_14086_, _08006_, \oc8051_golden_model_1.ACC [7]);
  or (_14087_, _08108_, \oc8051_golden_model_1.ACC [6]);
  nor (_14088_, _14087_, _08509_);
  or (_14089_, _14088_, _14086_);
  or (_14090_, _14089_, _14085_);
  nand (_14091_, _08256_, \oc8051_golden_model_1.ACC [3]);
  nor (_14092_, _08256_, \oc8051_golden_model_1.ACC [3]);
  nor (_14093_, _08396_, \oc8051_golden_model_1.ACC [2]);
  or (_14094_, _14093_, _14092_);
  and (_14095_, _14094_, _14091_);
  nor (_14096_, _08301_, \oc8051_golden_model_1.ACC [1]);
  nor (_14097_, _08351_, _05997_);
  nor (_14098_, _14097_, _11217_);
  or (_14099_, _14098_, _14096_);
  and (_14100_, _14099_, _12524_);
  or (_14101_, _14100_, _14095_);
  and (_14102_, _14101_, _12532_);
  or (_14103_, _14102_, _14090_);
  nor (_14104_, _12533_, _12536_);
  and (_14105_, _14104_, _14103_);
  or (_14106_, _14105_, _14079_);
  and (_14107_, _14106_, _12522_);
  and (_14108_, _06187_, _08506_);
  or (_14109_, _06326_, \oc8051_golden_model_1.ACC [6]);
  nor (_14110_, _14109_, _10942_);
  or (_14111_, _14110_, _14108_);
  not (_14112_, _12549_);
  nor (_14113_, _06230_, \oc8051_golden_model_1.ACC [4]);
  or (_14114_, _14113_, _12548_);
  and (_14115_, _14114_, _14112_);
  and (_14116_, _14115_, _12553_);
  or (_14117_, _14116_, _14111_);
  nor (_14118_, _06292_, \oc8051_golden_model_1.ACC [3]);
  nand (_14119_, _06292_, \oc8051_golden_model_1.ACC [3]);
  nor (_14120_, _06750_, \oc8051_golden_model_1.ACC [2]);
  and (_14121_, _14120_, _14119_);
  or (_14122_, _14121_, _14118_);
  nor (_14123_, _06155_, \oc8051_golden_model_1.ACC [1]);
  and (_14124_, _06155_, \oc8051_golden_model_1.ACC [1]);
  and (_14125_, _06802_, \oc8051_golden_model_1.ACC [0]);
  nor (_14126_, _14125_, _14124_);
  or (_14127_, _14126_, _14123_);
  and (_14128_, _14127_, _12543_);
  or (_14129_, _14128_, _14122_);
  and (_14130_, _14129_, _12554_);
  or (_14131_, _14130_, _14117_);
  nor (_14132_, _12555_, _12522_);
  and (_14133_, _14132_, _14131_);
  or (_14134_, _14133_, _12245_);
  or (_14135_, _14134_, _14107_);
  nand (_14136_, _12245_, \oc8051_golden_model_1.PSW [7]);
  and (_14137_, _14136_, _07164_);
  and (_14138_, _14137_, _14135_);
  nor (_14139_, _14138_, _14013_);
  nor (_14140_, _14139_, _06460_);
  and (_14141_, _06460_, \oc8051_golden_model_1.PSW [7]);
  and (_14142_, _14141_, _12954_);
  or (_14143_, _14142_, _14140_);
  nor (_14144_, _09487_, _06505_);
  and (_14145_, _14144_, _14143_);
  or (_14146_, _14145_, _14008_);
  and (_14147_, _14146_, _14006_);
  and (_14148_, _07492_, _05969_);
  nor (_14149_, _06359_, _06710_);
  or (_14150_, _14149_, _14148_);
  and (_14151_, _06361_, _05969_);
  nor (_14152_, _14151_, _14150_);
  or (_14153_, _12954_, \oc8051_golden_model_1.PSW [7]);
  nand (_14154_, _14153_, _06504_);
  nand (_14155_, _14154_, _14152_);
  or (_14156_, _14155_, _14147_);
  and (_14157_, _05969_, _06348_);
  and (_14158_, _10469_, _10465_);
  nor (_14159_, _14158_, _10463_);
  nand (_14160_, _10471_, _10465_);
  or (_14161_, _14160_, _10796_);
  and (_14162_, _14161_, _14159_);
  or (_14163_, _14162_, _10461_);
  nor (_14164_, _14163_, _14152_);
  nor (_14165_, _14164_, _14157_);
  and (_14166_, _14165_, _14156_);
  and (_14167_, _14163_, _14157_);
  or (_14168_, _14167_, _10610_);
  or (_14169_, _14168_, _14166_);
  and (_14170_, _10623_, _10618_);
  nor (_14171_, _14170_, _10616_);
  nand (_14172_, _10673_, _10618_);
  or (_14173_, _14172_, _10671_);
  and (_14174_, _14173_, _14171_);
  and (_14175_, _10612_, _08671_);
  or (_14176_, _14175_, _10611_);
  or (_14177_, _14176_, _14174_);
  and (_14178_, _14177_, _06516_);
  and (_14179_, _14178_, _14169_);
  or (_14180_, _14179_, _14005_);
  and (_14181_, _14180_, _10543_);
  and (_14182_, _10810_, _07910_);
  and (_14183_, _10822_, _10818_);
  nor (_14184_, _14183_, _10816_);
  nand (_14185_, _10868_, _10818_);
  or (_14186_, _14185_, _10866_);
  and (_14187_, _14186_, _14184_);
  or (_14188_, _14187_, _14182_);
  and (_14189_, _14188_, _10542_);
  or (_14190_, _14189_, _07187_);
  or (_14191_, _14190_, _14181_);
  and (_14192_, _14191_, _13997_);
  or (_14193_, _14192_, _07182_);
  and (_14194_, _08671_, _07907_);
  or (_14195_, _13987_, _07183_);
  or (_14196_, _14195_, _14194_);
  and (_14197_, _14196_, _06336_);
  and (_14198_, _14197_, _14193_);
  or (_14199_, _14198_, _13993_);
  nor (_14200_, _10046_, _06332_);
  and (_14201_, _14200_, _14199_);
  nor (_14202_, _12954_, _10854_);
  and (_14203_, _14202_, _06332_);
  or (_14204_, _14203_, _06371_);
  or (_14205_, _14204_, _14201_);
  and (_14206_, _08770_, _07907_);
  or (_14207_, _14206_, _13987_);
  or (_14208_, _14207_, _07198_);
  and (_14209_, _14208_, _14205_);
  or (_14210_, _14209_, _06331_);
  nand (_14211_, _12954_, _10854_);
  or (_14212_, _14211_, _06921_);
  and (_14213_, _14212_, _14210_);
  or (_14214_, _14213_, _06367_);
  and (_14215_, _08988_, _07907_);
  or (_14216_, _14215_, _13987_);
  or (_14217_, _14216_, _07218_);
  and (_14218_, _14217_, _07216_);
  and (_14219_, _14218_, _14214_);
  or (_14220_, _14219_, _13990_);
  and (_14221_, _14220_, _07213_);
  or (_14222_, _13987_, _08007_);
  and (_14223_, _14207_, _06366_);
  and (_14224_, _14223_, _14222_);
  or (_14225_, _14224_, _14221_);
  and (_14226_, _14225_, _07210_);
  and (_14227_, _14018_, _06541_);
  and (_14228_, _14227_, _14222_);
  or (_14229_, _14228_, _06383_);
  or (_14230_, _14229_, _14226_);
  and (_14231_, _08985_, _07907_);
  or (_14232_, _13987_, _07231_);
  or (_14233_, _14232_, _14231_);
  and (_14234_, _14233_, _07229_);
  and (_14235_, _14234_, _14230_);
  nor (_14236_, _08508_, _13994_);
  or (_14237_, _14236_, _13987_);
  and (_14238_, _14237_, _06528_);
  or (_14239_, _14238_, _11014_);
  or (_14240_, _14239_, _14235_);
  and (_14241_, _10462_, \oc8051_golden_model_1.ACC [7]);
  or (_14242_, _14241_, _10519_);
  or (_14243_, _14242_, _10461_);
  or (_14244_, _14243_, _10526_);
  and (_14245_, _14244_, _14240_);
  or (_14246_, _14245_, _10452_);
  or (_14247_, _14175_, _11022_);
  nor (_14248_, _10615_, _08506_);
  or (_14249_, _14248_, _11044_);
  or (_14250_, _14249_, _14247_);
  and (_14251_, _14250_, _06538_);
  and (_14252_, _14251_, _14246_);
  nor (_14253_, _10553_, _08506_);
  or (_14254_, _14253_, _11074_);
  or (_14255_, _11050_, _13998_);
  or (_14256_, _14255_, _14254_);
  and (_14257_, _14256_, _11052_);
  or (_14258_, _14257_, _14252_);
  nor (_14259_, _10815_, _08506_);
  or (_14260_, _14259_, _11104_);
  or (_14261_, _14182_, _11082_);
  or (_14262_, _14261_, _14260_);
  and (_14263_, _14262_, _11081_);
  and (_14264_, _14263_, _14258_);
  and (_14265_, _11080_, \oc8051_golden_model_1.ACC [7]);
  or (_14266_, _14265_, _12104_);
  or (_14267_, _14266_, _14264_);
  and (_14268_, _11148_, _10916_);
  nor (_14269_, _11117_, _10528_);
  nor (_14270_, _14269_, _10915_);
  or (_14271_, _14270_, _12103_);
  or (_14272_, _14271_, _14268_);
  and (_14273_, _14272_, _14267_);
  or (_14274_, _14273_, _11156_);
  and (_14275_, _11191_, _10935_);
  nor (_14276_, _11161_, _10934_);
  nor (_14277_, _14276_, _10933_);
  or (_14278_, _14277_, _11160_);
  or (_14279_, _14278_, _14275_);
  and (_14280_, _14279_, _06295_);
  and (_14281_, _14280_, _14274_);
  not (_14282_, _08508_);
  not (_14283_, _08507_);
  nand (_14284_, _11232_, _14283_);
  and (_14285_, _14284_, _06293_);
  and (_14286_, _14285_, _14282_);
  or (_14287_, _14286_, _10450_);
  or (_14288_, _14287_, _14281_);
  nor (_14289_, _11270_, _10940_);
  or (_14290_, _14289_, _10451_);
  or (_14291_, _14290_, _10941_);
  and (_14292_, _14291_, _14288_);
  or (_14293_, _14292_, _06563_);
  nor (_14294_, _14015_, _07241_);
  nor (_14295_, _14294_, _11284_);
  and (_14296_, _14295_, _14293_);
  and (_14297_, _11284_, \oc8051_golden_model_1.ACC [0]);
  or (_14298_, _14297_, _06199_);
  or (_14299_, _14298_, _14296_);
  and (_14300_, _14299_, _13986_);
  or (_14301_, _14300_, _06188_);
  and (_14302_, _08503_, _07907_);
  or (_14303_, _13987_, _06189_);
  or (_14304_, _14303_, _14302_);
  and (_14305_, _14304_, _01452_);
  and (_14306_, _14305_, _14301_);
  or (_14307_, _14306_, _13982_);
  and (_41203_, _14307_, _43223_);
  nor (_14308_, _07659_, _07508_);
  nor (_14309_, _07831_, _14308_);
  nor (_14310_, _07508_, _07263_);
  nor (_14311_, _07509_, _14310_);
  and (_14312_, _14311_, _07507_);
  and (_14313_, _14312_, _14309_);
  or (_14314_, _14313_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_14315_, _07844_, _07837_);
  nor (_14316_, _07845_, _14315_);
  and (_14317_, _07844_, _06236_);
  nand (_14318_, _14317_, _14316_);
  and (_14319_, _14318_, _14314_);
  not (_14320_, _14313_);
  not (_14321_, _06190_);
  nor (_14322_, _08351_, _14321_);
  nand (_14323_, _05912_, _05557_);
  not (_14324_, _07230_);
  or (_14325_, _08351_, _08908_);
  and (_14326_, _14325_, _07232_);
  nand (_14327_, _05895_, _05557_);
  or (_14328_, _08351_, _07523_);
  nor (_14329_, _12875_, _12851_);
  or (_14330_, _14329_, _08697_);
  nor (_14331_, _08351_, _08675_);
  nand (_14332_, _08572_, _07325_);
  nand (_14333_, _06705_, _05557_);
  or (_14334_, _06705_, \oc8051_golden_model_1.ACC [0]);
  and (_14335_, _14334_, _14333_);
  nor (_14336_, _14335_, _08572_);
  nor (_14337_, _14336_, _06253_);
  and (_14338_, _14337_, _14332_);
  or (_14339_, _14338_, _14331_);
  and (_14340_, _14339_, _08520_);
  nand (_14341_, _12875_, _12852_);
  and (_14342_, _14341_, _07139_);
  or (_14343_, _14342_, _07474_);
  or (_14344_, _14343_, _14340_);
  nor (_14345_, _05950_, \oc8051_golden_model_1.PC [0]);
  nor (_14346_, _14345_, _07143_);
  and (_14347_, _14346_, _14344_);
  and (_14348_, _07143_, _07325_);
  or (_14349_, _14348_, _07159_);
  or (_14350_, _14349_, _14347_);
  and (_14351_, _14350_, _14330_);
  or (_14352_, _14351_, _06247_);
  and (_14353_, _14352_, _14328_);
  or (_14354_, _14353_, _07165_);
  not (_14355_, _12876_);
  and (_14356_, _14341_, _14355_);
  or (_14357_, _14356_, _07270_);
  and (_14358_, _14357_, _05947_);
  and (_14359_, _14358_, _14354_);
  or (_14360_, _05947_, _05557_);
  nand (_14361_, _06497_, _14360_);
  or (_14362_, _14361_, _14359_);
  or (_14363_, _08351_, _06497_);
  and (_14364_, _14363_, _14362_);
  or (_14365_, _14364_, _07174_);
  and (_14366_, _09342_, _07904_);
  or (_14367_, _14366_, _08349_);
  or (_14368_, _14367_, _07369_);
  and (_14369_, _14368_, _08724_);
  and (_14370_, _14369_, _14365_);
  nand (_14371_, _12851_, _10854_);
  and (_14372_, _14371_, _14341_);
  and (_14373_, _14372_, _06243_);
  or (_14374_, _14373_, _05970_);
  or (_14375_, _14374_, _14370_);
  and (_14376_, _05970_, _05557_);
  nor (_14377_, _14376_, _07189_);
  and (_14378_, _14377_, _14375_);
  and (_14379_, _07189_, _07325_);
  or (_14380_, _14379_, _07184_);
  or (_14381_, _14380_, _14378_);
  or (_14382_, _09342_, _07185_);
  and (_14383_, _14382_, _08735_);
  and (_14384_, _14383_, _14381_);
  and (_14385_, _08769_, _07325_);
  and (_14386_, _08906_, \oc8051_golden_model_1.P0 [0]);
  and (_14387_, _08932_, \oc8051_golden_model_1.SBUF [0]);
  or (_14388_, _14387_, _14386_);
  and (_14389_, _08903_, \oc8051_golden_model_1.P1 [0]);
  and (_14390_, _08930_, \oc8051_golden_model_1.SCON [0]);
  or (_14391_, _14390_, _14389_);
  or (_14392_, _14391_, _14388_);
  and (_14393_, _08900_, \oc8051_golden_model_1.TCON [0]);
  and (_14394_, _08875_, \oc8051_golden_model_1.TL0 [0]);
  or (_14395_, _14394_, _14393_);
  and (_14396_, _08912_, \oc8051_golden_model_1.TMOD [0]);
  and (_14397_, _08894_, \oc8051_golden_model_1.PSW [0]);
  or (_14398_, _14397_, _14396_);
  or (_14399_, _14398_, _14395_);
  and (_14400_, _08884_, \oc8051_golden_model_1.B [0]);
  and (_14401_, _08890_, \oc8051_golden_model_1.ACC [0]);
  or (_14402_, _14401_, _14400_);
  and (_14403_, _08926_, \oc8051_golden_model_1.IE [0]);
  and (_14404_, _08917_, \oc8051_golden_model_1.P3 [0]);
  or (_14405_, _14404_, _14403_);
  and (_14406_, _08924_, \oc8051_golden_model_1.P2 [0]);
  and (_14407_, _08919_, \oc8051_golden_model_1.IP [0]);
  or (_14408_, _14407_, _14406_);
  or (_14409_, _14408_, _14405_);
  or (_14410_, _14409_, _14402_);
  or (_14411_, _14410_, _14399_);
  or (_14412_, _14411_, _14392_);
  and (_14413_, _08953_, \oc8051_golden_model_1.TH0 [0]);
  and (_14414_, _08943_, \oc8051_golden_model_1.DPL [0]);
  and (_14415_, _08960_, \oc8051_golden_model_1.SP [0]);
  or (_14416_, _14415_, _14414_);
  or (_14417_, _14416_, _14413_);
  and (_14418_, _08940_, \oc8051_golden_model_1.TL1 [0]);
  and (_14419_, _08958_, \oc8051_golden_model_1.DPH [0]);
  or (_14420_, _14419_, _14418_);
  and (_14421_, _08947_, \oc8051_golden_model_1.PCON [0]);
  and (_14422_, _08955_, \oc8051_golden_model_1.TH1 [0]);
  or (_14423_, _14422_, _14421_);
  or (_14424_, _14423_, _14420_);
  or (_14425_, _14424_, _14417_);
  or (_14426_, _14425_, _14412_);
  or (_14427_, _14426_, _14385_);
  and (_14428_, _14427_, _07186_);
  or (_14429_, _14428_, _08973_);
  or (_14430_, _14429_, _14384_);
  and (_14431_, _08973_, _06802_);
  nor (_14432_, _14431_, _07199_);
  and (_14433_, _14432_, _14430_);
  and (_14434_, _07199_, _08908_);
  or (_14435_, _14434_, _05895_);
  or (_14436_, _14435_, _14433_);
  and (_14437_, _14436_, _14327_);
  or (_14438_, _14437_, _07219_);
  not (_14439_, _07219_);
  and (_14440_, _08351_, _08908_);
  not (_14441_, _14440_);
  and (_14442_, _14441_, _14325_);
  or (_14443_, _14442_, _14439_);
  and (_14444_, _14443_, _08511_);
  and (_14445_, _14444_, _14438_);
  nor (_14446_, _12527_, _08511_);
  or (_14447_, _14446_, _07214_);
  or (_14448_, _14447_, _14445_);
  or (_14449_, _14440_, _07215_);
  and (_14450_, _14449_, _07212_);
  and (_14451_, _14450_, _14448_);
  and (_14452_, _11218_, _07211_);
  or (_14453_, _14452_, _07209_);
  or (_14454_, _14453_, _14451_);
  nor (_14455_, _05919_, \oc8051_golden_model_1.PC [0]);
  nor (_14456_, _14455_, _07232_);
  and (_14457_, _14456_, _14454_);
  or (_14458_, _14457_, _14326_);
  and (_14459_, _14458_, _14324_);
  nor (_14460_, _12526_, _14324_);
  or (_14461_, _14460_, _07228_);
  or (_14462_, _14461_, _14459_);
  or (_14463_, _05916_, \oc8051_golden_model_1.PC [0]);
  and (_14464_, _14463_, _12983_);
  and (_14465_, _14464_, _14462_);
  nor (_14466_, _12983_, _07325_);
  or (_14467_, _14466_, _07243_);
  or (_14468_, _14467_, _14465_);
  nand (_14469_, _09342_, _07243_);
  and (_14470_, _14469_, _14468_);
  or (_14471_, _14470_, _07242_);
  nand (_14472_, _08351_, _07242_);
  and (_14473_, _14472_, _08505_);
  and (_14474_, _14473_, _14471_);
  and (_14475_, _06378_, _05557_);
  or (_14476_, _14475_, _05912_);
  or (_14477_, _14476_, _14474_);
  and (_14478_, _14477_, _14323_);
  or (_14479_, _14478_, _07249_);
  or (_14480_, _14329_, _07265_);
  and (_14481_, _14480_, _09371_);
  and (_14482_, _14481_, _14479_);
  nor (_14483_, _09371_, _07325_);
  or (_14484_, _14483_, _07259_);
  or (_14485_, _14484_, _14482_);
  nand (_14486_, _09342_, _07259_);
  and (_14487_, _14486_, _14321_);
  and (_14488_, _14487_, _14485_);
  or (_14489_, _14488_, _14322_);
  or (_14490_, _14489_, _14320_);
  and (_14491_, _14490_, _14319_);
  and (_14492_, _14316_, _06236_);
  nand (_14493_, _12280_, _06378_);
  or (_14494_, _12185_, _06378_);
  and (_14495_, _14494_, _14493_);
  and (_14496_, _14495_, _07844_);
  and (_14497_, _14496_, _14492_);
  or (_41219_, _14497_, _14491_);
  or (_14498_, _14313_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_14499_, _14498_, _14318_);
  not (_14500_, _06976_);
  nor (_14501_, _09394_, _09343_);
  or (_14502_, _14501_, _14500_);
  nor (_14503_, _08678_, _08352_);
  nand (_14504_, _14503_, _07242_);
  not (_14505_, _06963_);
  and (_14506_, _07455_, _05911_);
  not (_14507_, _14506_);
  nor (_14508_, _05916_, \oc8051_golden_model_1.PC [1]);
  not (_14509_, _12822_);
  nand (_14510_, _12821_, _12799_);
  and (_14511_, _14510_, _07165_);
  and (_14512_, _14511_, _14509_);
  nor (_14513_, _12821_, _08134_);
  or (_14514_, _14513_, _08697_);
  nor (_14515_, _09382_, _08565_);
  nand (_14516_, _14515_, _08572_);
  and (_14517_, _06705_, _05550_);
  nor (_14518_, _06705_, _05937_);
  or (_14519_, _14518_, _14517_);
  or (_14520_, _14519_, _08572_);
  and (_14521_, _14520_, _14516_);
  or (_14522_, _14521_, _06253_);
  nand (_14523_, _14503_, _06253_);
  and (_14524_, _14523_, _14522_);
  or (_14525_, _14524_, _07139_);
  or (_14526_, _14510_, _08520_);
  and (_14527_, _14526_, _14525_);
  or (_14528_, _14527_, _07474_);
  nor (_14529_, _05950_, _05550_);
  nor (_14530_, _14529_, _07143_);
  and (_14531_, _14530_, _14528_);
  and (_14532_, _09381_, _07143_);
  or (_14533_, _14532_, _07159_);
  or (_14534_, _14533_, _14531_);
  and (_14535_, _14534_, _14514_);
  or (_14536_, _14535_, _06247_);
  nand (_14537_, _08301_, _06247_);
  and (_14538_, _14537_, _07270_);
  and (_14539_, _14538_, _14536_);
  or (_14540_, _14539_, _14512_);
  and (_14541_, _14540_, _05947_);
  or (_14542_, _05947_, \oc8051_golden_model_1.PC [1]);
  nand (_14543_, _06497_, _14542_);
  or (_14544_, _14543_, _14541_);
  nand (_14545_, _08301_, _06498_);
  and (_14546_, _14545_, _14544_);
  or (_14547_, _14546_, _07174_);
  nand (_14548_, _09297_, _07904_);
  nand (_14549_, _14548_, _08299_);
  or (_14550_, _14549_, _07369_);
  and (_14551_, _14550_, _08724_);
  and (_14552_, _14551_, _14547_);
  nand (_14553_, _08134_, _10854_);
  and (_14554_, _14553_, _06243_);
  and (_14555_, _14554_, _14510_);
  or (_14556_, _14555_, _05970_);
  or (_14557_, _14556_, _14552_);
  and (_14558_, _05970_, \oc8051_golden_model_1.PC [1]);
  nor (_14559_, _14558_, _07189_);
  and (_14560_, _14559_, _14557_);
  nor (_14561_, _07120_, _08512_);
  or (_14562_, _14561_, _07184_);
  or (_14563_, _14562_, _14560_);
  or (_14564_, _09297_, _07185_);
  and (_14565_, _14564_, _08735_);
  and (_14566_, _14565_, _14563_);
  nor (_14567_, _08770_, _07120_);
  and (_14568_, _08875_, \oc8051_golden_model_1.TL0 [1]);
  and (_14569_, _08884_, \oc8051_golden_model_1.B [1]);
  or (_14570_, _14569_, _14568_);
  and (_14571_, _08890_, \oc8051_golden_model_1.ACC [1]);
  and (_14572_, _08894_, \oc8051_golden_model_1.PSW [1]);
  or (_14573_, _14572_, _14571_);
  or (_14574_, _14573_, _14570_);
  and (_14575_, _08900_, \oc8051_golden_model_1.TCON [1]);
  and (_14576_, _08930_, \oc8051_golden_model_1.SCON [1]);
  or (_14577_, _14576_, _14575_);
  and (_14578_, _08906_, \oc8051_golden_model_1.P0 [1]);
  and (_14579_, _08912_, \oc8051_golden_model_1.TMOD [1]);
  or (_14580_, _14579_, _14578_);
  or (_14581_, _14580_, _14577_);
  and (_14582_, _08924_, \oc8051_golden_model_1.P2 [1]);
  and (_14583_, _08919_, \oc8051_golden_model_1.IP [1]);
  or (_14584_, _14583_, _14582_);
  and (_14585_, _08926_, \oc8051_golden_model_1.IE [1]);
  and (_14586_, _08917_, \oc8051_golden_model_1.P3 [1]);
  or (_14587_, _14586_, _14585_);
  or (_14588_, _14587_, _14584_);
  and (_14589_, _08903_, \oc8051_golden_model_1.P1 [1]);
  and (_14590_, _08932_, \oc8051_golden_model_1.SBUF [1]);
  or (_14591_, _14590_, _14589_);
  or (_14592_, _14591_, _14588_);
  or (_14593_, _14592_, _14581_);
  or (_14594_, _14593_, _14574_);
  and (_14595_, _08953_, \oc8051_golden_model_1.TH0 [1]);
  and (_14596_, _08943_, \oc8051_golden_model_1.DPL [1]);
  and (_14597_, _08958_, \oc8051_golden_model_1.DPH [1]);
  or (_14598_, _14597_, _14596_);
  or (_14599_, _14598_, _14595_);
  and (_14600_, _08940_, \oc8051_golden_model_1.TL1 [1]);
  and (_14601_, _08955_, \oc8051_golden_model_1.TH1 [1]);
  or (_14602_, _14601_, _14600_);
  and (_14603_, _08947_, \oc8051_golden_model_1.PCON [1]);
  and (_14604_, _08960_, \oc8051_golden_model_1.SP [1]);
  or (_14605_, _14604_, _14603_);
  or (_14606_, _14605_, _14602_);
  or (_14607_, _14606_, _14599_);
  or (_14608_, _14607_, _14594_);
  or (_14609_, _14608_, _14567_);
  and (_14610_, _14609_, _07186_);
  or (_14611_, _14610_, _08973_);
  or (_14612_, _14611_, _14566_);
  and (_14613_, _08973_, _06155_);
  nor (_14614_, _14613_, _07199_);
  and (_14615_, _14614_, _14612_);
  and (_14616_, _07199_, _08870_);
  or (_14617_, _14616_, _05895_);
  or (_14618_, _14617_, _14615_);
  and (_14619_, _05895_, \oc8051_golden_model_1.PC [1]);
  nor (_14620_, _14619_, _07219_);
  and (_14621_, _14620_, _14618_);
  nand (_14622_, _08301_, _07018_);
  nor (_14623_, _08301_, _07018_);
  not (_14624_, _14623_);
  and (_14625_, _14624_, _14622_);
  and (_14626_, _14625_, _07219_);
  or (_14627_, _14626_, _07217_);
  or (_14628_, _14627_, _14621_);
  or (_14629_, _11217_, _08511_);
  and (_14630_, _14629_, _07215_);
  and (_14631_, _14630_, _14628_);
  and (_14632_, _14623_, _07214_);
  or (_14633_, _14632_, _14631_);
  and (_14634_, _14633_, _07212_);
  and (_14635_, _11215_, _07211_);
  or (_14636_, _14635_, _07209_);
  or (_14637_, _14636_, _14634_);
  nor (_14638_, _05919_, _05550_);
  nor (_14639_, _14638_, _07232_);
  and (_14640_, _14639_, _14637_);
  and (_14641_, _14622_, _07232_);
  or (_14642_, _14641_, _07230_);
  or (_14643_, _14642_, _14640_);
  nand (_14644_, _11216_, _07230_);
  and (_14645_, _14644_, _05916_);
  and (_14646_, _14645_, _14643_);
  nor (_14647_, _14646_, _14508_);
  nor (_14648_, _14647_, _06690_);
  not (_14649_, _06690_);
  nor (_14650_, _14515_, _14649_);
  or (_14651_, _14650_, _06660_);
  or (_14652_, _14651_, _14648_);
  nand (_14653_, _14515_, _06660_);
  and (_14654_, _14653_, _07051_);
  and (_14655_, _14654_, _14652_);
  nor (_14656_, _14515_, _07051_);
  or (_14657_, _14656_, _07238_);
  or (_14658_, _14657_, _14655_);
  nand (_14659_, _14515_, _07238_);
  and (_14660_, _14659_, _14658_);
  and (_14661_, _14660_, _14507_);
  nor (_14662_, _14501_, _14507_);
  or (_14663_, _14662_, _14661_);
  and (_14664_, _14663_, _14505_);
  nor (_14665_, _14501_, _14505_);
  or (_14666_, _14665_, _07242_);
  or (_14667_, _14666_, _14664_);
  and (_14668_, _14667_, _14504_);
  or (_14669_, _14668_, _06378_);
  nand (_14670_, _06378_, _05978_);
  and (_14671_, _14670_, _05913_);
  and (_14672_, _14671_, _14669_);
  and (_14673_, _05912_, _05550_);
  or (_14674_, _07249_, _14673_);
  or (_14675_, _14674_, _14672_);
  or (_14676_, _14513_, _07265_);
  not (_14677_, _07433_);
  and (_14678_, _07055_, _14677_);
  and (_14679_, _14678_, _07457_);
  and (_14680_, _14679_, _14676_);
  and (_14681_, _14680_, _14675_);
  and (_14682_, _14501_, _07456_);
  and (_14683_, _14515_, _09372_);
  or (_14684_, _14683_, _06976_);
  or (_14685_, _14684_, _14682_);
  or (_14686_, _14685_, _14681_);
  and (_14687_, _14686_, _14502_);
  or (_14688_, _14687_, _06190_);
  or (_14689_, _14503_, _14321_);
  and (_14690_, _14689_, _07507_);
  and (_14691_, _14690_, _14688_);
  or (_14692_, _14691_, _14320_);
  and (_14693_, _14692_, _14499_);
  nand (_14694_, _12275_, _06378_);
  or (_14695_, _12133_, _06378_);
  and (_14696_, _14695_, _14694_);
  and (_14697_, _14696_, _07844_);
  and (_14698_, _14697_, _14492_);
  or (_41220_, _14698_, _14693_);
  or (_14699_, _14313_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_14700_, _14699_, _14318_);
  nor (_14701_, _06019_, _05916_);
  nand (_14702_, _12797_, _12775_);
  nand (_14703_, _07931_, _10854_);
  and (_14704_, _14703_, _06243_);
  and (_14705_, _14704_, _14702_);
  nor (_14706_, _12797_, _07931_);
  or (_14707_, _14706_, _08697_);
  or (_14708_, _14702_, _08520_);
  and (_14709_, _08396_, _08301_);
  and (_14710_, _14709_, _08677_);
  nor (_14711_, _08678_, _08396_);
  or (_14712_, _14711_, _14710_);
  and (_14713_, _14712_, _06253_);
  and (_14714_, _08565_, _07578_);
  nor (_14715_, _08565_, _07578_);
  or (_14716_, _14715_, _14714_);
  or (_14717_, _14716_, _08573_);
  nor (_14718_, _06705_, _10165_);
  and (_14719_, _06705_, _06018_);
  or (_14720_, _14719_, _14718_);
  nor (_14721_, _14720_, _08572_);
  nor (_14722_, _14721_, _06253_);
  and (_14723_, _14722_, _14717_);
  or (_14724_, _14723_, _07139_);
  or (_14725_, _14724_, _14713_);
  and (_14726_, _14725_, _14708_);
  or (_14727_, _14726_, _07474_);
  nor (_14728_, _06018_, _05950_);
  nor (_14729_, _14728_, _07143_);
  and (_14730_, _14729_, _14727_);
  and (_14731_, _09380_, _07143_);
  or (_14732_, _14731_, _07159_);
  or (_14733_, _14732_, _14730_);
  and (_14734_, _14733_, _14707_);
  or (_14735_, _14734_, _06247_);
  nand (_14736_, _08396_, _06247_);
  and (_14737_, _14736_, _07270_);
  and (_14738_, _14737_, _14735_);
  not (_14739_, _12798_);
  and (_14740_, _14702_, _14739_);
  and (_14741_, _14740_, _07165_);
  or (_14742_, _14741_, _14738_);
  and (_14743_, _14742_, _05947_);
  or (_14744_, _06019_, _05947_);
  nand (_14745_, _06497_, _14744_);
  or (_14746_, _14745_, _14743_);
  nand (_14747_, _08396_, _06498_);
  and (_14748_, _14747_, _14746_);
  or (_14749_, _14748_, _07174_);
  nand (_14750_, _09251_, _07904_);
  nand (_14751_, _14750_, _08394_);
  or (_14752_, _14751_, _07369_);
  and (_14753_, _14752_, _08724_);
  and (_14754_, _14753_, _14749_);
  or (_14755_, _14754_, _14705_);
  and (_14756_, _14755_, _08723_);
  and (_14757_, _06018_, _05970_);
  or (_14758_, _07189_, _14757_);
  or (_14759_, _14758_, _14756_);
  nand (_14760_, _07578_, _07189_);
  and (_14761_, _14760_, _14759_);
  or (_14762_, _14761_, _07184_);
  or (_14763_, _09251_, _07185_);
  and (_14764_, _14763_, _08735_);
  and (_14765_, _14764_, _14762_);
  nor (_14766_, _08770_, _07578_);
  and (_14767_, _08903_, \oc8051_golden_model_1.P1 [2]);
  and (_14768_, _08894_, \oc8051_golden_model_1.PSW [2]);
  or (_14769_, _14768_, _14767_);
  and (_14770_, _08900_, \oc8051_golden_model_1.TCON [2]);
  and (_14771_, _08875_, \oc8051_golden_model_1.TL0 [2]);
  or (_14772_, _14771_, _14770_);
  or (_14773_, _14772_, _14769_);
  and (_14774_, _08912_, \oc8051_golden_model_1.TMOD [2]);
  and (_14775_, _08890_, \oc8051_golden_model_1.ACC [2]);
  or (_14776_, _14775_, _14774_);
  and (_14777_, _08930_, \oc8051_golden_model_1.SCON [2]);
  and (_14778_, _08884_, \oc8051_golden_model_1.B [2]);
  or (_14779_, _14778_, _14777_);
  or (_14780_, _14779_, _14776_);
  and (_14781_, _08924_, \oc8051_golden_model_1.P2 [2]);
  and (_14782_, _08926_, \oc8051_golden_model_1.IE [2]);
  or (_14783_, _14782_, _14781_);
  and (_14784_, _08917_, \oc8051_golden_model_1.P3 [2]);
  and (_14785_, _08919_, \oc8051_golden_model_1.IP [2]);
  or (_14786_, _14785_, _14784_);
  or (_14787_, _14786_, _14783_);
  and (_14788_, _08906_, \oc8051_golden_model_1.P0 [2]);
  and (_14789_, _08932_, \oc8051_golden_model_1.SBUF [2]);
  or (_14790_, _14789_, _14788_);
  or (_14791_, _14790_, _14787_);
  or (_14792_, _14791_, _14780_);
  or (_14793_, _14792_, _14773_);
  and (_14794_, _08940_, \oc8051_golden_model_1.TL1 [2]);
  and (_14795_, _08953_, \oc8051_golden_model_1.TH0 [2]);
  and (_14796_, _08960_, \oc8051_golden_model_1.SP [2]);
  or (_14797_, _14796_, _14795_);
  or (_14798_, _14797_, _14794_);
  and (_14799_, _08943_, \oc8051_golden_model_1.DPL [2]);
  and (_14800_, _08958_, \oc8051_golden_model_1.DPH [2]);
  or (_14801_, _14800_, _14799_);
  and (_14802_, _08947_, \oc8051_golden_model_1.PCON [2]);
  and (_14803_, _08955_, \oc8051_golden_model_1.TH1 [2]);
  or (_14804_, _14803_, _14802_);
  or (_14805_, _14804_, _14801_);
  or (_14806_, _14805_, _14798_);
  or (_14807_, _14806_, _14793_);
  or (_14808_, _14807_, _14766_);
  and (_14809_, _14808_, _07186_);
  or (_14810_, _14809_, _08973_);
  or (_14811_, _14810_, _14765_);
  and (_14812_, _08973_, _06750_);
  nor (_14813_, _14812_, _07199_);
  and (_14814_, _14813_, _14811_);
  and (_14815_, _07199_, _08945_);
  or (_14816_, _14815_, _05895_);
  or (_14817_, _14816_, _14814_);
  and (_14818_, _06019_, _05895_);
  nor (_14819_, _14818_, _07219_);
  and (_14820_, _14819_, _14817_);
  nand (_14821_, _08396_, _06651_);
  nor (_14822_, _08396_, _06651_);
  not (_14823_, _14822_);
  and (_14824_, _14823_, _14821_);
  and (_14825_, _14824_, _07219_);
  or (_14826_, _14825_, _14820_);
  and (_14827_, _14826_, _08511_);
  and (_14828_, _11214_, _07217_);
  or (_14829_, _14828_, _14827_);
  and (_14830_, _14829_, _07215_);
  and (_14831_, _14822_, _07214_);
  or (_14832_, _14831_, _14830_);
  and (_14833_, _14832_, _07212_);
  and (_14834_, _11212_, _07211_);
  or (_14835_, _14834_, _07209_);
  or (_14836_, _14835_, _14833_);
  nor (_14837_, _06018_, _05919_);
  nor (_14838_, _14837_, _07232_);
  and (_14839_, _14838_, _14836_);
  and (_14840_, _14821_, _07232_);
  or (_14841_, _14840_, _07230_);
  or (_14842_, _14841_, _14839_);
  nand (_14843_, _11213_, _07230_);
  and (_14844_, _14843_, _05916_);
  and (_14845_, _14844_, _14842_);
  or (_14846_, _14845_, _14701_);
  and (_14847_, _14846_, _12983_);
  not (_14848_, _12983_);
  and (_14849_, _14716_, _14848_);
  or (_14850_, _14849_, _07243_);
  or (_14851_, _14850_, _14847_);
  nor (_14852_, _09343_, _09252_);
  or (_14853_, _09344_, _07403_);
  or (_14854_, _14853_, _14852_);
  and (_14855_, _14854_, _09021_);
  and (_14856_, _14855_, _14851_);
  and (_14857_, _14712_, _07242_);
  or (_14858_, _14857_, _06378_);
  or (_14859_, _14858_, _14856_);
  nand (_14860_, _12309_, _06378_);
  and (_14861_, _14860_, _05913_);
  and (_14862_, _14861_, _14859_);
  and (_14863_, _06018_, _05912_);
  or (_14864_, _07249_, _14863_);
  or (_14865_, _14864_, _14862_);
  or (_14866_, _14706_, _07265_);
  and (_14867_, _14866_, _09371_);
  and (_14868_, _14867_, _14865_);
  nor (_14869_, _09382_, _09380_);
  nor (_14870_, _14869_, _09383_);
  and (_14871_, _14870_, _09372_);
  or (_14872_, _14871_, _07456_);
  or (_14873_, _14872_, _14868_);
  not (_14874_, _07456_);
  nor (_14875_, _09394_, _09251_);
  nor (_14876_, _14875_, _09395_);
  or (_14877_, _14876_, _14874_);
  and (_14878_, _14877_, _14500_);
  and (_14879_, _14878_, _14873_);
  and (_14880_, _14876_, _06976_);
  or (_14881_, _14880_, _06190_);
  or (_14882_, _14881_, _14879_);
  nor (_14883_, _08397_, _08352_);
  nor (_14884_, _14883_, _08398_);
  or (_14885_, _14884_, _14321_);
  and (_14886_, _14885_, _07507_);
  and (_14887_, _14886_, _14882_);
  or (_14888_, _14887_, _14320_);
  and (_14889_, _14888_, _14700_);
  nand (_14890_, _12269_, _06378_);
  or (_14891_, _12127_, _06378_);
  and (_14892_, _14891_, _14890_);
  and (_14893_, _14892_, _07844_);
  and (_14894_, _14893_, _14492_);
  or (_41221_, _14894_, _14889_);
  or (_14895_, _14313_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_14896_, _14895_, _14318_);
  nor (_14897_, _14710_, _08256_);
  or (_14898_, _14897_, _08680_);
  or (_14899_, _14898_, _09021_);
  nor (_14900_, _14714_, _07713_);
  or (_14901_, _14900_, _08566_);
  or (_14902_, _14901_, _09012_);
  nand (_14903_, _06095_, _05895_);
  nor (_14904_, _12925_, _08150_);
  or (_14905_, _14904_, _08697_);
  nand (_14906_, _12925_, _12903_);
  or (_14907_, _14906_, _08520_);
  and (_14908_, _14898_, _06253_);
  or (_14909_, _14901_, _08573_);
  and (_14910_, _06705_, _06075_);
  nor (_14911_, _06705_, _10218_);
  or (_14912_, _14911_, _14910_);
  nor (_14913_, _14912_, _08572_);
  nor (_14914_, _14913_, _06253_);
  and (_14915_, _14914_, _14909_);
  or (_14916_, _14915_, _07139_);
  or (_14917_, _14916_, _14908_);
  and (_14918_, _14917_, _14907_);
  or (_14919_, _14918_, _07474_);
  nor (_14920_, _06075_, _05950_);
  nor (_14921_, _14920_, _07143_);
  and (_14922_, _14921_, _14919_);
  and (_14923_, _09379_, _07143_);
  or (_14924_, _14923_, _07159_);
  or (_14925_, _14924_, _14922_);
  and (_14926_, _14925_, _14905_);
  or (_14927_, _14926_, _06247_);
  nand (_14928_, _08256_, _06247_);
  and (_14929_, _14928_, _07270_);
  and (_14930_, _14929_, _14927_);
  not (_14931_, _12926_);
  and (_14932_, _14906_, _14931_);
  and (_14933_, _14932_, _07165_);
  or (_14934_, _14933_, _14930_);
  and (_14935_, _14934_, _05947_);
  or (_14936_, _06095_, _05947_);
  nand (_14937_, _06497_, _14936_);
  or (_14938_, _14937_, _14935_);
  nand (_14939_, _08256_, _06498_);
  and (_14940_, _14939_, _14938_);
  or (_14941_, _14940_, _07174_);
  nand (_14942_, _09205_, _07904_);
  nand (_14943_, _14942_, _08254_);
  or (_14944_, _14943_, _07369_);
  and (_14945_, _14944_, _08724_);
  and (_14946_, _14945_, _14941_);
  nand (_14947_, _08150_, _10854_);
  and (_14948_, _14947_, _06243_);
  and (_14949_, _14948_, _14906_);
  or (_14950_, _14949_, _05970_);
  or (_14951_, _14950_, _14946_);
  and (_14952_, _06095_, _05970_);
  nor (_14953_, _14952_, _07189_);
  and (_14954_, _14953_, _14951_);
  nor (_14955_, _07713_, _08512_);
  or (_14956_, _14955_, _07184_);
  or (_14957_, _14956_, _14954_);
  or (_14958_, _09205_, _07185_);
  and (_14959_, _14958_, _08735_);
  and (_14960_, _14959_, _14957_);
  nor (_14961_, _08770_, _07713_);
  and (_14962_, _08903_, \oc8051_golden_model_1.P1 [3]);
  and (_14963_, _08930_, \oc8051_golden_model_1.SCON [3]);
  or (_14964_, _14963_, _14962_);
  and (_14965_, _08912_, \oc8051_golden_model_1.TMOD [3]);
  and (_14966_, _08932_, \oc8051_golden_model_1.SBUF [3]);
  or (_14967_, _14966_, _14965_);
  or (_14968_, _14967_, _14964_);
  and (_14969_, _08906_, \oc8051_golden_model_1.P0 [3]);
  and (_14970_, _08875_, \oc8051_golden_model_1.TL0 [3]);
  or (_14971_, _14970_, _14969_);
  and (_14972_, _08900_, \oc8051_golden_model_1.TCON [3]);
  and (_14973_, _08894_, \oc8051_golden_model_1.PSW [3]);
  or (_14974_, _14973_, _14972_);
  or (_14975_, _14974_, _14971_);
  and (_14976_, _08890_, \oc8051_golden_model_1.ACC [3]);
  and (_14977_, _08884_, \oc8051_golden_model_1.B [3]);
  or (_14978_, _14977_, _14976_);
  and (_14979_, _08917_, \oc8051_golden_model_1.P3 [3]);
  and (_14980_, _08919_, \oc8051_golden_model_1.IP [3]);
  or (_14981_, _14980_, _14979_);
  and (_14982_, _08924_, \oc8051_golden_model_1.P2 [3]);
  and (_14983_, _08926_, \oc8051_golden_model_1.IE [3]);
  or (_14984_, _14983_, _14982_);
  or (_14985_, _14984_, _14981_);
  or (_14986_, _14985_, _14978_);
  or (_14987_, _14986_, _14975_);
  or (_14988_, _14987_, _14968_);
  and (_14989_, _08953_, \oc8051_golden_model_1.TH0 [3]);
  and (_14990_, _08947_, \oc8051_golden_model_1.PCON [3]);
  and (_14991_, _08955_, \oc8051_golden_model_1.TH1 [3]);
  or (_14992_, _14991_, _14990_);
  or (_14993_, _14992_, _14989_);
  and (_14994_, _08943_, \oc8051_golden_model_1.DPL [3]);
  and (_14995_, _08960_, \oc8051_golden_model_1.SP [3]);
  or (_14996_, _14995_, _14994_);
  and (_14997_, _08940_, \oc8051_golden_model_1.TL1 [3]);
  and (_14998_, _08958_, \oc8051_golden_model_1.DPH [3]);
  or (_14999_, _14998_, _14997_);
  or (_15000_, _14999_, _14996_);
  or (_15001_, _15000_, _14993_);
  or (_15002_, _15001_, _14988_);
  or (_15003_, _15002_, _14961_);
  and (_15004_, _15003_, _07186_);
  or (_15005_, _15004_, _08973_);
  or (_15006_, _15005_, _14960_);
  and (_15007_, _08973_, _06292_);
  nor (_15008_, _15007_, _07199_);
  and (_15009_, _15008_, _15006_);
  and (_15010_, _07199_, _08872_);
  or (_15011_, _15010_, _05895_);
  or (_15012_, _15011_, _15009_);
  and (_15013_, _15012_, _14903_);
  or (_15014_, _15013_, _07219_);
  nand (_15015_, _08256_, _06458_);
  nor (_15016_, _08256_, _06458_);
  not (_15017_, _15016_);
  and (_15018_, _15017_, _15015_);
  or (_15019_, _15018_, _14439_);
  and (_15020_, _15019_, _08511_);
  and (_15021_, _15020_, _15014_);
  and (_15022_, _12523_, _07217_);
  or (_15023_, _15022_, _07214_);
  or (_15024_, _15023_, _15021_);
  or (_15025_, _15016_, _07215_);
  and (_15026_, _15025_, _07212_);
  and (_15027_, _15026_, _15024_);
  and (_15028_, _11210_, _07211_);
  or (_15029_, _15028_, _07209_);
  or (_15030_, _15029_, _15027_);
  nor (_15031_, _06075_, _05919_);
  nor (_15032_, _15031_, _07232_);
  and (_15033_, _15032_, _15030_);
  and (_15034_, _15015_, _07232_);
  or (_15035_, _15034_, _07230_);
  or (_15036_, _15035_, _15033_);
  nand (_15037_, _11211_, _07230_);
  and (_15038_, _15037_, _05916_);
  and (_15039_, _15038_, _15036_);
  or (_15040_, _06095_, _05916_);
  nand (_15041_, _09012_, _15040_);
  or (_15042_, _15041_, _15039_);
  and (_15043_, _15042_, _14902_);
  or (_15044_, _15043_, _07238_);
  or (_15045_, _14901_, _07463_);
  and (_15046_, _15045_, _07403_);
  and (_15047_, _15046_, _15044_);
  nor (_15048_, _09344_, _09206_);
  or (_15049_, _15048_, _09345_);
  and (_15050_, _15049_, _07243_);
  or (_15051_, _15050_, _07242_);
  or (_15052_, _15051_, _15047_);
  and (_15053_, _15052_, _14899_);
  or (_15054_, _15053_, _06378_);
  nand (_15055_, _12304_, _06378_);
  and (_15056_, _15055_, _05913_);
  and (_15057_, _15056_, _15054_);
  and (_15058_, _06075_, _05912_);
  or (_15059_, _07249_, _15058_);
  or (_15060_, _15059_, _15057_);
  or (_15061_, _14904_, _07265_);
  and (_15062_, _15061_, _09371_);
  and (_15063_, _15062_, _15060_);
  nor (_15064_, _09383_, _09379_);
  nor (_15065_, _15064_, _09384_);
  and (_15066_, _15065_, _09372_);
  or (_15067_, _15066_, _07259_);
  or (_15068_, _15067_, _15063_);
  nor (_15069_, _09395_, _09205_);
  nor (_15070_, _15069_, _09396_);
  or (_15071_, _15070_, _07414_);
  and (_15072_, _15071_, _15068_);
  or (_15073_, _15072_, _06190_);
  nor (_15074_, _08398_, _08257_);
  nor (_15075_, _15074_, _08399_);
  or (_15076_, _15075_, _14321_);
  and (_15077_, _15076_, _07507_);
  and (_15078_, _15077_, _15073_);
  or (_15079_, _15078_, _14320_);
  and (_15080_, _15079_, _14896_);
  nand (_15081_, _12264_, _06378_);
  or (_15082_, _12122_, _06378_);
  and (_15083_, _15082_, _15081_);
  and (_15084_, _15083_, _07844_);
  and (_15085_, _15084_, _14492_);
  or (_41222_, _15085_, _15080_);
  or (_15086_, _14313_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_15087_, _15086_, _14318_);
  nor (_15088_, _12154_, _05916_);
  nor (_15089_, _12846_, _12845_);
  or (_15090_, _15089_, _08697_);
  nand (_15091_, _12847_, _12845_);
  or (_15092_, _15091_, _08520_);
  and (_15093_, _08566_, _08494_);
  nor (_15094_, _08566_, _08494_);
  or (_15095_, _15094_, _15093_);
  or (_15096_, _15095_, _08573_);
  and (_15097_, _12153_, _06705_);
  nor (_15098_, _06705_, _10087_);
  or (_15099_, _15098_, _15097_);
  or (_15100_, _15099_, _08572_);
  and (_15101_, _15100_, _15096_);
  or (_15102_, _15101_, _07134_);
  or (_15103_, _09159_, _07338_);
  and (_15104_, _15103_, _15102_);
  or (_15105_, _15104_, _06253_);
  and (_15106_, _08680_, _08496_);
  nor (_15107_, _08680_, _08496_);
  or (_15108_, _15107_, _15106_);
  or (_15109_, _15108_, _08675_);
  and (_15110_, _15109_, _15105_);
  or (_15111_, _15110_, _07139_);
  and (_15112_, _15111_, _15092_);
  or (_15113_, _15112_, _07474_);
  nor (_15114_, _12153_, _05950_);
  nor (_15115_, _15114_, _07143_);
  and (_15116_, _15115_, _15113_);
  and (_15117_, _09378_, _07143_);
  or (_15118_, _15117_, _07159_);
  or (_15119_, _15118_, _15116_);
  and (_15120_, _15119_, _15090_);
  or (_15121_, _15120_, _06247_);
  nand (_15122_, _08496_, _06247_);
  and (_15123_, _15122_, _07270_);
  and (_15124_, _15123_, _15121_);
  not (_15125_, _12848_);
  and (_15126_, _15091_, _15125_);
  and (_15127_, _15126_, _07165_);
  or (_15128_, _15127_, _15124_);
  and (_15129_, _15128_, _05947_);
  or (_15130_, _12154_, _05947_);
  nand (_15131_, _15130_, _06497_);
  or (_15132_, _15131_, _15129_);
  nand (_15133_, _08496_, _06498_);
  and (_15134_, _15133_, _15132_);
  or (_15135_, _15134_, _07174_);
  and (_15136_, _09159_, _07904_);
  nand (_15137_, _08441_, _07174_);
  or (_15138_, _15137_, _15136_);
  and (_15139_, _15138_, _08724_);
  and (_15140_, _15139_, _15135_);
  nand (_15141_, _12846_, _10854_);
  and (_15142_, _15141_, _06243_);
  and (_15143_, _15142_, _15091_);
  or (_15144_, _15143_, _05970_);
  or (_15146_, _15144_, _15140_);
  and (_15147_, _12154_, _05970_);
  nor (_15148_, _15147_, _07189_);
  and (_15149_, _15148_, _15146_);
  nor (_15150_, _08494_, _08512_);
  or (_15151_, _15150_, _07184_);
  or (_15152_, _15151_, _15149_);
  or (_15153_, _09159_, _07185_);
  and (_15154_, _15153_, _08735_);
  and (_15155_, _15154_, _15152_);
  nor (_15156_, _08770_, _08494_);
  and (_15157_, _08884_, \oc8051_golden_model_1.B [4]);
  and (_15158_, _08894_, \oc8051_golden_model_1.PSW [4]);
  or (_15159_, _15158_, _15157_);
  and (_15160_, _08903_, \oc8051_golden_model_1.P1 [4]);
  and (_15161_, _08932_, \oc8051_golden_model_1.SBUF [4]);
  or (_15162_, _15161_, _15160_);
  or (_15163_, _15162_, _15159_);
  and (_15164_, _08930_, \oc8051_golden_model_1.SCON [4]);
  and (_15165_, _08890_, \oc8051_golden_model_1.ACC [4]);
  or (_15166_, _15165_, _15164_);
  and (_15167_, _08906_, \oc8051_golden_model_1.P0 [4]);
  and (_15168_, _08875_, \oc8051_golden_model_1.TL0 [4]);
  or (_15169_, _15168_, _15167_);
  or (_15170_, _15169_, _15166_);
  and (_15171_, _08900_, \oc8051_golden_model_1.TCON [4]);
  and (_15172_, _08912_, \oc8051_golden_model_1.TMOD [4]);
  or (_15173_, _15172_, _15171_);
  and (_15174_, _08924_, \oc8051_golden_model_1.P2 [4]);
  and (_15175_, _08919_, \oc8051_golden_model_1.IP [4]);
  or (_15176_, _15175_, _15174_);
  and (_15177_, _08926_, \oc8051_golden_model_1.IE [4]);
  and (_15178_, _08917_, \oc8051_golden_model_1.P3 [4]);
  or (_15179_, _15178_, _15177_);
  or (_15180_, _15179_, _15176_);
  or (_15181_, _15180_, _15173_);
  or (_15182_, _15181_, _15170_);
  or (_15183_, _15182_, _15163_);
  and (_15184_, _08955_, \oc8051_golden_model_1.TH1 [4]);
  and (_15185_, _08953_, \oc8051_golden_model_1.TH0 [4]);
  and (_15186_, _08940_, \oc8051_golden_model_1.TL1 [4]);
  or (_15187_, _15186_, _15185_);
  or (_15188_, _15187_, _15184_);
  and (_15189_, _08943_, \oc8051_golden_model_1.DPL [4]);
  and (_15190_, _08947_, \oc8051_golden_model_1.PCON [4]);
  or (_15191_, _15190_, _15189_);
  and (_15192_, _08960_, \oc8051_golden_model_1.SP [4]);
  and (_15193_, _08958_, \oc8051_golden_model_1.DPH [4]);
  or (_15194_, _15193_, _15192_);
  or (_15195_, _15194_, _15191_);
  or (_15196_, _15195_, _15188_);
  or (_15197_, _15196_, _15183_);
  or (_15198_, _15197_, _15156_);
  and (_15199_, _15198_, _07186_);
  or (_15200_, _15199_, _08973_);
  or (_15201_, _15200_, _15155_);
  and (_15202_, _08973_, _06230_);
  nor (_15203_, _15202_, _07199_);
  and (_15204_, _15203_, _15201_);
  and (_15205_, _08892_, _07199_);
  or (_15206_, _15205_, _05895_);
  or (_15207_, _15206_, _15204_);
  and (_15208_, _12154_, _05895_);
  nor (_15209_, _15208_, _07219_);
  and (_15210_, _15209_, _15207_);
  nand (_15211_, _08834_, _08496_);
  nor (_15212_, _08834_, _08496_);
  not (_15213_, _15212_);
  and (_15214_, _15213_, _15211_);
  and (_15215_, _15214_, _07219_);
  or (_15216_, _15215_, _15210_);
  and (_15217_, _15216_, _08511_);
  and (_15218_, _11209_, _07217_);
  or (_15219_, _15218_, _07214_);
  or (_15220_, _15219_, _15217_);
  or (_15221_, _15212_, _07215_);
  and (_15222_, _15221_, _07212_);
  and (_15223_, _15222_, _15220_);
  and (_15224_, _11206_, _07211_);
  or (_15225_, _15224_, _07209_);
  or (_15226_, _15225_, _15223_);
  nor (_15227_, _12153_, _05919_);
  nor (_15228_, _15227_, _07232_);
  and (_15229_, _15228_, _15226_);
  and (_15230_, _15211_, _07232_);
  or (_15231_, _15230_, _07230_);
  or (_15232_, _15231_, _15229_);
  nand (_15233_, _11208_, _07230_);
  and (_15234_, _15233_, _05916_);
  and (_15235_, _15234_, _15232_);
  or (_15236_, _15235_, _15088_);
  and (_15237_, _15236_, _09012_);
  not (_15238_, _09012_);
  and (_15239_, _15095_, _15238_);
  or (_15240_, _15239_, _07238_);
  or (_15241_, _15240_, _15237_);
  nor (_15242_, _07238_, _14506_);
  and (_15243_, _15095_, _14507_);
  or (_15244_, _15243_, _15242_);
  and (_15245_, _15244_, _15241_);
  nor (_15246_, _09345_, _09160_);
  or (_15247_, _15246_, _09346_);
  or (_15248_, _15247_, _06963_);
  and (_15249_, _15248_, _07243_);
  or (_15250_, _15249_, _15245_);
  or (_15251_, _15247_, _14505_);
  and (_15252_, _15251_, _09021_);
  and (_15253_, _15252_, _15250_);
  and (_15254_, _15108_, _07242_);
  or (_15255_, _15254_, _06378_);
  or (_15256_, _15255_, _15253_);
  nand (_15257_, _12300_, _06378_);
  and (_15258_, _15257_, _05913_);
  and (_15259_, _15258_, _15256_);
  and (_15260_, _12153_, _05912_);
  or (_15261_, _15260_, _07249_);
  or (_15262_, _15261_, _15259_);
  or (_15263_, _15089_, _07265_);
  and (_15264_, _15263_, _09371_);
  and (_15265_, _15264_, _15262_);
  nor (_15266_, _09384_, _09378_);
  nor (_15267_, _15266_, _09385_);
  and (_15268_, _15267_, _09372_);
  or (_15269_, _15268_, _07456_);
  or (_15270_, _15269_, _15265_);
  nor (_15271_, _09396_, _09159_);
  nor (_15272_, _15271_, _09397_);
  or (_15273_, _15272_, _14874_);
  and (_15274_, _15273_, _14500_);
  and (_15275_, _15274_, _15270_);
  and (_15276_, _15272_, _06976_);
  or (_15277_, _15276_, _06190_);
  or (_15278_, _15277_, _15275_);
  nor (_15279_, _08497_, _08399_);
  nor (_15280_, _15279_, _08498_);
  or (_15281_, _15280_, _14321_);
  and (_15282_, _15281_, _07507_);
  and (_15283_, _15282_, _15278_);
  or (_15284_, _15283_, _14320_);
  and (_15285_, _15284_, _15087_);
  nand (_15286_, _12259_, _06378_);
  or (_15287_, _12117_, _06378_);
  and (_15288_, _15287_, _15286_);
  and (_15289_, _15288_, _07844_);
  and (_15290_, _15289_, _14492_);
  or (_41223_, _15290_, _15285_);
  or (_15291_, _14313_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_15292_, _15291_, _14318_);
  nor (_15293_, _12149_, _05916_);
  nor (_15294_, _12949_, _12948_);
  or (_15295_, _15294_, _08697_);
  nand (_15296_, _12950_, _12948_);
  or (_15297_, _15296_, _08520_);
  or (_15298_, _09113_, _07338_);
  nor (_15299_, _15093_, _08209_);
  or (_15300_, _15299_, _08567_);
  and (_15301_, _15300_, _08572_);
  nor (_15302_, _06705_, _10122_);
  and (_15303_, _12148_, _06705_);
  or (_15304_, _15303_, _15302_);
  and (_15305_, _15304_, _08573_);
  or (_15306_, _15305_, _07134_);
  or (_15307_, _15306_, _15301_);
  and (_15308_, _15307_, _15298_);
  or (_15309_, _15308_, _06253_);
  nor (_15310_, _15106_, _08211_);
  or (_15311_, _15310_, _08681_);
  or (_15312_, _15311_, _08675_);
  and (_15313_, _15312_, _15309_);
  or (_15314_, _15313_, _07139_);
  and (_15315_, _15314_, _15297_);
  or (_15316_, _15315_, _07474_);
  nor (_15317_, _12148_, _05950_);
  nor (_15318_, _15317_, _07143_);
  and (_15319_, _15318_, _15316_);
  and (_15320_, _09377_, _07143_);
  or (_15321_, _15320_, _07159_);
  or (_15322_, _15321_, _15319_);
  and (_15323_, _15322_, _15295_);
  or (_15324_, _15323_, _06247_);
  nand (_15325_, _08211_, _06247_);
  and (_15326_, _15325_, _07270_);
  and (_15327_, _15326_, _15324_);
  not (_15328_, _12951_);
  and (_15329_, _15296_, _07165_);
  and (_15330_, _15329_, _15328_);
  or (_15331_, _15330_, _15327_);
  and (_15332_, _15331_, _05947_);
  or (_15333_, _12149_, _05947_);
  nand (_15334_, _15333_, _06497_);
  or (_15335_, _15334_, _15332_);
  nand (_15336_, _08211_, _06498_);
  and (_15337_, _15336_, _15335_);
  or (_15338_, _15337_, _07174_);
  and (_15339_, _09113_, _07904_);
  nand (_15340_, _08156_, _07174_);
  or (_15341_, _15340_, _15339_);
  and (_15342_, _15341_, _08724_);
  and (_15343_, _15342_, _15338_);
  nand (_15344_, _12949_, _10854_);
  and (_15345_, _15344_, _06243_);
  and (_15346_, _15345_, _15296_);
  or (_15347_, _15346_, _05970_);
  or (_15348_, _15347_, _15343_);
  and (_15349_, _12149_, _05970_);
  nor (_15350_, _15349_, _07189_);
  and (_15351_, _15350_, _15348_);
  nor (_15352_, _08209_, _08512_);
  or (_15353_, _15352_, _07184_);
  or (_15354_, _15353_, _15351_);
  or (_15355_, _09113_, _07185_);
  and (_15356_, _15355_, _08735_);
  and (_15357_, _15356_, _15354_);
  nor (_15358_, _08770_, _08209_);
  and (_15359_, _08903_, \oc8051_golden_model_1.P1 [5]);
  and (_15360_, _08884_, \oc8051_golden_model_1.B [5]);
  or (_15361_, _15360_, _15359_);
  and (_15362_, _08906_, \oc8051_golden_model_1.P0 [5]);
  and (_15363_, _08890_, \oc8051_golden_model_1.ACC [5]);
  or (_15364_, _15363_, _15362_);
  or (_15365_, _15364_, _15361_);
  and (_15366_, _08900_, \oc8051_golden_model_1.TCON [5]);
  and (_15367_, _08912_, \oc8051_golden_model_1.TMOD [5]);
  or (_15368_, _15367_, _15366_);
  and (_15369_, _08875_, \oc8051_golden_model_1.TL0 [5]);
  and (_15370_, _08930_, \oc8051_golden_model_1.SCON [5]);
  or (_15371_, _15370_, _15369_);
  or (_15372_, _15371_, _15368_);
  and (_15373_, _08924_, \oc8051_golden_model_1.P2 [5]);
  and (_15374_, _08917_, \oc8051_golden_model_1.P3 [5]);
  or (_15375_, _15374_, _15373_);
  and (_15376_, _08926_, \oc8051_golden_model_1.IE [5]);
  and (_15377_, _08919_, \oc8051_golden_model_1.IP [5]);
  or (_15378_, _15377_, _15376_);
  or (_15379_, _15378_, _15375_);
  and (_15380_, _08932_, \oc8051_golden_model_1.SBUF [5]);
  and (_15381_, _08894_, \oc8051_golden_model_1.PSW [5]);
  or (_15382_, _15381_, _15380_);
  or (_15383_, _15382_, _15379_);
  or (_15384_, _15383_, _15372_);
  or (_15385_, _15384_, _15365_);
  and (_15386_, _08960_, \oc8051_golden_model_1.SP [5]);
  and (_15387_, _08943_, \oc8051_golden_model_1.DPL [5]);
  and (_15388_, _08955_, \oc8051_golden_model_1.TH1 [5]);
  or (_15389_, _15388_, _15387_);
  or (_15390_, _15389_, _15386_);
  and (_15391_, _08940_, \oc8051_golden_model_1.TL1 [5]);
  and (_15392_, _08958_, \oc8051_golden_model_1.DPH [5]);
  or (_15393_, _15392_, _15391_);
  and (_15394_, _08947_, \oc8051_golden_model_1.PCON [5]);
  and (_15395_, _08953_, \oc8051_golden_model_1.TH0 [5]);
  or (_15396_, _15395_, _15394_);
  or (_15397_, _15396_, _15393_);
  or (_15398_, _15397_, _15390_);
  or (_15399_, _15398_, _15385_);
  or (_15400_, _15399_, _15358_);
  and (_15401_, _15400_, _07186_);
  or (_15402_, _15401_, _08973_);
  or (_15403_, _15402_, _15357_);
  and (_15404_, _08973_, _06608_);
  nor (_15405_, _15404_, _07199_);
  and (_15406_, _15405_, _15403_);
  and (_15407_, _08888_, _07199_);
  or (_15408_, _15407_, _05895_);
  or (_15409_, _15408_, _15406_);
  and (_15410_, _12149_, _05895_);
  nor (_15411_, _15410_, _07219_);
  and (_15412_, _15411_, _15409_);
  nand (_15413_, _08867_, _08211_);
  nor (_15414_, _08867_, _08211_);
  not (_15415_, _15414_);
  and (_15416_, _15415_, _15413_);
  and (_15417_, _15416_, _07219_);
  or (_15418_, _15417_, _15412_);
  and (_15419_, _15418_, _08511_);
  and (_15420_, _11205_, _07217_);
  or (_15421_, _15420_, _15419_);
  and (_15422_, _15421_, _07215_);
  and (_15423_, _15414_, _07214_);
  or (_15424_, _15423_, _15422_);
  and (_15425_, _15424_, _07212_);
  and (_15426_, _11203_, _07211_);
  or (_15427_, _15426_, _07209_);
  or (_15428_, _15427_, _15425_);
  nor (_15429_, _12148_, _05919_);
  nor (_15430_, _15429_, _07232_);
  and (_15431_, _15430_, _15428_);
  and (_15432_, _15413_, _07232_);
  or (_15433_, _15432_, _07230_);
  or (_15434_, _15433_, _15431_);
  nand (_15435_, _11204_, _07230_);
  and (_15436_, _15435_, _05916_);
  and (_15437_, _15436_, _15434_);
  or (_15438_, _15437_, _15293_);
  and (_15439_, _15438_, _09012_);
  and (_15440_, _15300_, _15238_);
  or (_15441_, _15440_, _07238_);
  or (_15442_, _15441_, _15439_);
  or (_15443_, _15300_, _07463_);
  and (_15444_, _15443_, _14507_);
  and (_15445_, _15444_, _15442_);
  nor (_15446_, _09346_, _09114_);
  or (_15447_, _15446_, _09347_);
  or (_15448_, _15447_, _06963_);
  and (_15449_, _15448_, _07243_);
  or (_15450_, _15449_, _15445_);
  or (_15451_, _15447_, _14505_);
  and (_15452_, _15451_, _09021_);
  and (_15453_, _15452_, _15450_);
  and (_15454_, _15311_, _07242_);
  or (_15455_, _15454_, _06378_);
  or (_15456_, _15455_, _15453_);
  nand (_15457_, _12295_, _06378_);
  and (_15458_, _15457_, _05913_);
  and (_15459_, _15458_, _15456_);
  and (_15460_, _12148_, _05912_);
  or (_15461_, _15460_, _07249_);
  or (_15462_, _15461_, _15459_);
  or (_15463_, _15294_, _07265_);
  and (_15464_, _15463_, _09371_);
  and (_15465_, _15464_, _15462_);
  nor (_15466_, _09385_, _09377_);
  nor (_15467_, _15466_, _09386_);
  and (_15468_, _15467_, _09372_);
  or (_15469_, _15468_, _07259_);
  or (_15470_, _15469_, _15465_);
  nor (_15471_, _09397_, _09113_);
  nor (_15472_, _15471_, _09398_);
  or (_15473_, _15472_, _07414_);
  and (_15474_, _15473_, _15470_);
  or (_15475_, _15474_, _06190_);
  nor (_15476_, _08498_, _08212_);
  nor (_15477_, _15476_, _08499_);
  or (_15478_, _15477_, _14321_);
  and (_15479_, _15478_, _07507_);
  and (_15480_, _15479_, _15475_);
  or (_15481_, _15480_, _14320_);
  and (_15482_, _15481_, _15292_);
  not (_15483_, _12113_);
  nor (_15484_, _15483_, _06378_);
  and (_15485_, _12253_, _06378_);
  or (_15486_, _15485_, _15484_);
  and (_15487_, _15486_, _07844_);
  and (_15488_, _15487_, _14492_);
  or (_41225_, _15488_, _15482_);
  or (_15489_, _14313_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_15490_, _15489_, _14318_);
  nor (_15491_, _09386_, _09376_);
  nor (_15492_, _15491_, _09387_);
  and (_15493_, _15492_, _09372_);
  nor (_15494_, _08567_, _08106_);
  or (_15495_, _15494_, _08568_);
  or (_15496_, _15495_, _09012_);
  nor (_15497_, _12899_, _12898_);
  or (_15498_, _15497_, _08697_);
  nand (_15499_, _12900_, _12898_);
  or (_15500_, _15499_, _08520_);
  or (_15501_, _15495_, _08573_);
  nor (_15502_, _06705_, _10068_);
  and (_15503_, _12141_, _06705_);
  or (_15504_, _15503_, _08572_);
  or (_15505_, _15504_, _15502_);
  and (_15506_, _15505_, _15501_);
  or (_15507_, _15506_, _07134_);
  or (_15508_, _09067_, _07338_);
  and (_15509_, _15508_, _15507_);
  or (_15510_, _15509_, _06253_);
  nor (_15511_, _08681_, _08108_);
  or (_15512_, _15511_, _08682_);
  or (_15513_, _15512_, _08675_);
  and (_15514_, _15513_, _15510_);
  or (_15515_, _15514_, _07139_);
  and (_15516_, _15515_, _15500_);
  or (_15517_, _15516_, _07474_);
  nor (_15518_, _12141_, _05950_);
  nor (_15519_, _15518_, _07143_);
  and (_15520_, _15519_, _15517_);
  and (_15521_, _09376_, _07143_);
  or (_15522_, _15521_, _07159_);
  or (_15523_, _15522_, _15520_);
  and (_15524_, _15523_, _15498_);
  or (_15525_, _15524_, _06247_);
  nand (_15526_, _08108_, _06247_);
  and (_15527_, _15526_, _07270_);
  and (_15528_, _15527_, _15525_);
  not (_15529_, _12901_);
  and (_15530_, _15499_, _15529_);
  and (_15531_, _15530_, _07165_);
  or (_15532_, _15531_, _15528_);
  and (_15533_, _15532_, _05947_);
  or (_15534_, _12142_, _05947_);
  nand (_15535_, _15534_, _06497_);
  or (_15536_, _15535_, _15533_);
  nand (_15537_, _08108_, _06498_);
  and (_15538_, _15537_, _15536_);
  or (_15539_, _15538_, _07174_);
  and (_15540_, _09067_, _07904_);
  nand (_15541_, _08053_, _07174_);
  or (_15542_, _15541_, _15540_);
  and (_15543_, _15542_, _08724_);
  and (_15544_, _15543_, _15539_);
  nand (_15545_, _12899_, _10854_);
  and (_15546_, _15545_, _06243_);
  and (_15547_, _15546_, _15499_);
  or (_15548_, _15547_, _05970_);
  or (_15549_, _15548_, _15544_);
  and (_15550_, _12142_, _05970_);
  nor (_15551_, _15550_, _07189_);
  and (_15552_, _15551_, _15549_);
  nor (_15553_, _08106_, _08512_);
  or (_15554_, _15553_, _07184_);
  or (_15555_, _15554_, _15552_);
  or (_15556_, _09067_, _07185_);
  and (_15557_, _15556_, _08735_);
  and (_15558_, _15557_, _15555_);
  nor (_15559_, _08770_, _08106_);
  and (_15560_, _08875_, \oc8051_golden_model_1.TL0 [6]);
  and (_15561_, _08884_, \oc8051_golden_model_1.B [6]);
  or (_15562_, _15561_, _15560_);
  and (_15563_, _08890_, \oc8051_golden_model_1.ACC [6]);
  and (_15564_, _08894_, \oc8051_golden_model_1.PSW [6]);
  or (_15565_, _15564_, _15563_);
  or (_15566_, _15565_, _15562_);
  and (_15567_, _08900_, \oc8051_golden_model_1.TCON [6]);
  and (_15568_, _08932_, \oc8051_golden_model_1.SBUF [6]);
  or (_15569_, _15568_, _15567_);
  and (_15570_, _08906_, \oc8051_golden_model_1.P0 [6]);
  and (_15571_, _08912_, \oc8051_golden_model_1.TMOD [6]);
  or (_15572_, _15571_, _15570_);
  or (_15573_, _15572_, _15569_);
  and (_15574_, _08924_, \oc8051_golden_model_1.P2 [6]);
  and (_15575_, _08919_, \oc8051_golden_model_1.IP [6]);
  or (_15576_, _15575_, _15574_);
  and (_15577_, _08926_, \oc8051_golden_model_1.IE [6]);
  and (_15578_, _08917_, \oc8051_golden_model_1.P3 [6]);
  or (_15579_, _15578_, _15577_);
  or (_15580_, _15579_, _15576_);
  and (_15581_, _08903_, \oc8051_golden_model_1.P1 [6]);
  and (_15582_, _08930_, \oc8051_golden_model_1.SCON [6]);
  or (_15583_, _15582_, _15581_);
  or (_15584_, _15583_, _15580_);
  or (_15585_, _15584_, _15573_);
  or (_15586_, _15585_, _15566_);
  and (_15587_, _08953_, \oc8051_golden_model_1.TH0 [6]);
  and (_15588_, _08943_, \oc8051_golden_model_1.DPL [6]);
  and (_15589_, _08958_, \oc8051_golden_model_1.DPH [6]);
  or (_15590_, _15589_, _15588_);
  or (_15591_, _15590_, _15587_);
  and (_15592_, _08940_, \oc8051_golden_model_1.TL1 [6]);
  and (_15593_, _08955_, \oc8051_golden_model_1.TH1 [6]);
  or (_15594_, _15593_, _15592_);
  and (_15595_, _08947_, \oc8051_golden_model_1.PCON [6]);
  and (_15596_, _08960_, \oc8051_golden_model_1.SP [6]);
  or (_15597_, _15596_, _15595_);
  or (_15598_, _15597_, _15594_);
  or (_15599_, _15598_, _15591_);
  or (_15600_, _15599_, _15586_);
  or (_15601_, _15600_, _15559_);
  and (_15602_, _15601_, _07186_);
  or (_15603_, _15602_, _08973_);
  or (_15604_, _15603_, _15558_);
  and (_15605_, _08973_, _06326_);
  nor (_15606_, _15605_, _07199_);
  and (_15607_, _15606_, _15604_);
  not (_15608_, _08802_);
  and (_15609_, _15608_, _07199_);
  or (_15610_, _15609_, _05895_);
  or (_15611_, _15610_, _15607_);
  and (_15612_, _12142_, _05895_);
  nor (_15613_, _15612_, _07219_);
  and (_15614_, _15613_, _15611_);
  nand (_15615_, _08802_, _08108_);
  nor (_15616_, _08802_, _08108_);
  not (_15617_, _15616_);
  and (_15618_, _15617_, _15615_);
  and (_15619_, _15618_, _07219_);
  or (_15620_, _15619_, _15614_);
  and (_15621_, _15620_, _08511_);
  and (_15622_, _11202_, _07217_);
  or (_15623_, _15622_, _15621_);
  and (_15624_, _15623_, _07215_);
  and (_15625_, _15616_, _07214_);
  or (_15626_, _15625_, _15624_);
  and (_15627_, _15626_, _07212_);
  and (_15628_, _11199_, _07211_);
  or (_15629_, _15628_, _07209_);
  or (_15630_, _15629_, _15627_);
  nor (_15631_, _12141_, _05919_);
  nor (_15632_, _15631_, _07232_);
  and (_15633_, _15632_, _15630_);
  and (_15634_, _15615_, _07232_);
  or (_15635_, _15634_, _07230_);
  or (_15636_, _15635_, _15633_);
  nand (_15637_, _11201_, _07230_);
  and (_15638_, _15637_, _05916_);
  and (_15639_, _15638_, _15636_);
  or (_15640_, _12142_, _05916_);
  nand (_15641_, _15640_, _09012_);
  or (_15642_, _15641_, _15639_);
  and (_15643_, _15642_, _15496_);
  or (_15644_, _15643_, _07238_);
  and (_15645_, _15495_, _14507_);
  or (_15646_, _15645_, _15242_);
  and (_15647_, _15646_, _15644_);
  nor (_15648_, _09347_, _09068_);
  or (_15649_, _15648_, _09348_);
  or (_15650_, _15649_, _06963_);
  and (_15651_, _15650_, _07243_);
  or (_15652_, _15651_, _15647_);
  or (_15653_, _15649_, _14505_);
  and (_15654_, _15653_, _09021_);
  and (_15655_, _15654_, _15652_);
  and (_15656_, _15512_, _07242_);
  or (_15657_, _15656_, _06378_);
  or (_15658_, _15657_, _15655_);
  nand (_15659_, _12288_, _06378_);
  and (_15660_, _15659_, _05913_);
  and (_15661_, _15660_, _15658_);
  and (_15662_, _12141_, _05912_);
  or (_15663_, _15662_, _07249_);
  or (_15664_, _15663_, _15661_);
  or (_15665_, _15497_, _07265_);
  and (_15666_, _15665_, _09371_);
  and (_15667_, _15666_, _15664_);
  or (_15668_, _15667_, _15493_);
  and (_15669_, _15668_, _07414_);
  or (_15670_, _09398_, _09067_);
  nor (_15671_, _09399_, _07414_);
  and (_15672_, _15671_, _15670_);
  or (_15673_, _15672_, _06190_);
  or (_15674_, _15673_, _15669_);
  nor (_15675_, _08499_, _08109_);
  nor (_15676_, _15675_, _08500_);
  or (_15677_, _15676_, _14321_);
  and (_15678_, _15677_, _07507_);
  and (_15679_, _15678_, _15674_);
  or (_15680_, _15679_, _14320_);
  and (_15681_, _15680_, _15490_);
  not (_15682_, _12108_);
  nor (_15683_, _15682_, _06378_);
  and (_15684_, _12248_, _06378_);
  or (_15685_, _15684_, _15683_);
  and (_15686_, _15685_, _07844_);
  and (_15687_, _15686_, _14492_);
  or (_41226_, _15687_, _15681_);
  or (_15688_, _14313_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_15689_, _15688_, _14318_);
  nand (_15690_, _14313_, _09407_);
  and (_15691_, _15690_, _15689_);
  and (_15692_, _14492_, _09446_);
  or (_41227_, _15692_, _15691_);
  and (_15693_, _07509_, _07263_);
  and (_15694_, _15693_, _14309_);
  or (_15695_, _15694_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_15696_, _14489_, _07507_);
  not (_15697_, _15696_);
  nand (_15698_, _15697_, _15694_);
  and (_15699_, _15698_, _15695_);
  and (_15700_, _07844_, _07512_);
  and (_15701_, _15700_, _14316_);
  or (_15702_, _15701_, _15699_);
  not (_15703_, _07844_);
  nand (_15704_, _14316_, _07512_);
  or (_15705_, _15704_, _15703_);
  or (_15706_, _15705_, _14495_);
  and (_41230_, _15706_, _15702_);
  not (_15707_, _15694_);
  or (_15708_, _15707_, _14691_);
  or (_15709_, _15694_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_15710_, _15709_, _15705_);
  and (_15711_, _15710_, _15708_);
  and (_15712_, _15701_, _14697_);
  or (_41233_, _15712_, _15711_);
  or (_15713_, _15707_, _14887_);
  or (_15714_, _15694_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_15715_, _15714_, _15705_);
  and (_15716_, _15715_, _15713_);
  and (_15717_, _15701_, _14893_);
  or (_41234_, _15717_, _15716_);
  or (_15718_, _15707_, _15078_);
  or (_15719_, _15694_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_15720_, _15719_, _15705_);
  and (_15721_, _15720_, _15718_);
  and (_15722_, _15701_, _15084_);
  or (_41235_, _15722_, _15721_);
  or (_15723_, _15707_, _15283_);
  or (_15724_, _15694_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_15725_, _15724_, _15705_);
  and (_15726_, _15725_, _15723_);
  and (_15727_, _15701_, _15289_);
  or (_41236_, _15727_, _15726_);
  or (_15728_, _15707_, _15480_);
  or (_15729_, _15694_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_15730_, _15729_, _15705_);
  and (_15731_, _15730_, _15728_);
  and (_15732_, _15701_, _15487_);
  or (_41237_, _15732_, _15731_);
  or (_15733_, _15707_, _15679_);
  or (_15734_, _15694_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_15735_, _15734_, _15705_);
  and (_15736_, _15735_, _15733_);
  and (_15737_, _15701_, _15686_);
  or (_41239_, _15737_, _15736_);
  or (_15738_, _15707_, _09408_);
  or (_15739_, _15694_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_15740_, _15739_, _15705_);
  and (_15741_, _15740_, _15738_);
  and (_15742_, _15701_, _09446_);
  or (_41240_, _15742_, _15741_);
  and (_15743_, _14310_, _07419_);
  and (_15744_, _15743_, _14309_);
  or (_15745_, _15744_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_15746_, _15744_, _15697_);
  and (_15747_, _15746_, _15745_);
  and (_15748_, _08588_, _07844_);
  and (_15749_, _15748_, _14316_);
  or (_15750_, _15749_, _15747_);
  nand (_15751_, _14316_, _08588_);
  or (_15752_, _15751_, _15703_);
  or (_15753_, _15752_, _14495_);
  and (_41244_, _15753_, _15750_);
  not (_15754_, _15744_);
  or (_15755_, _15754_, _14691_);
  or (_15756_, _15744_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_15757_, _15756_, _15752_);
  and (_15758_, _15757_, _15755_);
  and (_15759_, _15749_, _14697_);
  or (_41245_, _15759_, _15758_);
  or (_15760_, _15754_, _14887_);
  or (_15761_, _15744_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_15762_, _15761_, _15752_);
  and (_15763_, _15762_, _15760_);
  and (_15764_, _15749_, _14893_);
  or (_41247_, _15764_, _15763_);
  or (_15765_, _15754_, _15078_);
  or (_15766_, _15744_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_15767_, _15766_, _15752_);
  and (_15768_, _15767_, _15765_);
  and (_15769_, _15749_, _15084_);
  or (_41248_, _15769_, _15768_);
  or (_15770_, _15754_, _15283_);
  or (_15771_, _15744_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_15772_, _15771_, _15752_);
  and (_15773_, _15772_, _15770_);
  and (_15774_, _15749_, _15289_);
  or (_41249_, _15774_, _15773_);
  or (_15775_, _15754_, _15480_);
  or (_15776_, _15744_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_15777_, _15776_, _15752_);
  and (_15778_, _15777_, _15775_);
  and (_15779_, _15749_, _15487_);
  or (_41250_, _15779_, _15778_);
  or (_15780_, _15754_, _15679_);
  or (_15781_, _15744_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_15782_, _15781_, _15752_);
  and (_15783_, _15782_, _15780_);
  and (_15784_, _15749_, _15686_);
  or (_41251_, _15784_, _15783_);
  or (_15785_, _15754_, _09408_);
  or (_15786_, _15744_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_15787_, _15786_, _15752_);
  and (_15788_, _15787_, _15785_);
  and (_15789_, _15749_, _09446_);
  or (_41253_, _15789_, _15788_);
  not (_15790_, _14310_);
  nor (_15791_, _15790_, _07419_);
  and (_15792_, _14309_, _15791_);
  nor (_15793_, _15792_, _07279_);
  nand (_15794_, _14316_, _06234_);
  or (_15795_, _15794_, _15703_);
  nand (_15796_, _15792_, _15696_);
  nand (_15797_, _15796_, _15795_);
  or (_15798_, _15797_, _15793_);
  or (_15799_, _15795_, _14495_);
  and (_41255_, _15799_, _15798_);
  or (_15800_, _15792_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_15801_, _15800_, _15795_);
  not (_15802_, _15792_);
  or (_15803_, _15802_, _14691_);
  and (_15804_, _15803_, _15801_);
  and (_15805_, _07844_, _06234_);
  and (_15806_, _15805_, _14316_);
  and (_15807_, _15806_, _14697_);
  or (_41256_, _15807_, _15804_);
  or (_15808_, _15792_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_15809_, _15808_, _15795_);
  or (_15810_, _15802_, _14887_);
  and (_15811_, _15810_, _15809_);
  and (_15812_, _15806_, _14893_);
  or (_41257_, _15812_, _15811_);
  or (_15813_, _15792_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_15814_, _15813_, _15795_);
  or (_15815_, _15802_, _15078_);
  and (_15816_, _15815_, _15814_);
  and (_15817_, _15806_, _15084_);
  or (_41258_, _15817_, _15816_);
  or (_15818_, _15792_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_15819_, _15818_, _15795_);
  or (_15820_, _15802_, _15283_);
  and (_15821_, _15820_, _15819_);
  and (_15822_, _15806_, _15289_);
  or (_41259_, _15822_, _15821_);
  or (_15823_, _15792_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_15824_, _15823_, _15795_);
  or (_15825_, _15802_, _15480_);
  and (_15826_, _15825_, _15824_);
  and (_15827_, _15806_, _15487_);
  or (_41260_, _15827_, _15826_);
  or (_15828_, _15792_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_15829_, _15828_, _15795_);
  or (_15830_, _15802_, _15679_);
  and (_15831_, _15830_, _15829_);
  and (_15832_, _15806_, _15686_);
  or (_41262_, _15832_, _15831_);
  or (_15833_, _15792_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_15834_, _15833_, _15795_);
  or (_15835_, _15802_, _09408_);
  and (_15836_, _15835_, _15834_);
  and (_15837_, _15806_, _09446_);
  or (_41263_, _15837_, _15836_);
  and (_15838_, _14308_, _07830_);
  and (_15839_, _15838_, _14311_);
  nand (_15840_, _15839_, _15697_);
  not (_15841_, _07840_);
  and (_15842_, _14315_, _15841_);
  and (_15843_, _15842_, _06236_);
  not (_15844_, _15843_);
  or (_15845_, _15839_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_15846_, _15845_, _15844_);
  and (_15847_, _15846_, _15840_);
  and (_15848_, _15843_, _14496_);
  or (_41266_, _15848_, _15847_);
  not (_15849_, _15839_);
  or (_15850_, _15849_, _14691_);
  or (_15851_, _15839_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_15852_, _15851_, _15844_);
  and (_15853_, _15852_, _15850_);
  and (_15854_, _15843_, _14697_);
  or (_41267_, _15854_, _15853_);
  or (_15855_, _15849_, _14887_);
  or (_15856_, _15839_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_15857_, _15856_, _15844_);
  and (_15858_, _15857_, _15855_);
  and (_15859_, _15843_, _14893_);
  or (_41269_, _15859_, _15858_);
  or (_15860_, _15849_, _15078_);
  or (_15861_, _15839_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_15862_, _15861_, _15844_);
  and (_15863_, _15862_, _15860_);
  and (_15864_, _15843_, _15084_);
  or (_41270_, _15864_, _15863_);
  or (_15865_, _15849_, _15283_);
  or (_15866_, _15839_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_15867_, _15866_, _15844_);
  and (_15868_, _15867_, _15865_);
  and (_15869_, _15843_, _15289_);
  or (_41271_, _15869_, _15868_);
  or (_15870_, _15849_, _15480_);
  or (_15871_, _15839_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_15872_, _15871_, _15844_);
  and (_15873_, _15872_, _15870_);
  and (_15874_, _15843_, _15487_);
  or (_41272_, _15874_, _15873_);
  or (_15875_, _15849_, _15679_);
  or (_15876_, _15839_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_15877_, _15876_, _15844_);
  and (_15878_, _15877_, _15875_);
  and (_15879_, _15843_, _15686_);
  or (_41273_, _15879_, _15878_);
  or (_15880_, _15849_, _09408_);
  or (_15881_, _15839_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_15882_, _15881_, _15844_);
  and (_15883_, _15882_, _15880_);
  and (_15884_, _15843_, _09446_);
  or (_41275_, _15884_, _15883_);
  and (_15885_, _15838_, _15693_);
  nand (_15886_, _15885_, _15697_);
  and (_15887_, _15842_, _07512_);
  not (_15888_, _15887_);
  or (_15889_, _15885_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_15890_, _15889_, _15888_);
  and (_15891_, _15890_, _15886_);
  and (_15892_, _15887_, _14496_);
  or (_41277_, _15892_, _15891_);
  not (_15893_, _15885_);
  or (_15894_, _15893_, _14691_);
  or (_15895_, _15885_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_15896_, _15895_, _15888_);
  and (_15897_, _15896_, _15894_);
  and (_15898_, _15887_, _14697_);
  or (_41278_, _15898_, _15897_);
  or (_15899_, _15893_, _14887_);
  or (_15900_, _15885_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_15901_, _15900_, _15888_);
  and (_15902_, _15901_, _15899_);
  and (_15903_, _15887_, _14893_);
  or (_41281_, _15903_, _15902_);
  or (_15904_, _15893_, _15078_);
  or (_15905_, _15885_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_15906_, _15905_, _15888_);
  and (_15907_, _15906_, _15904_);
  and (_15908_, _15887_, _15084_);
  or (_41282_, _15908_, _15907_);
  or (_15909_, _15893_, _15283_);
  or (_15910_, _15885_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_15911_, _15910_, _15888_);
  and (_15912_, _15911_, _15909_);
  and (_15913_, _15887_, _15289_);
  or (_41283_, _15913_, _15912_);
  or (_15914_, _15893_, _15480_);
  or (_15915_, _15885_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_15916_, _15915_, _15888_);
  and (_15917_, _15916_, _15914_);
  and (_15918_, _15887_, _15487_);
  or (_41284_, _15918_, _15917_);
  or (_15919_, _15893_, _15679_);
  or (_15920_, _15885_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_15921_, _15920_, _15888_);
  and (_15922_, _15921_, _15919_);
  and (_15923_, _15887_, _15686_);
  or (_41285_, _15923_, _15922_);
  or (_15924_, _15893_, _09408_);
  or (_15925_, _15885_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_15926_, _15925_, _15888_);
  and (_15927_, _15926_, _15924_);
  and (_15928_, _15887_, _09446_);
  or (_41287_, _15928_, _15927_);
  and (_15929_, _15838_, _15743_);
  nand (_15930_, _15929_, _15697_);
  or (_15931_, _15929_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_15932_, _15842_, _08588_);
  not (_15933_, _15932_);
  and (_15934_, _15933_, _15931_);
  and (_15935_, _15934_, _15930_);
  and (_15936_, _15932_, _14496_);
  or (_41289_, _15936_, _15935_);
  not (_15937_, _15929_);
  or (_15938_, _15937_, _14691_);
  or (_15939_, _15929_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_15940_, _15939_, _15933_);
  and (_15941_, _15940_, _15938_);
  and (_15942_, _15932_, _14697_);
  or (_41292_, _15942_, _15941_);
  or (_15943_, _15937_, _14887_);
  or (_15944_, _15929_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_15945_, _15944_, _15933_);
  and (_15946_, _15945_, _15943_);
  and (_15947_, _15932_, _14893_);
  or (_41293_, _15947_, _15946_);
  or (_15948_, _15937_, _15078_);
  or (_15949_, _15929_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_15950_, _15949_, _15933_);
  and (_15951_, _15950_, _15948_);
  and (_15952_, _15932_, _15084_);
  or (_41294_, _15952_, _15951_);
  or (_15953_, _15937_, _15283_);
  or (_15954_, _15929_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_15955_, _15954_, _15933_);
  and (_15956_, _15955_, _15953_);
  and (_15957_, _15932_, _15289_);
  or (_41295_, _15957_, _15956_);
  or (_15958_, _15937_, _15480_);
  or (_15959_, _15929_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_15960_, _15959_, _15933_);
  and (_15961_, _15960_, _15958_);
  and (_15962_, _15932_, _15487_);
  or (_41296_, _15962_, _15961_);
  or (_15963_, _15937_, _15679_);
  or (_15964_, _15929_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_15965_, _15964_, _15933_);
  and (_15966_, _15965_, _15963_);
  and (_15967_, _15932_, _15686_);
  or (_41298_, _15967_, _15966_);
  or (_15968_, _15937_, _09408_);
  or (_15969_, _15929_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_15970_, _15969_, _15933_);
  and (_15971_, _15970_, _15968_);
  and (_15972_, _15932_, _09446_);
  or (_41299_, _15972_, _15971_);
  and (_15973_, _15842_, _06234_);
  not (_15974_, _15973_);
  or (_15975_, _15974_, _14496_);
  and (_15976_, _15838_, _15791_);
  nor (_15977_, _15976_, _07287_);
  and (_15978_, _15976_, _15696_);
  or (_15979_, _15978_, _15973_);
  or (_15980_, _15979_, _15977_);
  and (_41302_, _15980_, _15975_);
  not (_15981_, _15976_);
  or (_15982_, _15981_, _14691_);
  or (_15983_, _15976_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_15984_, _15983_, _15974_);
  and (_15985_, _15984_, _15982_);
  and (_15986_, _15973_, _14697_);
  or (_41304_, _15986_, _15985_);
  or (_15987_, _15981_, _14887_);
  or (_15988_, _15976_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_15989_, _15988_, _15974_);
  and (_15990_, _15989_, _15987_);
  and (_15991_, _15973_, _14893_);
  or (_41305_, _15991_, _15990_);
  or (_15992_, _15981_, _15078_);
  or (_15993_, _15976_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_15994_, _15993_, _15974_);
  and (_15995_, _15994_, _15992_);
  and (_15996_, _15973_, _15084_);
  or (_41306_, _15996_, _15995_);
  or (_15997_, _15981_, _15283_);
  or (_15998_, _15976_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_15999_, _15998_, _15974_);
  and (_16000_, _15999_, _15997_);
  and (_16001_, _15973_, _15289_);
  or (_41307_, _16001_, _16000_);
  or (_16002_, _15981_, _15480_);
  or (_16003_, _15976_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_16004_, _16003_, _15974_);
  and (_16005_, _16004_, _16002_);
  and (_16006_, _15973_, _15487_);
  or (_41308_, _16006_, _16005_);
  or (_16007_, _15981_, _15679_);
  or (_16008_, _15976_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_16009_, _16008_, _15974_);
  and (_16010_, _16009_, _16007_);
  and (_16011_, _15973_, _15686_);
  or (_41310_, _16011_, _16010_);
  or (_16012_, _15981_, _09408_);
  or (_16013_, _15976_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_16014_, _16013_, _15974_);
  and (_16015_, _16014_, _16012_);
  and (_16016_, _15973_, _09446_);
  or (_41311_, _16016_, _16015_);
  and (_16017_, _07831_, _07659_);
  and (_16018_, _16017_, _14311_);
  or (_16019_, _16018_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_16020_, _16018_, _15697_);
  and (_16021_, _16020_, _16019_);
  not (_16022_, _07837_);
  and (_16023_, _07845_, _16022_);
  and (_16024_, _16023_, _06236_);
  or (_16025_, _16024_, _16021_);
  not (_16026_, _07845_);
  or (_16027_, _16026_, _07835_);
  or (_16028_, _16027_, _14495_);
  and (_41315_, _16028_, _16025_);
  not (_16029_, _16018_);
  or (_16030_, _16029_, _14691_);
  or (_16031_, _16018_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_16032_, _16031_, _16027_);
  and (_16033_, _16032_, _16030_);
  and (_16034_, _16024_, _14697_);
  or (_41316_, _16034_, _16033_);
  or (_16035_, _16029_, _14887_);
  or (_16036_, _16018_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_16037_, _16036_, _16027_);
  and (_16038_, _16037_, _16035_);
  and (_16039_, _16024_, _14893_);
  or (_41318_, _16039_, _16038_);
  or (_16040_, _16029_, _15078_);
  or (_16041_, _16018_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_16042_, _16041_, _16027_);
  and (_16043_, _16042_, _16040_);
  and (_16044_, _16024_, _15084_);
  or (_41319_, _16044_, _16043_);
  or (_16045_, _16029_, _15283_);
  or (_16046_, _16018_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_16047_, _16046_, _16027_);
  and (_16048_, _16047_, _16045_);
  and (_16049_, _16024_, _15289_);
  or (_41320_, _16049_, _16048_);
  or (_16050_, _16029_, _15480_);
  or (_16051_, _16018_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_16052_, _16051_, _16027_);
  and (_16053_, _16052_, _16050_);
  and (_16054_, _16024_, _15487_);
  or (_41321_, _16054_, _16053_);
  or (_16055_, _16029_, _15679_);
  or (_16056_, _16018_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_16057_, _16056_, _16027_);
  and (_16058_, _16057_, _16055_);
  and (_16059_, _16024_, _15686_);
  or (_41322_, _16059_, _16058_);
  or (_16060_, _16029_, _09408_);
  or (_16061_, _16018_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_16062_, _16061_, _16027_);
  and (_16063_, _16062_, _16060_);
  and (_16064_, _16024_, _09446_);
  or (_41324_, _16064_, _16063_);
  and (_16065_, _16017_, _15693_);
  or (_16066_, _16065_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_16067_, _16065_, _15697_);
  and (_16068_, _16067_, _16066_);
  and (_16069_, _16023_, _07512_);
  or (_16070_, _16069_, _16068_);
  nand (_16071_, _07845_, _07513_);
  or (_16072_, _16071_, _14495_);
  and (_41327_, _16072_, _16070_);
  not (_16073_, _16065_);
  or (_16074_, _16073_, _14691_);
  or (_16075_, _16065_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_16076_, _16075_, _16071_);
  and (_16077_, _16076_, _16074_);
  and (_16078_, _16069_, _14697_);
  or (_41328_, _16078_, _16077_);
  or (_16079_, _16073_, _14887_);
  or (_16080_, _16065_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_16081_, _16080_, _16071_);
  and (_16082_, _16081_, _16079_);
  and (_16083_, _16069_, _14893_);
  or (_41330_, _16083_, _16082_);
  or (_16084_, _16073_, _15078_);
  or (_16085_, _16065_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_16086_, _16085_, _16071_);
  and (_16087_, _16086_, _16084_);
  and (_16088_, _16069_, _15084_);
  or (_41331_, _16088_, _16087_);
  or (_16089_, _16073_, _15283_);
  or (_16090_, _16065_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_16091_, _16090_, _16071_);
  and (_16092_, _16091_, _16089_);
  and (_16093_, _16069_, _15289_);
  or (_41332_, _16093_, _16092_);
  or (_16094_, _16073_, _15480_);
  or (_16095_, _16065_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_16096_, _16095_, _16071_);
  and (_16097_, _16096_, _16094_);
  and (_16098_, _16069_, _15487_);
  or (_41333_, _16098_, _16097_);
  or (_16099_, _16073_, _15679_);
  or (_16100_, _16065_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_16101_, _16100_, _16071_);
  and (_16102_, _16101_, _16099_);
  and (_16103_, _16069_, _15686_);
  or (_41334_, _16103_, _16102_);
  or (_16104_, _16073_, _09408_);
  or (_16105_, _16065_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_16106_, _16105_, _16071_);
  and (_16107_, _16106_, _16104_);
  and (_16108_, _16069_, _09446_);
  or (_41336_, _16108_, _16107_);
  and (_16109_, _16017_, _15743_);
  nor (_16110_, _16109_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_16111_, _16109_, _15697_);
  or (_16112_, _16111_, _16110_);
  and (_16113_, _16023_, _08588_);
  not (_16114_, _16113_);
  nand (_16115_, _16114_, _16112_);
  or (_16116_, _16114_, _14496_);
  and (_41339_, _16116_, _16115_);
  not (_16117_, _16109_);
  or (_16118_, _16117_, _14691_);
  or (_16119_, _16109_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_16120_, _16119_, _16114_);
  and (_16121_, _16120_, _16118_);
  and (_16122_, _16113_, _14697_);
  or (_41341_, _16122_, _16121_);
  or (_16123_, _16117_, _14887_);
  or (_16124_, _16109_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_16125_, _16124_, _16114_);
  and (_16126_, _16125_, _16123_);
  and (_16127_, _16113_, _14893_);
  or (_41342_, _16127_, _16126_);
  or (_16128_, _16117_, _15078_);
  or (_16129_, _16109_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_16130_, _16129_, _16114_);
  and (_16131_, _16130_, _16128_);
  and (_16132_, _16113_, _15084_);
  or (_41343_, _16132_, _16131_);
  or (_16133_, _16117_, _15283_);
  or (_16134_, _16109_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_16135_, _16134_, _16114_);
  and (_16136_, _16135_, _16133_);
  and (_16137_, _16113_, _15289_);
  or (_41344_, _16137_, _16136_);
  or (_16138_, _16117_, _15480_);
  or (_16139_, _16109_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_16140_, _16139_, _16114_);
  and (_16141_, _16140_, _16138_);
  and (_16142_, _16113_, _15487_);
  or (_41345_, _16142_, _16141_);
  or (_16143_, _16117_, _15679_);
  or (_16144_, _16109_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_16145_, _16144_, _16114_);
  and (_16146_, _16145_, _16143_);
  and (_16147_, _16113_, _15686_);
  or (_41347_, _16147_, _16146_);
  or (_16148_, _16117_, _09408_);
  or (_16149_, _16109_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_16150_, _16149_, _16114_);
  and (_16151_, _16150_, _16148_);
  and (_16152_, _16113_, _09446_);
  or (_41348_, _16152_, _16151_);
  and (_16153_, _16017_, _07510_);
  or (_16154_, _16153_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_16155_, _16153_, _15697_);
  and (_16156_, _16155_, _16154_);
  and (_16157_, _16023_, _06234_);
  or (_16158_, _16157_, _16156_);
  not (_16159_, _16157_);
  or (_16160_, _16159_, _14496_);
  and (_41351_, _16160_, _16158_);
  and (_16161_, _16017_, _15791_);
  or (_16162_, _16161_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_16163_, _16162_, _16159_);
  not (_16164_, _16161_);
  or (_16165_, _16164_, _14691_);
  and (_16166_, _16165_, _16163_);
  and (_16167_, _16157_, _14697_);
  or (_41353_, _16167_, _16166_);
  or (_16168_, _16161_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_16169_, _16168_, _16159_);
  or (_16170_, _16164_, _14887_);
  and (_16171_, _16170_, _16169_);
  and (_16172_, _16157_, _14893_);
  or (_41354_, _16172_, _16171_);
  or (_16173_, _16161_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_16174_, _16173_, _16159_);
  or (_16175_, _16164_, _15078_);
  and (_16176_, _16175_, _16174_);
  and (_16177_, _16157_, _15084_);
  or (_41355_, _16177_, _16176_);
  or (_16178_, _16161_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_16179_, _16178_, _16159_);
  or (_16180_, _16164_, _15283_);
  and (_16181_, _16180_, _16179_);
  and (_16182_, _16157_, _15289_);
  or (_41356_, _16182_, _16181_);
  or (_16183_, _16161_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_16184_, _16183_, _16159_);
  or (_16185_, _16164_, _15480_);
  and (_16186_, _16185_, _16184_);
  and (_16187_, _16157_, _15487_);
  or (_41357_, _16187_, _16186_);
  or (_16188_, _16161_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_16189_, _16188_, _16159_);
  or (_16190_, _16164_, _15679_);
  and (_16191_, _16190_, _16189_);
  and (_16192_, _16157_, _15686_);
  or (_41359_, _16192_, _16191_);
  nor (_16193_, _16161_, \oc8051_golden_model_1.IRAM[11] [7]);
  not (_16194_, _16153_);
  nor (_16195_, _16194_, _09408_);
  or (_16196_, _16195_, _16193_);
  nor (_16197_, _16196_, _16157_);
  and (_16198_, _16157_, _09446_);
  or (_41360_, _16198_, _16197_);
  and (_16199_, _14311_, _07832_);
  nand (_16200_, _16199_, _15697_);
  and (_16201_, _07846_, _06236_);
  not (_16202_, _16201_);
  or (_16203_, _16199_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_16204_, _16203_, _16202_);
  and (_16205_, _16204_, _16200_);
  and (_16206_, _16201_, _14496_);
  or (_41364_, _16206_, _16205_);
  not (_16207_, _16199_);
  or (_16208_, _16207_, _14691_);
  or (_16209_, _16199_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_16210_, _16209_, _16202_);
  and (_16211_, _16210_, _16208_);
  and (_16212_, _16201_, _14697_);
  or (_41365_, _16212_, _16211_);
  or (_16213_, _16199_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_16214_, _16213_, _16202_);
  or (_16215_, _16207_, _14887_);
  and (_16216_, _16215_, _16214_);
  and (_16217_, _16201_, _14893_);
  or (_41366_, _16217_, _16216_);
  or (_16218_, _16199_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_16219_, _16218_, _16202_);
  or (_16220_, _16207_, _15078_);
  and (_16221_, _16220_, _16219_);
  and (_16222_, _16201_, _15084_);
  or (_41367_, _16222_, _16221_);
  or (_16223_, _16207_, _15283_);
  or (_16224_, _16199_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_16225_, _16224_, _16202_);
  and (_16226_, _16225_, _16223_);
  and (_16227_, _16201_, _15289_);
  or (_41369_, _16227_, _16226_);
  or (_16228_, _16207_, _15480_);
  or (_16229_, _16199_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_16230_, _16229_, _16202_);
  and (_16231_, _16230_, _16228_);
  and (_16232_, _16201_, _15487_);
  or (_41370_, _16232_, _16231_);
  or (_16233_, _16207_, _15679_);
  or (_16234_, _16199_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_16235_, _16234_, _16202_);
  and (_16236_, _16235_, _16233_);
  and (_16237_, _16201_, _15686_);
  or (_41371_, _16237_, _16236_);
  or (_16238_, _16207_, _09408_);
  or (_16239_, _16199_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_16240_, _16239_, _16202_);
  and (_16241_, _16240_, _16238_);
  and (_16242_, _16201_, _09446_);
  or (_41372_, _16242_, _16241_);
  and (_16243_, _15693_, _07832_);
  nand (_16244_, _16243_, _15697_);
  and (_16245_, _07846_, _07512_);
  not (_16246_, _16245_);
  or (_16247_, _16243_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_16248_, _16247_, _16246_);
  and (_16249_, _16248_, _16244_);
  and (_16250_, _16245_, _14496_);
  or (_41376_, _16250_, _16249_);
  and (_16251_, _16245_, _14697_);
  or (_16252_, _16243_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_16253_, _16252_, _16246_);
  not (_16254_, _16243_);
  or (_16255_, _16254_, _14691_);
  and (_16256_, _16255_, _16253_);
  or (_41377_, _16256_, _16251_);
  and (_16257_, _16245_, _14893_);
  or (_16258_, _16243_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_16259_, _16258_, _16246_);
  or (_16260_, _16254_, _14887_);
  and (_16261_, _16260_, _16259_);
  or (_41378_, _16261_, _16257_);
  and (_16262_, _16245_, _15084_);
  or (_16263_, _16243_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_16264_, _16263_, _16246_);
  or (_16265_, _16254_, _15078_);
  and (_16266_, _16265_, _16264_);
  or (_41379_, _16266_, _16262_);
  or (_16267_, _16243_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_16268_, _16267_, _16246_);
  or (_16269_, _16254_, _15283_);
  and (_16270_, _16269_, _16268_);
  and (_16271_, _16245_, _15289_);
  or (_41381_, _16271_, _16270_);
  and (_16272_, _16245_, _15487_);
  or (_16273_, _16243_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_16274_, _16273_, _16246_);
  or (_16275_, _16254_, _15480_);
  and (_16276_, _16275_, _16274_);
  or (_41382_, _16276_, _16272_);
  or (_16277_, _16243_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_16278_, _16277_, _16246_);
  or (_16279_, _16254_, _15679_);
  and (_16280_, _16279_, _16278_);
  and (_16281_, _16245_, _15686_);
  or (_41383_, _16281_, _16280_);
  or (_16282_, _16243_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_16283_, _16282_, _16246_);
  or (_16284_, _16254_, _09408_);
  and (_16285_, _16284_, _16283_);
  and (_16286_, _16245_, _09446_);
  or (_41384_, _16286_, _16285_);
  and (_16287_, _15743_, _07832_);
  or (_16288_, _16287_, \oc8051_golden_model_1.IRAM[14] [0]);
  nand (_16289_, _16287_, _15697_);
  and (_16290_, _16289_, _16288_);
  and (_16291_, _08588_, _07846_);
  or (_16292_, _16291_, _16290_);
  not (_16293_, _16291_);
  or (_16294_, _16293_, _14496_);
  and (_41388_, _16294_, _16292_);
  or (_16295_, _16287_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_16296_, _16295_, _16293_);
  not (_16297_, _16287_);
  or (_16298_, _16297_, _14691_);
  and (_16299_, _16298_, _16296_);
  and (_16300_, _16291_, _14697_);
  or (_41389_, _16300_, _16299_);
  or (_16301_, _16287_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_16302_, _16301_, _16293_);
  or (_16303_, _16297_, _14887_);
  and (_16304_, _16303_, _16302_);
  and (_16305_, _16291_, _14893_);
  or (_41390_, _16305_, _16304_);
  or (_16306_, _16287_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_16307_, _16306_, _16293_);
  or (_16308_, _16297_, _15078_);
  and (_16309_, _16308_, _16307_);
  and (_16310_, _16291_, _15084_);
  or (_41391_, _16310_, _16309_);
  or (_16311_, _16287_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_16312_, _16311_, _16293_);
  or (_16313_, _16297_, _15283_);
  and (_16314_, _16313_, _16312_);
  and (_16315_, _16291_, _15289_);
  or (_41392_, _16315_, _16314_);
  or (_16316_, _16287_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_16317_, _16316_, _16293_);
  or (_16318_, _16297_, _15480_);
  and (_16319_, _16318_, _16317_);
  and (_16320_, _16291_, _15487_);
  or (_41393_, _16320_, _16319_);
  or (_16321_, _16287_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_16322_, _16321_, _16293_);
  or (_16323_, _16297_, _15679_);
  and (_16324_, _16323_, _16322_);
  and (_16325_, _16291_, _15686_);
  or (_41394_, _16325_, _16324_);
  or (_16326_, _16287_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_16327_, _16326_, _16293_);
  or (_16328_, _16297_, _09408_);
  and (_16329_, _16328_, _16327_);
  and (_16330_, _16291_, _09446_);
  or (_41395_, _16330_, _16329_);
  or (_16331_, _07833_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_16332_, _15697_, _07833_);
  and (_16333_, _16332_, _16331_);
  or (_16334_, _16333_, _07847_);
  or (_16335_, _14496_, _07848_);
  and (_41399_, _16335_, _16334_);
  or (_16336_, _07833_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_16337_, _16336_, _07848_);
  or (_16338_, _14691_, _07850_);
  and (_16339_, _16338_, _16337_);
  and (_16340_, _14697_, _07847_);
  or (_41400_, _16340_, _16339_);
  or (_16341_, _07833_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_16342_, _16341_, _07848_);
  or (_16343_, _14887_, _07850_);
  and (_16344_, _16343_, _16342_);
  and (_16345_, _14893_, _07847_);
  or (_41401_, _16345_, _16344_);
  or (_16346_, _07833_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_16347_, _16346_, _07848_);
  or (_16348_, _15078_, _07850_);
  and (_16349_, _16348_, _16347_);
  and (_16350_, _15084_, _07847_);
  or (_41403_, _16350_, _16349_);
  or (_16351_, _07833_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_16352_, _16351_, _07848_);
  or (_16353_, _15283_, _07850_);
  and (_16354_, _16353_, _16352_);
  and (_16355_, _15289_, _07847_);
  or (_41404_, _16355_, _16354_);
  or (_16356_, _07833_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_16357_, _16356_, _07848_);
  or (_16358_, _15480_, _07850_);
  and (_16359_, _16358_, _16357_);
  and (_16360_, _15487_, _07847_);
  or (_41405_, _16360_, _16359_);
  or (_16361_, _07833_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_16362_, _16361_, _07848_);
  or (_16363_, _15679_, _07850_);
  and (_16364_, _16363_, _16362_);
  and (_16365_, _15686_, _07847_);
  or (_41406_, _16365_, _16364_);
  nor (_16366_, _01452_, _10058_);
  nand (_16367_, _11218_, _07911_);
  nor (_16368_, _07911_, _10058_);
  nor (_16369_, _16368_, _07210_);
  nand (_16370_, _16369_, _16367_);
  and (_16371_, _07911_, _08908_);
  or (_16372_, _16371_, _16368_);
  or (_16373_, _16372_, _07198_);
  and (_16374_, _07911_, _07325_);
  or (_16375_, _16374_, _16368_);
  or (_16376_, _16375_, _07188_);
  nor (_16377_, _08351_, _09454_);
  or (_16378_, _16377_, _16368_);
  and (_16379_, _16378_, _06251_);
  nor (_16380_, _07123_, _10058_);
  and (_16381_, _07911_, \oc8051_golden_model_1.ACC [0]);
  or (_16382_, _16381_, _16368_);
  and (_16383_, _16382_, _07123_);
  or (_16384_, _16383_, _16380_);
  and (_16385_, _16384_, _06252_);
  or (_16386_, _16385_, _06475_);
  or (_16387_, _16386_, _16379_);
  and (_16388_, _14341_, _08547_);
  nor (_16389_, _08547_, _10058_);
  or (_16390_, _16389_, _06476_);
  or (_16391_, _16390_, _16388_);
  and (_16392_, _16391_, _16387_);
  or (_16393_, _16392_, _06468_);
  or (_16394_, _16375_, _07142_);
  and (_16395_, _16394_, _16393_);
  or (_16396_, _16395_, _06466_);
  or (_16397_, _16382_, _06801_);
  and (_16398_, _16397_, _06484_);
  and (_16399_, _16398_, _16396_);
  and (_16400_, _16368_, _06483_);
  or (_16401_, _16400_, _06461_);
  or (_16402_, _16401_, _16399_);
  or (_16403_, _16378_, _07164_);
  and (_16404_, _16403_, _16402_);
  or (_16405_, _16404_, _09487_);
  nor (_16406_, _09997_, _09995_);
  nor (_16407_, _16406_, _09998_);
  or (_16408_, _16407_, _09494_);
  and (_16409_, _16408_, _06242_);
  and (_16410_, _16409_, _16405_);
  and (_16411_, _14372_, _08547_);
  or (_16412_, _16411_, _16389_);
  and (_16413_, _16412_, _06241_);
  or (_16414_, _16413_, _07187_);
  or (_16415_, _16414_, _16410_);
  and (_16416_, _16415_, _16376_);
  or (_16417_, _16416_, _07182_);
  and (_16418_, _09342_, _07911_);
  or (_16419_, _16368_, _07183_);
  or (_16420_, _16419_, _16418_);
  and (_16421_, _16420_, _16417_);
  or (_16422_, _16421_, _05968_);
  and (_16423_, _14427_, _07911_);
  or (_16424_, _16368_, _06336_);
  or (_16425_, _16424_, _16423_);
  and (_16426_, _16425_, _10052_);
  and (_16427_, _16426_, _16422_);
  or (_16428_, _10392_, _10347_);
  or (_16429_, _10398_, _16428_);
  nand (_16430_, _10398_, _05997_);
  and (_16431_, _16430_, _10046_);
  and (_16432_, _16431_, _16429_);
  or (_16433_, _16432_, _06371_);
  or (_16434_, _16433_, _16427_);
  and (_16435_, _16434_, _16373_);
  or (_16436_, _16435_, _06367_);
  and (_16437_, _14442_, _07911_);
  or (_16438_, _16437_, _16368_);
  or (_16439_, _16438_, _07218_);
  and (_16440_, _16439_, _07216_);
  and (_16441_, _16440_, _16436_);
  nor (_16442_, _12526_, _09454_);
  or (_16443_, _16442_, _16368_);
  and (_16444_, _16367_, _06533_);
  and (_16445_, _16444_, _16443_);
  or (_16446_, _16445_, _16441_);
  and (_16447_, _16446_, _07213_);
  nand (_16448_, _16372_, _06366_);
  nor (_16449_, _16448_, _16377_);
  or (_16450_, _16449_, _06541_);
  or (_16451_, _16450_, _16447_);
  and (_16452_, _16451_, _16370_);
  or (_16453_, _16452_, _06383_);
  and (_16454_, _14325_, _07911_);
  or (_16455_, _16368_, _07231_);
  or (_16456_, _16455_, _16454_);
  and (_16457_, _16456_, _07229_);
  and (_16458_, _16457_, _16453_);
  and (_16459_, _16443_, _06528_);
  or (_16460_, _16459_, _06563_);
  or (_16461_, _16460_, _16458_);
  or (_16462_, _16378_, _07241_);
  and (_16463_, _16462_, _16461_);
  or (_16464_, _16463_, _06199_);
  or (_16465_, _16368_, _06571_);
  and (_16466_, _16465_, _16464_);
  or (_16467_, _16466_, _06188_);
  or (_16468_, _16378_, _06189_);
  and (_16469_, _16468_, _01452_);
  and (_16470_, _16469_, _16467_);
  or (_16471_, _16470_, _16366_);
  and (_43761_, _16471_, _43223_);
  nor (_16472_, _01452_, _10053_);
  nor (_16473_, _07911_, _10053_);
  nor (_16474_, _11216_, _09454_);
  or (_16475_, _16474_, _16473_);
  or (_16476_, _16475_, _07229_);
  or (_16477_, _07911_, \oc8051_golden_model_1.B [1]);
  nand (_16478_, _07911_, _07018_);
  and (_16479_, _16478_, _06371_);
  and (_16480_, _16479_, _16477_);
  nor (_16481_, _09454_, _07120_);
  or (_16482_, _16481_, _16473_);
  or (_16483_, _16482_, _07142_);
  and (_16484_, _14503_, _07911_);
  not (_16485_, _16484_);
  and (_16486_, _16485_, _16477_);
  or (_16487_, _16486_, _06252_);
  and (_16488_, _07911_, \oc8051_golden_model_1.ACC [1]);
  or (_16489_, _16488_, _16473_);
  and (_16490_, _16489_, _07123_);
  nor (_16491_, _07123_, _10053_);
  or (_16492_, _16491_, _06251_);
  or (_16493_, _16492_, _16490_);
  and (_16494_, _16493_, _06476_);
  and (_16495_, _16494_, _16487_);
  nor (_16496_, _08547_, _10053_);
  and (_16497_, _14510_, _08547_);
  or (_16498_, _16497_, _16496_);
  and (_16499_, _16498_, _06475_);
  or (_16500_, _16499_, _06468_);
  or (_16501_, _16500_, _16495_);
  and (_16502_, _16501_, _16483_);
  or (_16503_, _16502_, _06466_);
  or (_16504_, _16489_, _06801_);
  and (_16505_, _16504_, _16503_);
  or (_16506_, _16505_, _06483_);
  and (_16507_, _14513_, _08547_);
  or (_16508_, _16507_, _16496_);
  or (_16509_, _16508_, _06484_);
  and (_16510_, _16509_, _07164_);
  and (_16511_, _16510_, _16506_);
  or (_16512_, _16496_, _14509_);
  and (_16513_, _16512_, _06461_);
  and (_16514_, _16513_, _16498_);
  or (_16515_, _16514_, _09487_);
  or (_16516_, _16515_, _16511_);
  or (_16517_, _09941_, _09940_);
  nand (_16518_, _16517_, _09999_);
  or (_16519_, _16517_, _09999_);
  and (_16520_, _16519_, _16518_);
  or (_16521_, _16520_, _09494_);
  and (_16522_, _16521_, _06242_);
  and (_16523_, _16522_, _16516_);
  or (_16524_, _16496_, _14553_);
  and (_16525_, _16524_, _06241_);
  and (_16526_, _16525_, _16498_);
  or (_16527_, _16526_, _07187_);
  or (_16528_, _16527_, _16523_);
  or (_16529_, _16482_, _07188_);
  and (_16530_, _16529_, _16528_);
  or (_16531_, _16530_, _07182_);
  and (_16532_, _09297_, _07911_);
  or (_16533_, _16473_, _07183_);
  or (_16534_, _16533_, _16532_);
  and (_16535_, _16534_, _06336_);
  and (_16536_, _16535_, _16531_);
  or (_16537_, _14609_, _09454_);
  and (_16538_, _16477_, _05968_);
  and (_16539_, _16538_, _16537_);
  or (_16540_, _16539_, _10046_);
  or (_16541_, _16540_, _16536_);
  nor (_16542_, _10393_, _10391_);
  or (_16543_, _16542_, _10394_);
  nor (_16544_, _16543_, _10398_);
  and (_16545_, _10398_, _10344_);
  or (_16546_, _16545_, _16544_);
  or (_16547_, _16546_, _10052_);
  and (_16548_, _16547_, _07198_);
  and (_16549_, _16548_, _16541_);
  or (_16550_, _16549_, _16480_);
  and (_16551_, _16550_, _07218_);
  or (_16552_, _14625_, _09454_);
  and (_16553_, _16477_, _06367_);
  and (_16554_, _16553_, _16552_);
  or (_16555_, _16554_, _06533_);
  or (_16556_, _16555_, _16551_);
  and (_16557_, _11217_, _07911_);
  or (_16558_, _16557_, _16473_);
  or (_16559_, _16558_, _07216_);
  and (_16560_, _16559_, _07213_);
  and (_16561_, _16560_, _16556_);
  or (_16562_, _14623_, _09454_);
  and (_16563_, _16477_, _06366_);
  and (_16564_, _16563_, _16562_);
  or (_16565_, _16564_, _06541_);
  or (_16566_, _16565_, _16561_);
  and (_16567_, _16488_, _08302_);
  or (_16568_, _16473_, _07210_);
  or (_16569_, _16568_, _16567_);
  and (_16570_, _16569_, _07231_);
  and (_16571_, _16570_, _16566_);
  or (_16572_, _16478_, _08302_);
  and (_16573_, _16477_, _06383_);
  and (_16574_, _16573_, _16572_);
  or (_16575_, _16574_, _06528_);
  or (_16576_, _16575_, _16571_);
  and (_16577_, _16576_, _16476_);
  or (_16578_, _16577_, _06563_);
  or (_16579_, _16486_, _07241_);
  and (_16580_, _16579_, _06571_);
  and (_16581_, _16580_, _16578_);
  and (_16582_, _16508_, _06199_);
  or (_16583_, _16582_, _06188_);
  or (_16584_, _16583_, _16581_);
  or (_16585_, _16473_, _06189_);
  or (_16586_, _16585_, _16484_);
  and (_16587_, _16586_, _01452_);
  and (_16588_, _16587_, _16584_);
  or (_16589_, _16588_, _16472_);
  and (_43762_, _16589_, _43223_);
  nor (_16590_, _01452_, _10111_);
  nor (_16591_, _07911_, _10111_);
  and (_16592_, _07911_, _08945_);
  or (_16593_, _16592_, _16591_);
  or (_16594_, _16593_, _07198_);
  nor (_16595_, _09454_, _07578_);
  or (_16596_, _16595_, _16591_);
  or (_16597_, _16596_, _07188_);
  and (_16598_, _07911_, \oc8051_golden_model_1.ACC [2]);
  or (_16599_, _16598_, _16591_);
  or (_16600_, _16599_, _06801_);
  and (_16601_, _14712_, _07911_);
  or (_16602_, _16601_, _16591_);
  or (_16603_, _16602_, _06252_);
  and (_16604_, _16599_, _07123_);
  nor (_16605_, _07123_, _10111_);
  or (_16606_, _16605_, _06251_);
  or (_16607_, _16606_, _16604_);
  and (_16608_, _16607_, _06476_);
  and (_16609_, _16608_, _16603_);
  nor (_16610_, _08547_, _10111_);
  and (_16611_, _14702_, _08547_);
  or (_16612_, _16611_, _16610_);
  and (_16613_, _16612_, _06475_);
  or (_16614_, _16613_, _06468_);
  or (_16615_, _16614_, _16609_);
  or (_16616_, _16596_, _07142_);
  and (_16617_, _16616_, _16615_);
  or (_16618_, _16617_, _06466_);
  and (_16619_, _16618_, _16600_);
  or (_16620_, _16619_, _06483_);
  and (_16621_, _14706_, _08547_);
  or (_16622_, _16621_, _16610_);
  or (_16623_, _16622_, _06484_);
  and (_16624_, _16623_, _07164_);
  and (_16625_, _16624_, _16620_);
  or (_16626_, _16610_, _14739_);
  and (_16627_, _16626_, _06461_);
  and (_16628_, _16627_, _16612_);
  or (_16629_, _16628_, _09487_);
  or (_16630_, _16629_, _16625_);
  or (_16631_, _10001_, _09897_);
  and (_16632_, _16631_, _10002_);
  or (_16633_, _16632_, _09494_);
  and (_16634_, _16633_, _06242_);
  and (_16635_, _16634_, _16630_);
  or (_16636_, _16610_, _14703_);
  and (_16637_, _16636_, _06241_);
  and (_16638_, _16637_, _16612_);
  or (_16639_, _16638_, _07187_);
  or (_16640_, _16639_, _16635_);
  and (_16641_, _16640_, _16597_);
  or (_16642_, _16641_, _07182_);
  and (_16643_, _09251_, _07911_);
  or (_16644_, _16591_, _07183_);
  or (_16645_, _16644_, _16643_);
  and (_16646_, _16645_, _16642_);
  or (_16647_, _16646_, _05968_);
  and (_16648_, _14808_, _07911_);
  or (_16649_, _16591_, _06336_);
  or (_16650_, _16649_, _16648_);
  and (_16651_, _16650_, _10052_);
  and (_16652_, _16651_, _16647_);
  nand (_16653_, _10398_, _10335_);
  nor (_16654_, _10394_, _10345_);
  not (_16655_, _16654_);
  and (_16656_, _16655_, _10338_);
  nor (_16657_, _16655_, _10338_);
  nor (_16658_, _16657_, _16656_);
  or (_16659_, _16658_, _10398_);
  and (_16660_, _16659_, _10046_);
  and (_16661_, _16660_, _16653_);
  or (_16662_, _16661_, _06371_);
  or (_16663_, _16662_, _16652_);
  and (_16664_, _16663_, _16594_);
  or (_16665_, _16664_, _06367_);
  and (_16666_, _14824_, _07911_);
  or (_16667_, _16666_, _16591_);
  or (_16668_, _16667_, _07218_);
  and (_16669_, _16668_, _07216_);
  and (_16670_, _16669_, _16665_);
  and (_16671_, _11214_, _07911_);
  or (_16672_, _16671_, _16591_);
  and (_16673_, _16672_, _06533_);
  or (_16674_, _16673_, _16670_);
  and (_16675_, _16674_, _07213_);
  or (_16676_, _16591_, _08397_);
  and (_16677_, _16593_, _06366_);
  and (_16678_, _16677_, _16676_);
  or (_16679_, _16678_, _16675_);
  and (_16680_, _16679_, _07210_);
  and (_16681_, _16599_, _06541_);
  and (_16682_, _16681_, _16676_);
  or (_16683_, _16682_, _06383_);
  or (_16684_, _16683_, _16680_);
  and (_16685_, _14821_, _07911_);
  or (_16686_, _16591_, _07231_);
  or (_16687_, _16686_, _16685_);
  and (_16688_, _16687_, _07229_);
  and (_16689_, _16688_, _16684_);
  nor (_16690_, _11213_, _09454_);
  or (_16691_, _16690_, _16591_);
  and (_16692_, _16691_, _06528_);
  or (_16693_, _16692_, _06563_);
  or (_16694_, _16693_, _16689_);
  or (_16695_, _16602_, _07241_);
  and (_16696_, _16695_, _06571_);
  and (_16697_, _16696_, _16694_);
  and (_16698_, _16622_, _06199_);
  or (_16699_, _16698_, _06188_);
  or (_16700_, _16699_, _16697_);
  and (_16701_, _14884_, _07911_);
  or (_16702_, _16591_, _06189_);
  or (_16703_, _16702_, _16701_);
  and (_16704_, _16703_, _01452_);
  and (_16705_, _16704_, _16700_);
  or (_16706_, _16705_, _16590_);
  and (_43763_, _16706_, _43223_);
  nor (_16707_, _01452_, _10097_);
  nor (_16708_, _07911_, _10097_);
  and (_16709_, _07911_, _08872_);
  or (_16710_, _16709_, _16708_);
  or (_16711_, _16710_, _07198_);
  and (_16712_, _15003_, _07911_);
  or (_16713_, _16712_, _16708_);
  and (_16714_, _16713_, _05968_);
  nor (_16715_, _08547_, _10097_);
  and (_16716_, _14906_, _08547_);
  or (_16717_, _16716_, _16715_);
  or (_16718_, _16715_, _14931_);
  and (_16719_, _16718_, _16717_);
  or (_16720_, _16719_, _07164_);
  and (_16721_, _14898_, _07911_);
  or (_16722_, _16721_, _16708_);
  or (_16723_, _16722_, _06252_);
  and (_16724_, _07911_, \oc8051_golden_model_1.ACC [3]);
  or (_16725_, _16724_, _16708_);
  and (_16726_, _16725_, _07123_);
  nor (_16727_, _07123_, _10097_);
  or (_16728_, _16727_, _06251_);
  or (_16729_, _16728_, _16726_);
  and (_16730_, _16729_, _06476_);
  and (_16731_, _16730_, _16723_);
  and (_16732_, _16717_, _06475_);
  or (_16733_, _16732_, _06468_);
  or (_16734_, _16733_, _16731_);
  nor (_16735_, _09454_, _07713_);
  or (_16736_, _16735_, _16708_);
  or (_16737_, _16736_, _07142_);
  and (_16738_, _16737_, _16734_);
  or (_16739_, _16738_, _06466_);
  or (_16740_, _16725_, _06801_);
  and (_16741_, _16740_, _06484_);
  and (_16742_, _16741_, _16739_);
  and (_16743_, _14904_, _08547_);
  or (_16744_, _16743_, _16715_);
  and (_16745_, _16744_, _06483_);
  or (_16746_, _16745_, _06461_);
  or (_16747_, _16746_, _16742_);
  and (_16748_, _16747_, _16720_);
  or (_16749_, _16748_, _09487_);
  nor (_16750_, _10004_, _09839_);
  nor (_16751_, _16750_, _10005_);
  or (_16752_, _16751_, _09494_);
  and (_16753_, _16752_, _06242_);
  and (_16754_, _16753_, _16749_);
  or (_16755_, _16715_, _14947_);
  and (_16756_, _16755_, _06241_);
  and (_16757_, _16756_, _16717_);
  or (_16758_, _16757_, _07187_);
  or (_16759_, _16758_, _16754_);
  or (_16760_, _16736_, _07188_);
  and (_16761_, _16760_, _16759_);
  or (_16762_, _16761_, _07182_);
  and (_16763_, _09205_, _07911_);
  or (_16764_, _16708_, _07183_);
  or (_16765_, _16764_, _16763_);
  and (_16766_, _16765_, _06336_);
  and (_16767_, _16766_, _16762_);
  or (_16768_, _16767_, _16714_);
  and (_16769_, _16768_, _10052_);
  nor (_16770_, _16656_, _10337_);
  nor (_16771_, _16770_, _10329_);
  and (_16772_, _16770_, _10329_);
  or (_16773_, _16772_, _16771_);
  or (_16774_, _16773_, _10398_);
  not (_16775_, _10398_);
  or (_16776_, _16775_, _10326_);
  and (_16777_, _16776_, _10046_);
  and (_16778_, _16777_, _16774_);
  or (_16779_, _16778_, _06371_);
  or (_16780_, _16779_, _16769_);
  and (_16781_, _16780_, _16711_);
  or (_16782_, _16781_, _06367_);
  and (_16783_, _15018_, _07911_);
  or (_16784_, _16783_, _16708_);
  or (_16785_, _16784_, _07218_);
  and (_16786_, _16785_, _07216_);
  and (_16787_, _16786_, _16782_);
  and (_16788_, _12523_, _07911_);
  or (_16789_, _16788_, _16708_);
  and (_16790_, _16789_, _06533_);
  or (_16791_, _16790_, _16787_);
  and (_16792_, _16791_, _07213_);
  or (_16793_, _16708_, _08257_);
  and (_16794_, _16710_, _06366_);
  and (_16795_, _16794_, _16793_);
  or (_16796_, _16795_, _16792_);
  and (_16797_, _16796_, _07210_);
  and (_16798_, _16725_, _06541_);
  and (_16799_, _16798_, _16793_);
  or (_16800_, _16799_, _06383_);
  or (_16801_, _16800_, _16797_);
  and (_16802_, _15015_, _07911_);
  or (_16803_, _16708_, _07231_);
  or (_16804_, _16803_, _16802_);
  and (_16805_, _16804_, _07229_);
  and (_16806_, _16805_, _16801_);
  nor (_16807_, _11211_, _09454_);
  or (_16808_, _16807_, _16708_);
  and (_16809_, _16808_, _06528_);
  or (_16810_, _16809_, _06563_);
  or (_16811_, _16810_, _16806_);
  or (_16812_, _16722_, _07241_);
  and (_16813_, _16812_, _06571_);
  and (_16814_, _16813_, _16811_);
  and (_16815_, _16744_, _06199_);
  or (_16816_, _16815_, _06188_);
  or (_16817_, _16816_, _16814_);
  and (_16818_, _15075_, _07911_);
  or (_16819_, _16708_, _06189_);
  or (_16820_, _16819_, _16818_);
  and (_16821_, _16820_, _01452_);
  and (_16822_, _16821_, _16817_);
  or (_16823_, _16822_, _16707_);
  and (_43764_, _16823_, _43223_);
  nor (_16824_, _01452_, _10190_);
  nor (_16825_, _07911_, _10190_);
  and (_16826_, _08892_, _07911_);
  or (_16827_, _16826_, _16825_);
  or (_16828_, _16827_, _07198_);
  and (_16829_, _15198_, _07911_);
  or (_16830_, _16829_, _16825_);
  and (_16831_, _16830_, _05968_);
  nor (_16832_, _08494_, _09454_);
  or (_16833_, _16832_, _16825_);
  or (_16834_, _16833_, _07188_);
  nor (_16835_, _08547_, _10190_);
  and (_16836_, _15089_, _08547_);
  or (_16837_, _16836_, _16835_);
  and (_16838_, _16837_, _06483_);
  or (_16839_, _16833_, _07142_);
  and (_16840_, _15108_, _07911_);
  or (_16841_, _16840_, _16825_);
  or (_16842_, _16841_, _06252_);
  and (_16843_, _07911_, \oc8051_golden_model_1.ACC [4]);
  or (_16844_, _16843_, _16825_);
  and (_16845_, _16844_, _07123_);
  nor (_16846_, _07123_, _10190_);
  or (_16847_, _16846_, _06251_);
  or (_16848_, _16847_, _16845_);
  and (_16849_, _16848_, _06476_);
  and (_16850_, _16849_, _16842_);
  and (_16851_, _15091_, _08547_);
  or (_16852_, _16851_, _16835_);
  and (_16853_, _16852_, _06475_);
  or (_16854_, _16853_, _06468_);
  or (_16855_, _16854_, _16850_);
  and (_16856_, _16855_, _16839_);
  or (_16857_, _16856_, _06466_);
  or (_16858_, _16844_, _06801_);
  and (_16859_, _16858_, _06484_);
  and (_16860_, _16859_, _16857_);
  or (_16861_, _16860_, _16838_);
  and (_16862_, _16861_, _07164_);
  or (_16863_, _16835_, _15125_);
  and (_16864_, _16863_, _06461_);
  and (_16865_, _16864_, _16852_);
  or (_16866_, _16865_, _09487_);
  or (_16867_, _16866_, _16862_);
  or (_16868_, _10008_, _10006_);
  and (_16869_, _16868_, _10009_);
  or (_16870_, _16869_, _09494_);
  and (_16871_, _16870_, _06242_);
  and (_16872_, _16871_, _16867_);
  or (_16873_, _16835_, _15141_);
  and (_16874_, _16873_, _06241_);
  and (_16875_, _16874_, _16852_);
  or (_16876_, _16875_, _07187_);
  or (_16877_, _16876_, _16872_);
  and (_16878_, _16877_, _16834_);
  or (_16879_, _16878_, _07182_);
  and (_16880_, _09159_, _07911_);
  or (_16881_, _16825_, _07183_);
  or (_16882_, _16881_, _16880_);
  and (_16883_, _16882_, _06336_);
  and (_16884_, _16883_, _16879_);
  or (_16885_, _16884_, _16831_);
  and (_16886_, _16885_, _10052_);
  nor (_16887_, _16770_, _10328_);
  or (_16888_, _16887_, _10327_);
  nand (_16889_, _16888_, _10364_);
  or (_16890_, _16888_, _10364_);
  and (_16891_, _16890_, _16889_);
  or (_16892_, _16891_, _10398_);
  nand (_16893_, _10398_, _10361_);
  and (_16894_, _16893_, _10046_);
  and (_16895_, _16894_, _16892_);
  or (_16896_, _16895_, _06371_);
  or (_16897_, _16896_, _16886_);
  and (_16898_, _16897_, _16828_);
  or (_16899_, _16898_, _06367_);
  and (_16900_, _15214_, _07911_);
  or (_16901_, _16900_, _16825_);
  or (_16902_, _16901_, _07218_);
  and (_16903_, _16902_, _07216_);
  and (_16904_, _16903_, _16899_);
  and (_16905_, _11209_, _07911_);
  or (_16906_, _16905_, _16825_);
  and (_16907_, _16906_, _06533_);
  or (_16908_, _16907_, _16904_);
  and (_16909_, _16908_, _07213_);
  or (_16910_, _16825_, _08497_);
  and (_16911_, _16827_, _06366_);
  and (_16912_, _16911_, _16910_);
  or (_16913_, _16912_, _16909_);
  and (_16914_, _16913_, _07210_);
  and (_16915_, _16844_, _06541_);
  and (_16916_, _16915_, _16910_);
  or (_16917_, _16916_, _06383_);
  or (_16918_, _16917_, _16914_);
  and (_16919_, _15211_, _07911_);
  or (_16920_, _16825_, _07231_);
  or (_16921_, _16920_, _16919_);
  and (_16922_, _16921_, _07229_);
  and (_16923_, _16922_, _16918_);
  nor (_16924_, _11208_, _09454_);
  or (_16925_, _16924_, _16825_);
  and (_16926_, _16925_, _06528_);
  or (_16927_, _16926_, _06563_);
  or (_16928_, _16927_, _16923_);
  or (_16929_, _16841_, _07241_);
  and (_16930_, _16929_, _06571_);
  and (_16931_, _16930_, _16928_);
  and (_16932_, _16837_, _06199_);
  or (_16933_, _16932_, _06188_);
  or (_16934_, _16933_, _16931_);
  and (_16935_, _15280_, _07911_);
  or (_16936_, _16825_, _06189_);
  or (_16937_, _16936_, _16935_);
  and (_16938_, _16937_, _01452_);
  and (_16939_, _16938_, _16934_);
  or (_16940_, _16939_, _16824_);
  and (_43765_, _16940_, _43223_);
  nor (_16941_, _01452_, _10181_);
  nor (_16942_, _07911_, _10181_);
  and (_16943_, _08888_, _07911_);
  or (_16944_, _16943_, _16942_);
  or (_16945_, _16944_, _07198_);
  and (_16946_, _15400_, _07911_);
  or (_16947_, _16946_, _16942_);
  and (_16948_, _16947_, _05968_);
  nor (_16949_, _08209_, _09454_);
  or (_16950_, _16949_, _16942_);
  or (_16951_, _16950_, _07188_);
  or (_16952_, _16950_, _07142_);
  and (_16953_, _15311_, _07911_);
  or (_16954_, _16953_, _16942_);
  or (_16955_, _16954_, _06252_);
  and (_16956_, _07911_, \oc8051_golden_model_1.ACC [5]);
  or (_16957_, _16956_, _16942_);
  and (_16958_, _16957_, _07123_);
  nor (_16959_, _07123_, _10181_);
  or (_16960_, _16959_, _06251_);
  or (_16961_, _16960_, _16958_);
  and (_16962_, _16961_, _06476_);
  and (_16963_, _16962_, _16955_);
  nor (_16964_, _08547_, _10181_);
  and (_16965_, _15296_, _08547_);
  or (_16966_, _16965_, _16964_);
  and (_16967_, _16966_, _06475_);
  or (_16968_, _16967_, _06468_);
  or (_16969_, _16968_, _16963_);
  and (_16970_, _16969_, _16952_);
  or (_16971_, _16970_, _06466_);
  or (_16972_, _16957_, _06801_);
  and (_16973_, _16972_, _06484_);
  and (_16974_, _16973_, _16971_);
  and (_16975_, _15294_, _08547_);
  or (_16976_, _16975_, _16964_);
  and (_16977_, _16976_, _06483_);
  or (_16978_, _16977_, _16974_);
  and (_16979_, _16978_, _07164_);
  or (_16980_, _16964_, _15328_);
  and (_16981_, _16980_, _06461_);
  and (_16982_, _16981_, _16966_);
  or (_16983_, _16982_, _09487_);
  or (_16984_, _16983_, _16979_);
  nor (_16985_, _10011_, _09700_);
  nor (_16986_, _16985_, _10012_);
  or (_16987_, _16986_, _09494_);
  and (_16988_, _16987_, _06242_);
  and (_16989_, _16988_, _16984_);
  or (_16990_, _16964_, _15344_);
  and (_16991_, _16990_, _06241_);
  and (_16992_, _16991_, _16966_);
  or (_16993_, _16992_, _07187_);
  or (_16994_, _16993_, _16989_);
  and (_16995_, _16994_, _16951_);
  or (_16996_, _16995_, _07182_);
  and (_16997_, _09113_, _07911_);
  or (_16998_, _16942_, _07183_);
  or (_16999_, _16998_, _16997_);
  and (_17000_, _16999_, _06336_);
  and (_17001_, _17000_, _16996_);
  or (_17002_, _17001_, _16948_);
  and (_17003_, _17002_, _10052_);
  nand (_17004_, _10398_, _10371_);
  not (_17005_, _10363_);
  and (_17006_, _16889_, _17005_);
  nor (_17007_, _17006_, _10374_);
  and (_17008_, _17006_, _10374_);
  or (_17009_, _17008_, _17007_);
  or (_17010_, _17009_, _10398_);
  and (_17011_, _17010_, _10046_);
  and (_17012_, _17011_, _17004_);
  or (_17013_, _17012_, _06371_);
  or (_17014_, _17013_, _17003_);
  and (_17015_, _17014_, _16945_);
  or (_17016_, _17015_, _06367_);
  and (_17017_, _15416_, _07911_);
  or (_17018_, _17017_, _16942_);
  or (_17019_, _17018_, _07218_);
  and (_17020_, _17019_, _07216_);
  and (_17021_, _17020_, _17016_);
  and (_17022_, _11205_, _07911_);
  or (_17023_, _17022_, _16942_);
  and (_17024_, _17023_, _06533_);
  or (_17025_, _17024_, _17021_);
  and (_17026_, _17025_, _07213_);
  or (_17027_, _16942_, _08212_);
  and (_17028_, _16944_, _06366_);
  and (_17029_, _17028_, _17027_);
  or (_17030_, _17029_, _17026_);
  and (_17031_, _17030_, _07210_);
  and (_17032_, _16957_, _06541_);
  and (_17033_, _17032_, _17027_);
  or (_17034_, _17033_, _06383_);
  or (_17035_, _17034_, _17031_);
  and (_17036_, _15413_, _07911_);
  or (_17037_, _16942_, _07231_);
  or (_17038_, _17037_, _17036_);
  and (_17039_, _17038_, _07229_);
  and (_17040_, _17039_, _17035_);
  nor (_17041_, _11204_, _09454_);
  or (_17042_, _17041_, _16942_);
  and (_17043_, _17042_, _06528_);
  or (_17044_, _17043_, _06563_);
  or (_17045_, _17044_, _17040_);
  or (_17046_, _16954_, _07241_);
  and (_17047_, _17046_, _06571_);
  and (_17048_, _17047_, _17045_);
  and (_17049_, _16976_, _06199_);
  or (_17050_, _17049_, _06188_);
  or (_17051_, _17050_, _17048_);
  and (_17052_, _15477_, _07911_);
  or (_17053_, _16942_, _06189_);
  or (_17054_, _17053_, _17052_);
  and (_17055_, _17054_, _01452_);
  and (_17056_, _17055_, _17051_);
  or (_17057_, _17056_, _16941_);
  and (_43767_, _17057_, _43223_);
  nor (_17058_, _01452_, _10310_);
  nor (_17059_, _07911_, _10310_);
  and (_17060_, _15608_, _07911_);
  or (_17061_, _17060_, _17059_);
  or (_17062_, _17061_, _07198_);
  and (_17063_, _15601_, _07911_);
  or (_17064_, _17063_, _17059_);
  and (_17065_, _17064_, _05968_);
  nor (_17066_, _08106_, _09454_);
  or (_17067_, _17066_, _17059_);
  or (_17068_, _17067_, _07188_);
  or (_17069_, _17067_, _07142_);
  and (_17070_, _15512_, _07911_);
  or (_17071_, _17070_, _17059_);
  or (_17072_, _17071_, _06252_);
  and (_17073_, _07911_, \oc8051_golden_model_1.ACC [6]);
  or (_17074_, _17073_, _17059_);
  and (_17075_, _17074_, _07123_);
  nor (_17076_, _07123_, _10310_);
  or (_17077_, _17076_, _06251_);
  or (_17078_, _17077_, _17075_);
  and (_17079_, _17078_, _06476_);
  and (_17080_, _17079_, _17072_);
  nor (_17081_, _08547_, _10310_);
  and (_17082_, _15499_, _08547_);
  or (_17083_, _17082_, _17081_);
  and (_17084_, _17083_, _06475_);
  or (_17085_, _17084_, _06468_);
  or (_17086_, _17085_, _17080_);
  and (_17087_, _17086_, _17069_);
  or (_17088_, _17087_, _06466_);
  or (_17089_, _17074_, _06801_);
  and (_17090_, _17089_, _06484_);
  and (_17091_, _17090_, _17088_);
  and (_17092_, _15497_, _08547_);
  or (_17093_, _17092_, _17081_);
  and (_17094_, _17093_, _06483_);
  or (_17095_, _17094_, _17091_);
  and (_17096_, _17095_, _07164_);
  or (_17097_, _17081_, _15529_);
  and (_17098_, _17097_, _06461_);
  and (_17099_, _17098_, _17083_);
  or (_17100_, _17099_, _09487_);
  or (_17101_, _17100_, _17096_);
  nor (_17102_, _10026_, _10013_);
  nor (_17103_, _17102_, _10027_);
  or (_17104_, _17103_, _09494_);
  and (_17105_, _17104_, _06242_);
  and (_17106_, _17105_, _17101_);
  or (_17107_, _17081_, _15545_);
  and (_17108_, _17107_, _06241_);
  and (_17109_, _17108_, _17083_);
  or (_17110_, _17109_, _07187_);
  or (_17111_, _17110_, _17106_);
  and (_17112_, _17111_, _17068_);
  or (_17113_, _17112_, _07182_);
  and (_17114_, _09067_, _07911_);
  or (_17115_, _17059_, _07183_);
  or (_17116_, _17115_, _17114_);
  and (_17117_, _17116_, _06336_);
  and (_17118_, _17117_, _17113_);
  or (_17119_, _17118_, _17065_);
  and (_17120_, _17119_, _10052_);
  nor (_17121_, _17006_, _10372_);
  or (_17122_, _17121_, _10373_);
  and (_17123_, _17122_, _10378_);
  nor (_17124_, _17122_, _10378_);
  or (_17125_, _17124_, _17123_);
  or (_17126_, _17125_, _10398_);
  or (_17127_, _16775_, _10316_);
  and (_17128_, _17127_, _10046_);
  and (_17129_, _17128_, _17126_);
  or (_17130_, _17129_, _06371_);
  or (_17131_, _17130_, _17120_);
  and (_17132_, _17131_, _17062_);
  or (_17133_, _17132_, _06367_);
  and (_17134_, _15618_, _07911_);
  or (_17135_, _17134_, _17059_);
  or (_17136_, _17135_, _07218_);
  and (_17137_, _17136_, _07216_);
  and (_17138_, _17137_, _17133_);
  and (_17139_, _11202_, _07911_);
  or (_17140_, _17139_, _17059_);
  and (_17141_, _17140_, _06533_);
  or (_17142_, _17141_, _17138_);
  and (_17143_, _17142_, _07213_);
  or (_17144_, _17059_, _08109_);
  and (_17145_, _17061_, _06366_);
  and (_17146_, _17145_, _17144_);
  or (_17147_, _17146_, _17143_);
  and (_17148_, _17147_, _07210_);
  and (_17149_, _17074_, _06541_);
  and (_17150_, _17149_, _17144_);
  or (_17151_, _17150_, _06383_);
  or (_17152_, _17151_, _17148_);
  and (_17153_, _15615_, _07911_);
  or (_17154_, _17059_, _07231_);
  or (_17155_, _17154_, _17153_);
  and (_17156_, _17155_, _07229_);
  and (_17157_, _17156_, _17152_);
  nor (_17158_, _11201_, _09454_);
  or (_17159_, _17158_, _17059_);
  and (_17160_, _17159_, _06528_);
  or (_17161_, _17160_, _06563_);
  or (_17162_, _17161_, _17157_);
  or (_17163_, _17071_, _07241_);
  and (_17164_, _17163_, _06571_);
  and (_17165_, _17164_, _17162_);
  and (_17166_, _17093_, _06199_);
  or (_17167_, _17166_, _06188_);
  or (_17168_, _17167_, _17165_);
  and (_17169_, _15676_, _07911_);
  or (_17170_, _17059_, _06189_);
  or (_17171_, _17170_, _17169_);
  and (_17172_, _17171_, _01452_);
  and (_17173_, _17172_, _17168_);
  or (_17174_, _17173_, _17058_);
  and (_43768_, _17174_, _43223_);
  nor (_17175_, _01452_, _05997_);
  nand (_17176_, _10448_, _08506_);
  nand (_17177_, _11080_, _10854_);
  nor (_17178_, _10661_, _05997_);
  or (_17179_, _17178_, _10662_);
  or (_17180_, _17179_, _11022_);
  nand (_17181_, _11004_, _12544_);
  and (_17182_, _07129_, _06382_);
  nor (_17183_, _09342_, \oc8051_golden_model_1.ACC [0]);
  nor (_17184_, _17183_, _11179_);
  or (_17185_, _10930_, _17184_);
  nor (_17186_, _07325_, \oc8051_golden_model_1.ACC [0]);
  nor (_17187_, _11135_, _17186_);
  and (_17188_, _07053_, _05888_);
  nor (_17189_, _17188_, _06697_);
  not (_17190_, _17189_);
  and (_17191_, _17190_, _17187_);
  nor (_17192_, _07914_, _05997_);
  and (_17193_, _07914_, _07325_);
  or (_17194_, _17193_, _17192_);
  or (_17195_, _17194_, _07188_);
  nor (_17196_, _10591_, _05997_);
  or (_17197_, _17196_, _10592_);
  or (_17198_, _17197_, _06516_);
  and (_17199_, _17198_, _10543_);
  not (_17200_, _10682_);
  or (_17201_, _17200_, _07325_);
  nor (_17202_, _10687_, _07134_);
  or (_17203_, _17202_, _09342_);
  not (_17204_, _10704_);
  and (_17205_, _17204_, _07325_);
  or (_17206_, _06808_, \oc8051_golden_model_1.ACC [0]);
  nand (_17207_, _06808_, \oc8051_golden_model_1.ACC [0]);
  and (_17208_, _17207_, _17206_);
  and (_17209_, _17208_, _10704_);
  or (_17210_, _17209_, _10687_);
  or (_17211_, _17210_, _17205_);
  and (_17212_, _17211_, _05955_);
  or (_17213_, _17212_, _07134_);
  and (_17214_, _17213_, _06252_);
  and (_17215_, _17214_, _17203_);
  nor (_17216_, _08351_, _10538_);
  or (_17217_, _17216_, _17192_);
  and (_17218_, _17217_, _06251_);
  or (_17219_, _17218_, _06475_);
  or (_17220_, _17219_, _17215_);
  and (_17221_, _14341_, _08545_);
  nor (_17222_, _08545_, _05997_);
  or (_17223_, _17222_, _06476_);
  or (_17224_, _17223_, _17221_);
  and (_17225_, _17224_, _07142_);
  and (_17226_, _17225_, _17220_);
  and (_17227_, _17194_, _06468_);
  or (_17228_, _17227_, _10682_);
  or (_17229_, _17228_, _17226_);
  and (_17230_, _17229_, _17201_);
  or (_17231_, _17230_, _07153_);
  or (_17232_, _09342_, _07353_);
  and (_17233_, _17232_, _06801_);
  and (_17234_, _17233_, _17231_);
  and (_17235_, _08351_, _06466_);
  or (_17236_, _17235_, _10759_);
  or (_17237_, _17236_, _17234_);
  nand (_17238_, _10759_, _10087_);
  and (_17239_, _17238_, _17237_);
  or (_17240_, _17239_, _06483_);
  or (_17241_, _17192_, _06484_);
  and (_17242_, _17241_, _07164_);
  and (_17243_, _17242_, _17240_);
  and (_17244_, _17217_, _06461_);
  or (_17245_, _17244_, _09487_);
  or (_17246_, _17245_, _17243_);
  nand (_17247_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nand (_17248_, _17247_, _09487_);
  and (_17249_, _17248_, _10779_);
  and (_17250_, _17249_, _17246_);
  nor (_17251_, _10505_, _05997_);
  or (_17252_, _17251_, _10788_);
  and (_17253_, _17252_, _12236_);
  or (_17254_, _17253_, _10610_);
  or (_17255_, _17254_, _17250_);
  or (_17256_, _17179_, _10611_);
  and (_17257_, _17256_, _17255_);
  or (_17258_, _17257_, _06510_);
  and (_17259_, _17258_, _17199_);
  nor (_17260_, _12545_, _10854_);
  and (_17261_, _12545_, _10854_);
  or (_17262_, _17261_, _17260_);
  and (_17263_, _17262_, _10542_);
  or (_17264_, _17263_, _05976_);
  or (_17265_, _17264_, _17259_);
  or (_17266_, _06799_, _05977_);
  and (_17267_, _17266_, _06242_);
  and (_17268_, _17267_, _17265_);
  and (_17269_, _14372_, _08545_);
  or (_17270_, _17269_, _17222_);
  and (_17271_, _17270_, _06241_);
  or (_17272_, _17271_, _07187_);
  or (_17273_, _17272_, _17268_);
  and (_17274_, _17273_, _17195_);
  or (_17275_, _17274_, _07182_);
  and (_17276_, _09342_, _07914_);
  or (_17277_, _17192_, _07183_);
  or (_17278_, _17277_, _17276_);
  and (_17279_, _17278_, _06336_);
  and (_17280_, _17279_, _17275_);
  and (_17281_, _14427_, _07914_);
  or (_17282_, _17281_, _17192_);
  and (_17283_, _17282_, _05968_);
  or (_17284_, _17283_, _10046_);
  or (_17285_, _17284_, _17280_);
  nand (_17286_, _10398_, _10046_);
  and (_17287_, _17286_, _05975_);
  and (_17288_, _17287_, _17285_);
  and (_17289_, _06799_, _05935_);
  or (_17290_, _17289_, _06371_);
  or (_17291_, _17290_, _17288_);
  and (_17292_, _07914_, _08908_);
  or (_17293_, _17292_, _17192_);
  or (_17294_, _17293_, _07198_);
  and (_17295_, _17294_, _10905_);
  and (_17296_, _17295_, _17291_);
  and (_17297_, _10904_, _06799_);
  or (_17298_, _17297_, _10912_);
  or (_17299_, _17298_, _17296_);
  and (_17300_, _17189_, _10917_);
  and (_17301_, _17189_, _17187_);
  or (_17302_, _17301_, _17300_);
  and (_17303_, _17302_, _17299_);
  nor (_17304_, _17303_, _17191_);
  nor (_17305_, _10530_, _06924_);
  nor (_17306_, _17305_, _17304_);
  and (_17307_, _17305_, _17187_);
  or (_17308_, _17307_, _10929_);
  or (_17309_, _17308_, _17306_);
  and (_17310_, _17309_, _17185_);
  or (_17311_, _17310_, _06531_);
  nand (_17312_, _12527_, _06531_);
  and (_17313_, _17312_, _10534_);
  and (_17314_, _17313_, _17311_);
  and (_17315_, _12545_, _10533_);
  or (_17316_, _17315_, _06367_);
  or (_17317_, _17316_, _17314_);
  and (_17318_, _14442_, _07914_);
  or (_17319_, _17318_, _17192_);
  or (_17320_, _17319_, _07218_);
  and (_17321_, _17320_, _17317_);
  or (_17322_, _17321_, _06533_);
  nor (_17323_, _17192_, _07216_);
  nor (_17324_, _17323_, _12223_);
  and (_17325_, _17324_, _17322_);
  and (_17327_, _12223_, _11135_);
  nor (_17328_, _17327_, _17325_);
  nor (_17329_, _17328_, _12222_);
  and (_17330_, _12222_, _11135_);
  or (_17331_, _17330_, _17329_);
  and (_17332_, _17331_, _12220_);
  and (_17333_, _11135_, _12219_);
  or (_17334_, _17333_, _10960_);
  or (_17335_, _17334_, _17332_);
  or (_17336_, _10962_, _11179_);
  and (_17338_, _17336_, _06540_);
  and (_17339_, _17338_, _17335_);
  or (_17340_, _10966_, _11218_);
  and (_17341_, _17340_, _10968_);
  or (_17342_, _17341_, _17339_);
  or (_17343_, _10972_, _11256_);
  and (_17344_, _17343_, _07213_);
  and (_17345_, _17344_, _17342_);
  nand (_17346_, _17293_, _06366_);
  nor (_17347_, _17346_, _17216_);
  or (_17349_, _17347_, _07032_);
  or (_17350_, _17349_, _17345_);
  not (_17351_, _10980_);
  nand (_17352_, _17186_, _07032_);
  and (_17353_, _17352_, _17351_);
  and (_17354_, _17353_, _17350_);
  nor (_17355_, _17186_, _17351_);
  or (_17356_, _17355_, _07020_);
  or (_17357_, _17356_, _17354_);
  nand (_17358_, _17186_, _07020_);
  nand (_17360_, _17358_, _17357_);
  nor (_17361_, _17360_, _17182_);
  not (_17362_, _17186_);
  and (_17363_, _17362_, _17182_);
  or (_17364_, _17363_, _10998_);
  or (_17365_, _17364_, _17361_);
  nand (_17366_, _10998_, _17183_);
  and (_17367_, _17366_, _06527_);
  and (_17368_, _17367_, _17365_);
  nand (_17369_, _11007_, _12526_);
  and (_17371_, _17369_, _11006_);
  or (_17372_, _17371_, _17368_);
  and (_17373_, _17372_, _17181_);
  or (_17374_, _17373_, _06383_);
  and (_17375_, _14325_, _07914_);
  or (_17376_, _17192_, _07231_);
  or (_17377_, _17376_, _17375_);
  and (_17378_, _17377_, _10526_);
  and (_17379_, _17378_, _17374_);
  and (_17380_, _17252_, _10522_);
  and (_17382_, _17252_, _10525_);
  or (_17383_, _17382_, _10452_);
  or (_17384_, _17383_, _17380_);
  or (_17385_, _17384_, _17379_);
  and (_17386_, _17385_, _17180_);
  or (_17387_, _17386_, _06537_);
  or (_17388_, _17197_, _06538_);
  and (_17389_, _17388_, _11082_);
  and (_17390_, _17389_, _17387_);
  and (_17391_, _11050_, _17262_);
  or (_17392_, _17391_, _11080_);
  or (_17393_, _17392_, _17390_);
  and (_17394_, _17393_, _17177_);
  or (_17395_, _17394_, _06684_);
  not (_17396_, _06684_);
  nor (_17397_, _17187_, _17396_);
  nor (_17398_, _17397_, _06661_);
  and (_17399_, _17398_, _17395_);
  and (_17400_, _17187_, _06661_);
  and (_17401_, _06259_, _06347_);
  or (_17402_, _17401_, _17400_);
  or (_17403_, _17402_, _17399_);
  not (_17404_, _17401_);
  or (_17405_, _17404_, _17187_);
  and (_17406_, _17405_, _11160_);
  and (_17407_, _17406_, _17403_);
  and (_17408_, _11156_, _17184_);
  or (_17409_, _17408_, _06293_);
  or (_17410_, _17409_, _17407_);
  nand (_17411_, _12527_, _06293_);
  and (_17412_, _17411_, _10451_);
  and (_17413_, _17412_, _17410_);
  and (_17414_, _12545_, _10450_);
  or (_17415_, _17414_, _10448_);
  or (_17416_, _17415_, _17413_);
  and (_17417_, _17416_, _17176_);
  or (_17418_, _17417_, _06563_);
  or (_17419_, _17217_, _07241_);
  and (_17420_, _17419_, _11280_);
  and (_17421_, _17420_, _17418_);
  nor (_17422_, _11284_, _05997_);
  nor (_17423_, _17422_, _12991_);
  or (_17424_, _17423_, _17421_);
  nand (_17425_, _11284_, _05937_);
  and (_17426_, _17425_, _06571_);
  and (_17427_, _17426_, _17424_);
  and (_17428_, _17192_, _06199_);
  or (_17429_, _17428_, _06188_);
  or (_17430_, _17429_, _17427_);
  or (_17431_, _17217_, _06189_);
  and (_17432_, _17431_, _11303_);
  and (_17433_, _17432_, _17430_);
  and (_17434_, _11302_, _05997_);
  or (_17435_, _17434_, _11309_);
  or (_17436_, _17435_, _17433_);
  nand (_17437_, _11309_, _05937_);
  and (_17438_, _17437_, _01452_);
  and (_17439_, _17438_, _17436_);
  or (_17440_, _17439_, _17175_);
  and (_43769_, _17440_, _43223_);
  nor (_17441_, _01452_, _05937_);
  and (_17442_, _06810_, _06259_);
  and (_17443_, _07455_, _06259_);
  not (_17444_, _17443_);
  nor (_17445_, _11179_, _11178_);
  nor (_17446_, _17445_, _11180_);
  or (_17447_, _17446_, _17444_);
  or (_17448_, _11061_, _11060_);
  nor (_17449_, _11062_, _06538_);
  and (_17450_, _17449_, _17448_);
  and (_17451_, _07492_, _06365_);
  nor (_17452_, _07914_, _05937_);
  nor (_17453_, _10538_, _07120_);
  or (_17454_, _17453_, _17452_);
  or (_17455_, _17454_, _07188_);
  nor (_17456_, _08545_, _05937_);
  and (_17457_, _14510_, _08545_);
  or (_17458_, _17457_, _17456_);
  or (_17459_, _17456_, _14509_);
  and (_17460_, _17459_, _06461_);
  and (_17461_, _17460_, _17458_);
  nand (_17462_, _10682_, _07120_);
  nor (_17463_, _10722_, \oc8051_golden_model_1.PSW [6]);
  nor (_17464_, _17463_, \oc8051_golden_model_1.ACC [1]);
  and (_17465_, _17463_, \oc8051_golden_model_1.ACC [1]);
  nor (_17466_, _17465_, _17464_);
  nand (_17467_, _17466_, _10718_);
  or (_17468_, _17202_, _09297_);
  nor (_17469_, _10704_, _07120_);
  or (_17470_, _06808_, \oc8051_golden_model_1.ACC [1]);
  nand (_17471_, _06808_, \oc8051_golden_model_1.ACC [1]);
  and (_17472_, _17471_, _17470_);
  and (_17473_, _17472_, _10704_);
  or (_17474_, _17473_, _10687_);
  or (_17475_, _17474_, _17469_);
  and (_17476_, _17475_, _05955_);
  or (_17477_, _17476_, _07134_);
  and (_17478_, _17477_, _17468_);
  or (_17479_, _17478_, _06251_);
  or (_17480_, _07914_, \oc8051_golden_model_1.ACC [1]);
  and (_17481_, _14503_, _07914_);
  not (_17482_, _17481_);
  and (_17483_, _17482_, _17480_);
  or (_17484_, _17483_, _06252_);
  and (_17485_, _17484_, _17479_);
  or (_17486_, _17485_, _10718_);
  and (_17487_, _17486_, _17467_);
  or (_17488_, _17487_, _06475_);
  or (_17489_, _17458_, _06476_);
  and (_17490_, _17489_, _07142_);
  and (_17491_, _17490_, _17488_);
  and (_17492_, _17454_, _06468_);
  or (_17493_, _17492_, _10682_);
  or (_17494_, _17493_, _17491_);
  and (_17495_, _17494_, _17462_);
  or (_17496_, _17495_, _07153_);
  or (_17497_, _09297_, _07353_);
  and (_17498_, _17497_, _06801_);
  and (_17499_, _17498_, _17496_);
  nor (_17500_, _08301_, _06801_);
  or (_17501_, _17500_, _10759_);
  or (_17502_, _17501_, _17499_);
  nand (_17503_, _10759_, _10122_);
  and (_17504_, _17503_, _17502_);
  or (_17505_, _17504_, _06483_);
  and (_17506_, _14513_, _08545_);
  or (_17507_, _17506_, _17456_);
  or (_17508_, _17507_, _06484_);
  and (_17509_, _17508_, _07164_);
  and (_17510_, _17509_, _17505_);
  or (_17511_, _17510_, _17461_);
  and (_17512_, _17511_, _09494_);
  nor (_17513_, _09976_, _09975_);
  nor (_17514_, _17513_, _09977_);
  and (_17515_, _17514_, _09487_);
  or (_17516_, _17515_, _12236_);
  or (_17517_, _17516_, _17512_);
  nor (_17518_, _10453_, _05997_);
  or (_17519_, _17518_, _10504_);
  and (_17520_, _17519_, _11134_);
  nor (_17521_, _17519_, _11134_);
  or (_17522_, _17521_, _17520_);
  or (_17523_, _17522_, _10779_);
  and (_17524_, _17523_, _10611_);
  and (_17525_, _17524_, _17517_);
  nor (_17526_, _10654_, _05997_);
  or (_17527_, _17526_, _10660_);
  not (_17528_, _17527_);
  nand (_17529_, _17528_, _11178_);
  or (_17530_, _17528_, _11178_);
  and (_17531_, _17530_, _10610_);
  and (_17532_, _17531_, _17529_);
  or (_17533_, _17532_, _06510_);
  or (_17534_, _17533_, _17525_);
  nor (_17535_, _10544_, _05997_);
  or (_17536_, _17535_, _10590_);
  nor (_17537_, _17536_, _11217_);
  and (_17538_, _17536_, _11217_);
  or (_17539_, _17538_, _17537_);
  or (_17540_, _17539_, _06516_);
  and (_17541_, _17540_, _10543_);
  and (_17542_, _17541_, _17534_);
  and (_17543_, _06799_, _05997_);
  nor (_17544_, _17543_, _11255_);
  and (_17545_, _17543_, _11255_);
  or (_17546_, _17545_, _17544_);
  not (_17547_, _17546_);
  nand (_17548_, _17260_, _17547_);
  or (_17549_, _17260_, _17547_);
  and (_17550_, _17549_, _10542_);
  and (_17551_, _17550_, _17548_);
  or (_17552_, _17551_, _05976_);
  or (_17553_, _17552_, _17542_);
  nand (_17554_, _06155_, _05976_);
  and (_17555_, _17554_, _06242_);
  and (_17556_, _17555_, _17553_);
  or (_17557_, _17456_, _14553_);
  and (_17558_, _17557_, _06241_);
  and (_17559_, _17558_, _17458_);
  or (_17560_, _17559_, _07187_);
  or (_17561_, _17560_, _17556_);
  and (_17562_, _17561_, _17455_);
  or (_17563_, _17562_, _07182_);
  and (_17564_, _09297_, _07914_);
  or (_17565_, _17452_, _07183_);
  or (_17566_, _17565_, _17564_);
  and (_17567_, _17566_, _06336_);
  and (_17568_, _17567_, _17563_);
  or (_17569_, _14609_, _10538_);
  and (_17570_, _17480_, _05968_);
  and (_17571_, _17570_, _17569_);
  or (_17572_, _17571_, _10046_);
  or (_17573_, _17572_, _17568_);
  or (_17574_, _10305_, _10052_);
  and (_17575_, _17574_, _17573_);
  or (_17576_, _17575_, _05935_);
  nand (_17577_, _06155_, _05935_);
  and (_17578_, _17577_, _07198_);
  and (_17579_, _17578_, _17576_);
  nand (_17580_, _07914_, _07018_);
  and (_17581_, _17580_, _06371_);
  and (_17582_, _17581_, _17480_);
  or (_17583_, _17582_, _10904_);
  or (_17584_, _17583_, _17579_);
  nand (_17585_, _10904_, _06155_);
  and (_17586_, _17585_, _10917_);
  and (_17587_, _17586_, _17584_);
  and (_17588_, _10912_, _11134_);
  or (_17589_, _17588_, _17587_);
  and (_17590_, _17589_, _10920_);
  and (_17591_, _10919_, _11134_);
  or (_17592_, _17591_, _10924_);
  or (_17593_, _17592_, _17590_);
  and (_17594_, _10930_, _11134_);
  or (_17595_, _17594_, _12230_);
  and (_17596_, _17595_, _17593_);
  and (_17597_, _10929_, _11178_);
  or (_17598_, _17597_, _06531_);
  or (_17599_, _17598_, _17596_);
  or (_17600_, _11217_, _06532_);
  and (_17601_, _17600_, _17599_);
  or (_17602_, _17601_, _10533_);
  or (_17603_, _11255_, _10534_);
  and (_17604_, _17603_, _07218_);
  and (_17605_, _17604_, _17602_);
  or (_17606_, _14625_, _10538_);
  and (_17607_, _17606_, _06367_);
  and (_17608_, _17607_, _17480_);
  or (_17609_, _17608_, _06533_);
  or (_17610_, _17609_, _17605_);
  or (_17611_, _17452_, _07216_);
  and (_17612_, _17611_, _17610_);
  or (_17613_, _17612_, _17451_);
  nor (_17614_, _10692_, _05918_);
  nor (_17615_, _17614_, _10531_);
  not (_17616_, _17451_);
  or (_17617_, _17616_, _11132_);
  and (_17618_, _17617_, _17615_);
  and (_17619_, _17618_, _17613_);
  not (_17620_, _17615_);
  and (_17621_, _17620_, _11132_);
  or (_17622_, _17621_, _10960_);
  or (_17623_, _17622_, _17619_);
  or (_17624_, _10962_, _11176_);
  and (_17625_, _17624_, _06540_);
  and (_17626_, _17625_, _17623_);
  or (_17627_, _10966_, _11215_);
  and (_17628_, _17627_, _10968_);
  or (_17629_, _17628_, _17626_);
  or (_17630_, _10972_, _11253_);
  and (_17631_, _17630_, _07213_);
  and (_17632_, _17631_, _17629_);
  or (_17633_, _14623_, _10538_);
  and (_17634_, _17480_, _06366_);
  and (_17635_, _17634_, _17633_);
  or (_17636_, _17635_, _17632_);
  nor (_17637_, _10981_, _06654_);
  and (_17638_, _17637_, _17636_);
  nor (_17639_, _17637_, _11133_);
  or (_17640_, _17639_, _10988_);
  or (_17641_, _17640_, _17638_);
  nand (_17642_, _10988_, _11133_);
  and (_17643_, _17642_, _10993_);
  and (_17644_, _17643_, _17641_);
  nor (_17645_, _11133_, _10993_);
  or (_17646_, _17645_, _10998_);
  or (_17647_, _17646_, _17644_);
  nand (_17648_, _10998_, _11177_);
  and (_17649_, _17648_, _06527_);
  and (_17650_, _17649_, _17647_);
  nand (_17651_, _11007_, _11216_);
  and (_17652_, _17651_, _11006_);
  or (_17653_, _17652_, _17650_);
  nand (_17654_, _11004_, _11254_);
  and (_17655_, _17654_, _07231_);
  and (_17656_, _17655_, _17653_);
  or (_17657_, _17580_, _08302_);
  and (_17658_, _17480_, _06383_);
  and (_17659_, _17658_, _17657_);
  nor (_17660_, _17659_, _17656_);
  nor (_17661_, _17660_, _10525_);
  nor (_17662_, _10506_, _10503_);
  nor (_17663_, _17662_, _10507_);
  and (_17664_, _17663_, _10525_);
  or (_17665_, _17664_, _10522_);
  or (_17666_, _17665_, _17661_);
  and (_17667_, _07455_, _06380_);
  nor (_17668_, _17667_, _10522_);
  not (_17669_, _17667_);
  and (_17670_, _17663_, _17669_);
  or (_17671_, _17670_, _17668_);
  and (_17672_, _17671_, _17666_);
  and (_17673_, _06810_, _06380_);
  nor (_17674_, _11031_, _11030_);
  nor (_17675_, _17674_, _11032_);
  and (_17676_, _17675_, _10452_);
  or (_17677_, _17676_, _17673_);
  or (_17678_, _17677_, _17672_);
  not (_17679_, _17673_);
  or (_17680_, _17675_, _17679_);
  and (_17681_, _17680_, _06538_);
  and (_17682_, _17681_, _17678_);
  or (_17683_, _17682_, _17450_);
  and (_17684_, _17683_, _11082_);
  or (_17685_, _11091_, _11090_);
  nor (_17686_, _11092_, _11082_);
  and (_17687_, _17686_, _17685_);
  or (_17688_, _17687_, _11080_);
  or (_17689_, _17688_, _17684_);
  nand (_17690_, _11080_, _05997_);
  and (_17691_, _17690_, _12103_);
  and (_17692_, _17691_, _17689_);
  or (_17693_, _11135_, _11134_);
  nor (_17694_, _12103_, _11136_);
  and (_17695_, _17694_, _17693_);
  or (_17696_, _17695_, _17443_);
  or (_17697_, _17696_, _17692_);
  and (_17698_, _17697_, _17447_);
  or (_17699_, _17698_, _17442_);
  not (_17700_, _17442_);
  or (_17701_, _17446_, _17700_);
  and (_17702_, _17701_, _06295_);
  and (_17703_, _17702_, _17699_);
  nor (_17704_, _11218_, _11217_);
  nor (_17705_, _17704_, _11219_);
  or (_17706_, _17705_, _10450_);
  and (_17707_, _17706_, _12964_);
  or (_17708_, _17707_, _17703_);
  nor (_17709_, _11256_, _11255_);
  nor (_17710_, _17709_, _11257_);
  or (_17711_, _17710_, _10451_);
  and (_17712_, _17711_, _12966_);
  and (_17713_, _17712_, _17708_);
  and (_17714_, _10448_, \oc8051_golden_model_1.ACC [0]);
  or (_17715_, _17714_, _06563_);
  or (_17716_, _17715_, _17713_);
  or (_17717_, _17483_, _07241_);
  and (_17718_, _17717_, _11280_);
  and (_17719_, _17718_, _17716_);
  nor (_17720_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor (_17721_, _11310_, _17720_);
  nor (_17722_, _17721_, _11280_);
  or (_17723_, _17722_, _11284_);
  or (_17724_, _17723_, _17719_);
  nand (_17725_, _11284_, _10165_);
  and (_17726_, _17725_, _06571_);
  and (_17727_, _17726_, _17724_);
  and (_17728_, _17507_, _06199_);
  or (_17729_, _17728_, _06188_);
  or (_17730_, _17729_, _17727_);
  or (_17731_, _17481_, _17452_);
  or (_17732_, _17731_, _06189_);
  and (_17733_, _17732_, _11303_);
  and (_17734_, _17733_, _17730_);
  nor (_17735_, _17721_, _11309_);
  nor (_17736_, _17735_, _13013_);
  or (_17737_, _17736_, _17734_);
  nand (_17738_, _11309_, _10165_);
  and (_17739_, _17738_, _01452_);
  and (_17740_, _17739_, _17737_);
  or (_17741_, _17740_, _17441_);
  and (_43771_, _17741_, _43223_);
  nor (_17742_, _01452_, _10165_);
  nand (_17743_, _10448_, _05937_);
  nand (_17744_, _11004_, _11251_);
  or (_17745_, _11214_, _06532_);
  and (_17746_, _17745_, _10534_);
  and (_17747_, _06361_, _05888_);
  not (_17748_, _17747_);
  nor (_17749_, _10905_, _06750_);
  nand (_17750_, _06750_, _05935_);
  nor (_17751_, _07914_, _10165_);
  nor (_17752_, _10538_, _07578_);
  or (_17753_, _17752_, _17751_);
  or (_17754_, _17753_, _07188_);
  and (_17755_, _06810_, _05969_);
  nand (_17756_, _10682_, _07578_);
  nor (_17757_, _17464_, _10165_);
  and (_17758_, _10721_, \oc8051_golden_model_1.PSW [6]);
  nor (_17759_, _17758_, _17757_);
  nand (_17760_, _17759_, _10718_);
  or (_17761_, _17202_, _09251_);
  nor (_17762_, _10704_, _07578_);
  or (_17763_, _06808_, \oc8051_golden_model_1.ACC [2]);
  nand (_17764_, _06808_, \oc8051_golden_model_1.ACC [2]);
  and (_17765_, _17764_, _17763_);
  and (_17766_, _17765_, _10704_);
  or (_17767_, _17766_, _10687_);
  or (_17768_, _17767_, _17762_);
  and (_17769_, _17768_, _05955_);
  or (_17770_, _17769_, _07134_);
  and (_17771_, _17770_, _17761_);
  or (_17772_, _17771_, _06251_);
  and (_17773_, _14712_, _07914_);
  or (_17774_, _17773_, _17751_);
  or (_17775_, _17774_, _06252_);
  and (_17776_, _17775_, _17772_);
  or (_17777_, _17776_, _10718_);
  and (_17778_, _17777_, _17760_);
  or (_17779_, _17778_, _06475_);
  nor (_17780_, _08545_, _10165_);
  and (_17781_, _14702_, _08545_);
  or (_17782_, _17781_, _17780_);
  or (_17783_, _17782_, _06476_);
  and (_17784_, _17783_, _07142_);
  and (_17785_, _17784_, _17779_);
  and (_17786_, _17753_, _06468_);
  or (_17787_, _17786_, _10682_);
  or (_17788_, _17787_, _17785_);
  and (_17789_, _17788_, _17756_);
  or (_17790_, _17789_, _07153_);
  or (_17791_, _09251_, _07353_);
  and (_17792_, _17791_, _06801_);
  and (_17793_, _17792_, _17790_);
  nor (_17794_, _08396_, _06801_);
  or (_17795_, _17794_, _10759_);
  or (_17796_, _17795_, _17793_);
  nand (_17797_, _10759_, _10068_);
  and (_17798_, _17797_, _17796_);
  or (_17799_, _17798_, _06483_);
  and (_17800_, _14706_, _08545_);
  or (_17801_, _17800_, _17780_);
  or (_17802_, _17801_, _06484_);
  and (_17803_, _17802_, _07164_);
  and (_17804_, _17803_, _17799_);
  or (_17805_, _17780_, _14739_);
  and (_17806_, _17782_, _06461_);
  and (_17807_, _17806_, _17805_);
  or (_17808_, _17807_, _09487_);
  or (_17809_, _17808_, _17804_);
  nor (_17810_, _09979_, _09977_);
  or (_17811_, _17810_, _09980_);
  nand (_17812_, _17811_, _09487_);
  and (_17813_, _17812_, _10779_);
  and (_17814_, _17813_, _17809_);
  and (_17815_, _07455_, _05969_);
  and (_17816_, _07120_, \oc8051_golden_model_1.ACC [1]);
  and (_17817_, _07325_, _05997_);
  nor (_17818_, _17817_, _11134_);
  nor (_17819_, _17818_, _17816_);
  nor (_17820_, _11131_, _17819_);
  and (_17821_, _11131_, _17819_);
  nor (_17822_, _17821_, _17820_);
  nor (_17823_, _17187_, _11134_);
  and (_17824_, _17823_, \oc8051_golden_model_1.PSW [7]);
  or (_17825_, _17824_, _17822_);
  nand (_17826_, _17824_, _17822_);
  and (_17827_, _17826_, _12236_);
  and (_17828_, _17827_, _17825_);
  or (_17829_, _17828_, _17815_);
  or (_17830_, _17829_, _17814_);
  nor (_17831_, _09297_, _05937_);
  and (_17832_, _09342_, _05997_);
  nor (_17833_, _17832_, _11178_);
  nor (_17834_, _17833_, _17831_);
  nor (_17835_, _11175_, _17834_);
  and (_17836_, _11175_, _17834_);
  nor (_17837_, _17836_, _17835_);
  nor (_17838_, _17184_, _11178_);
  not (_17839_, _17838_);
  or (_17840_, _17839_, _17837_);
  and (_17841_, _17840_, \oc8051_golden_model_1.PSW [7]);
  nor (_17842_, _17837_, \oc8051_golden_model_1.PSW [7]);
  nor (_17843_, _17842_, _17841_);
  and (_17844_, _17839_, _17837_);
  or (_17845_, _17844_, _17843_);
  or (_17846_, _17845_, _10611_);
  and (_17847_, _17846_, _17830_);
  or (_17848_, _17847_, _17755_);
  not (_17849_, _17755_);
  or (_17850_, _17845_, _17849_);
  and (_17851_, _17850_, _06516_);
  and (_17852_, _17851_, _17848_);
  and (_17853_, _08301_, \oc8051_golden_model_1.ACC [1]);
  and (_17854_, _08351_, _05997_);
  nor (_17855_, _14096_, _17854_);
  nor (_17856_, _17855_, _17853_);
  nor (_17857_, _11214_, _17856_);
  and (_17858_, _11214_, _17856_);
  nor (_17859_, _17858_, _17857_);
  not (_17860_, _17859_);
  and (_17861_, _12528_, \oc8051_golden_model_1.PSW [7]);
  or (_17862_, _17861_, _17860_);
  nand (_17863_, _17861_, _17860_);
  nand (_17864_, _17863_, _17862_);
  and (_17865_, _17864_, _06510_);
  or (_17866_, _17865_, _10542_);
  or (_17867_, _17866_, _17852_);
  nor (_17868_, _17544_, _14124_);
  nor (_17869_, _11252_, _17868_);
  and (_17870_, _11252_, _17868_);
  nor (_17871_, _17870_, _17869_);
  and (_17872_, _12546_, \oc8051_golden_model_1.PSW [7]);
  nand (_17873_, _17872_, _17871_);
  or (_17874_, _17872_, _17871_);
  and (_17875_, _17874_, _17873_);
  or (_17876_, _17875_, _10543_);
  and (_17877_, _17876_, _17867_);
  or (_17878_, _17877_, _05976_);
  nand (_17879_, _06750_, _05976_);
  and (_17880_, _17879_, _06242_);
  and (_17881_, _17880_, _17878_);
  or (_17882_, _17780_, _14703_);
  and (_17883_, _17882_, _06241_);
  and (_17884_, _17883_, _17782_);
  or (_17885_, _17884_, _07187_);
  or (_17886_, _17885_, _17881_);
  and (_17887_, _17886_, _17754_);
  or (_17888_, _17887_, _07182_);
  and (_17889_, _09251_, _07914_);
  or (_17890_, _17751_, _07183_);
  or (_17891_, _17890_, _17889_);
  and (_17892_, _17891_, _06336_);
  and (_17893_, _17892_, _17888_);
  and (_17894_, _14808_, _07914_);
  or (_17895_, _17894_, _17751_);
  and (_17896_, _17895_, _05968_);
  or (_17897_, _17896_, _10046_);
  or (_17898_, _17897_, _17893_);
  or (_17899_, _10242_, _10052_);
  and (_17900_, _17899_, _17898_);
  or (_17901_, _17900_, _05935_);
  and (_17902_, _17901_, _17750_);
  or (_17903_, _17902_, _06371_);
  and (_17904_, _07914_, _08945_);
  or (_17905_, _17904_, _17751_);
  or (_17906_, _17905_, _07198_);
  and (_17907_, _17906_, _10905_);
  and (_17908_, _17907_, _17903_);
  or (_17909_, _17908_, _17749_);
  and (_17910_, _17909_, _12231_);
  not (_17911_, _12231_);
  and (_17912_, _17911_, _11131_);
  or (_17913_, _17912_, _17910_);
  and (_17914_, _17913_, _17748_);
  and (_17915_, _05888_, _06348_);
  and (_17916_, _17747_, _11131_);
  or (_17917_, _17916_, _17915_);
  or (_17918_, _17917_, _17914_);
  not (_17919_, _17915_);
  or (_17920_, _11131_, _17919_);
  and (_17921_, _17920_, _10930_);
  and (_17922_, _17921_, _17918_);
  and (_17923_, _10929_, _11175_);
  or (_17924_, _17923_, _06531_);
  or (_17925_, _17924_, _17922_);
  and (_17926_, _17925_, _17746_);
  and (_17927_, _11252_, _10533_);
  or (_17928_, _17927_, _06367_);
  or (_17929_, _17928_, _17926_);
  and (_17930_, _14824_, _07914_);
  or (_17931_, _17930_, _17751_);
  or (_17932_, _17931_, _07218_);
  and (_17933_, _17932_, _17929_);
  or (_17934_, _17933_, _06533_);
  or (_17935_, _17751_, _07216_);
  and (_17936_, _17935_, _12225_);
  and (_17937_, _17936_, _17934_);
  not (_17938_, _12225_);
  and (_17939_, _17938_, _11129_);
  or (_17940_, _17939_, _10960_);
  or (_17941_, _17940_, _17937_);
  or (_17942_, _10962_, _11173_);
  and (_17943_, _17942_, _06540_);
  and (_17944_, _17943_, _17941_);
  or (_17945_, _10966_, _11212_);
  and (_17946_, _17945_, _10968_);
  or (_17947_, _17946_, _17944_);
  or (_17948_, _10972_, _11250_);
  and (_17949_, _17948_, _07213_);
  and (_17951_, _17949_, _17947_);
  nand (_17952_, _17905_, _06366_);
  nor (_17953_, _17952_, _11213_);
  or (_17954_, _17953_, _17951_);
  and (_17955_, _17954_, _17637_);
  nor (_17956_, _17637_, _11130_);
  or (_17957_, _17956_, _10988_);
  or (_17958_, _17957_, _17955_);
  nand (_17959_, _10988_, _11130_);
  and (_17960_, _17959_, _10993_);
  and (_17961_, _17960_, _17958_);
  nor (_17962_, _11130_, _10993_);
  or (_17963_, _17962_, _10998_);
  or (_17964_, _17963_, _17961_);
  nand (_17965_, _10998_, _11174_);
  and (_17966_, _17965_, _06527_);
  and (_17967_, _17966_, _17964_);
  nand (_17968_, _11007_, _11213_);
  and (_17969_, _17968_, _11006_);
  or (_17970_, _17969_, _17967_);
  and (_17971_, _17970_, _17744_);
  or (_17972_, _17971_, _06383_);
  and (_17973_, _14821_, _07914_);
  or (_17974_, _17751_, _07231_);
  or (_17975_, _17974_, _17973_);
  and (_17976_, _17975_, _10526_);
  and (_17977_, _17976_, _17972_);
  and (_17978_, _10508_, _10496_);
  nor (_17979_, _17978_, _10509_);
  and (_17980_, _17979_, _11014_);
  or (_17981_, _17980_, _17667_);
  or (_17982_, _17981_, _17977_);
  and (_17983_, _11033_, _10652_);
  nor (_17984_, _17983_, _11034_);
  or (_17985_, _17984_, _11022_);
  and (_17986_, _17985_, _17679_);
  and (_17987_, _17986_, _17982_);
  nand (_17988_, _17984_, _17673_);
  nand (_17989_, _17988_, _06538_);
  or (_17990_, _17989_, _17987_);
  and (_17991_, _11063_, _10584_);
  nor (_17992_, _17991_, _11064_);
  or (_17993_, _17992_, _06538_);
  and (_17994_, _17993_, _11082_);
  and (_17995_, _17994_, _17990_);
  and (_17996_, _11093_, _10847_);
  nor (_17997_, _17996_, _11094_);
  and (_17998_, _17997_, _11050_);
  or (_17999_, _17998_, _11080_);
  or (_18000_, _17999_, _17995_);
  nand (_18001_, _11080_, _05937_);
  and (_18002_, _18001_, _12103_);
  and (_18003_, _18002_, _18000_);
  or (_18004_, _11138_, _11131_);
  nor (_18005_, _12103_, _11139_);
  and (_18006_, _18005_, _18004_);
  or (_18007_, _18006_, _17443_);
  or (_18008_, _18007_, _18003_);
  nor (_18009_, _11182_, _11175_);
  nor (_18010_, _18009_, _11183_);
  and (_18011_, _18010_, _05932_);
  or (_18012_, _18011_, _11160_);
  and (_18013_, _18012_, _18008_);
  and (_18014_, _18010_, _17442_);
  or (_18015_, _18014_, _18013_);
  or (_18016_, _18015_, _06293_);
  nor (_18017_, _11221_, _11214_);
  nor (_18018_, _18017_, _11222_);
  or (_18019_, _18018_, _06295_);
  and (_18020_, _18019_, _10451_);
  and (_18021_, _18020_, _18016_);
  or (_18022_, _11259_, _11252_);
  nor (_18023_, _11260_, _10451_);
  and (_18024_, _18023_, _18022_);
  or (_18025_, _18024_, _10448_);
  or (_18026_, _18025_, _18021_);
  and (_18027_, _18026_, _17743_);
  or (_18028_, _18027_, _06563_);
  or (_18029_, _17774_, _07241_);
  and (_18030_, _18029_, _11280_);
  and (_18031_, _18030_, _18028_);
  nor (_18032_, _17720_, _10165_);
  or (_18033_, _18032_, _11285_);
  and (_18034_, _18033_, _11279_);
  or (_18035_, _18034_, _11284_);
  or (_18036_, _18035_, _18031_);
  nand (_18037_, _11284_, _10218_);
  and (_18038_, _18037_, _06571_);
  and (_18039_, _18038_, _18036_);
  and (_18040_, _17801_, _06199_);
  or (_18041_, _18040_, _06188_);
  or (_18042_, _18041_, _18039_);
  and (_18043_, _14884_, _07914_);
  or (_18044_, _18043_, _17751_);
  or (_18045_, _18044_, _06189_);
  and (_18046_, _18045_, _11303_);
  and (_18047_, _18046_, _18042_);
  nor (_18048_, _11310_, \oc8051_golden_model_1.ACC [2]);
  nor (_18049_, _18048_, _11311_);
  and (_18050_, _18049_, _11302_);
  or (_18051_, _18050_, _11309_);
  or (_18052_, _18051_, _18047_);
  nand (_18053_, _11309_, _10218_);
  and (_18054_, _18053_, _01452_);
  and (_18055_, _18054_, _18052_);
  or (_18056_, _18055_, _17742_);
  and (_43772_, _18056_, _43223_);
  nor (_18057_, _01452_, _10218_);
  nand (_18058_, _10448_, _10165_);
  nor (_18059_, _11223_, _12523_);
  and (_18060_, _11223_, _12523_);
  or (_18061_, _18060_, _18059_);
  and (_18062_, _18061_, _06293_);
  and (_18063_, _10510_, _10490_);
  nor (_18064_, _18063_, _10511_);
  or (_18065_, _18064_, _10526_);
  or (_18066_, _11210_, _06540_);
  and (_18067_, _06810_, _05888_);
  nand (_18068_, _06292_, _05935_);
  nor (_18069_, _07914_, _10218_);
  nor (_18070_, _10538_, _07713_);
  or (_18071_, _18070_, _18069_);
  or (_18072_, _18071_, _07188_);
  nor (_18073_, _08545_, _10218_);
  and (_18074_, _14906_, _08545_);
  or (_18075_, _18074_, _18073_);
  or (_18076_, _18073_, _14931_);
  and (_18077_, _18076_, _06461_);
  and (_18078_, _18077_, _18075_);
  nand (_18079_, _10682_, _07713_);
  and (_18080_, _14898_, _07914_);
  or (_18081_, _18080_, _18069_);
  and (_18082_, _18081_, _06251_);
  or (_18083_, _17202_, _09205_);
  nor (_18084_, _10704_, _07713_);
  nor (_18085_, _06808_, _10218_);
  and (_18086_, _06808_, _10218_);
  or (_18087_, _18086_, _18085_);
  and (_18088_, _18087_, _10704_);
  or (_18089_, _18088_, _10687_);
  or (_18090_, _18089_, _18084_);
  and (_18091_, _18090_, _05955_);
  or (_18092_, _18091_, _07134_);
  and (_18093_, _18092_, _06252_);
  and (_18094_, _18093_, _18083_);
  or (_18095_, _18094_, _18082_);
  and (_18096_, _18095_, _10719_);
  not (_18097_, \oc8051_golden_model_1.PSW [6]);
  nor (_18098_, _10721_, _18097_);
  nor (_18099_, _18098_, \oc8051_golden_model_1.ACC [3]);
  nor (_18100_, _18099_, _10722_);
  and (_18101_, _18100_, _10718_);
  or (_18102_, _18101_, _06475_);
  or (_18103_, _18102_, _18096_);
  or (_18104_, _18075_, _06476_);
  and (_18105_, _18104_, _07142_);
  and (_18106_, _18105_, _18103_);
  and (_18107_, _18071_, _06468_);
  or (_18108_, _18107_, _10682_);
  or (_18109_, _18108_, _18106_);
  and (_18110_, _18109_, _18079_);
  or (_18111_, _18110_, _07153_);
  or (_18112_, _09205_, _07353_);
  and (_18113_, _18112_, _06801_);
  and (_18114_, _18113_, _18111_);
  nor (_18115_, _08256_, _06801_);
  or (_18116_, _18115_, _10759_);
  or (_18117_, _18116_, _18114_);
  nand (_18118_, _10759_, _08506_);
  and (_18119_, _18118_, _18117_);
  or (_18120_, _18119_, _06483_);
  and (_18121_, _14904_, _08545_);
  or (_18122_, _18121_, _18073_);
  or (_18123_, _18122_, _06484_);
  and (_18124_, _18123_, _07164_);
  and (_18125_, _18124_, _18120_);
  or (_18126_, _18125_, _18078_);
  and (_18127_, _18126_, _09494_);
  or (_18128_, _09982_, _09980_);
  nor (_18129_, _09983_, _09494_);
  and (_18130_, _18129_, _18128_);
  or (_18131_, _18130_, _12236_);
  or (_18132_, _18131_, _18127_);
  and (_18133_, _07578_, \oc8051_golden_model_1.ACC [2]);
  nor (_18134_, _17820_, _18133_);
  nor (_18135_, _11127_, _11128_);
  nor (_18136_, _18135_, _18134_);
  and (_18137_, _18135_, _18134_);
  nor (_18138_, _18137_, _18136_);
  and (_18139_, _18138_, \oc8051_golden_model_1.PSW [7]);
  nor (_18140_, _18138_, \oc8051_golden_model_1.PSW [7]);
  nor (_18141_, _18140_, _18139_);
  and (_18142_, _17822_, \oc8051_golden_model_1.PSW [7]);
  nor (_18143_, _17823_, _10854_);
  nor (_18144_, _18143_, _18142_);
  not (_18145_, _18144_);
  and (_18146_, _18145_, _18141_);
  nor (_18147_, _18145_, _18141_);
  nor (_18148_, _18147_, _18146_);
  or (_18149_, _18148_, _10779_);
  and (_18150_, _18149_, _18132_);
  or (_18151_, _18150_, _10610_);
  nor (_18152_, _09251_, _10165_);
  nor (_18153_, _17835_, _18152_);
  nor (_18154_, _11172_, _11171_);
  nor (_18155_, _18154_, _18153_);
  and (_18156_, _18154_, _18153_);
  nor (_18157_, _18156_, _18155_);
  and (_18158_, _18157_, \oc8051_golden_model_1.PSW [7]);
  nor (_18159_, _18157_, \oc8051_golden_model_1.PSW [7]);
  nor (_18160_, _18159_, _18158_);
  nand (_18161_, _18160_, _17841_);
  or (_18162_, _18160_, _17841_);
  and (_18163_, _18162_, _18161_);
  or (_18164_, _18163_, _10611_);
  and (_18165_, _18164_, _06516_);
  and (_18166_, _18165_, _18151_);
  and (_18167_, _12529_, \oc8051_golden_model_1.PSW [7]);
  and (_18168_, _08396_, \oc8051_golden_model_1.ACC [2]);
  nor (_18169_, _17857_, _18168_);
  nor (_18170_, _12523_, _18169_);
  and (_18171_, _12523_, _18169_);
  nor (_18172_, _18171_, _18170_);
  and (_18173_, _17863_, _18172_);
  or (_18174_, _18173_, _10542_);
  or (_18175_, _18174_, _18167_);
  and (_18176_, _18175_, _12589_);
  or (_18177_, _18176_, _18166_);
  and (_18178_, _12547_, \oc8051_golden_model_1.PSW [7]);
  and (_18179_, _06750_, \oc8051_golden_model_1.ACC [2]);
  nor (_18180_, _17869_, _18179_);
  nor (_18181_, _12542_, _18180_);
  and (_18182_, _12542_, _18180_);
  nor (_18183_, _18182_, _18181_);
  not (_18184_, _12546_);
  or (_18185_, _18184_, _17871_);
  or (_18186_, _18185_, _10854_);
  and (_18187_, _18186_, _18183_);
  or (_18188_, _18187_, _10543_);
  or (_18189_, _18188_, _18178_);
  and (_18190_, _18189_, _18177_);
  or (_18191_, _18190_, _05976_);
  nand (_18192_, _06292_, _05976_);
  and (_18193_, _18192_, _06242_);
  and (_18194_, _18193_, _18191_);
  or (_18195_, _18073_, _14947_);
  and (_18196_, _18195_, _06241_);
  and (_18197_, _18196_, _18075_);
  or (_18198_, _18197_, _07187_);
  or (_18199_, _18198_, _18194_);
  and (_18200_, _18199_, _18072_);
  or (_18201_, _18200_, _07182_);
  and (_18202_, _09205_, _07914_);
  or (_18203_, _18069_, _07183_);
  or (_18204_, _18203_, _18202_);
  and (_18205_, _18204_, _06336_);
  and (_18206_, _18205_, _18201_);
  and (_18207_, _15003_, _07914_);
  or (_18208_, _18207_, _18069_);
  and (_18209_, _18208_, _05968_);
  or (_18210_, _18209_, _10046_);
  or (_18211_, _18210_, _18206_);
  or (_18212_, _10187_, _10052_);
  and (_18213_, _18212_, _18211_);
  or (_18214_, _18213_, _05935_);
  and (_18215_, _18214_, _18068_);
  or (_18216_, _18215_, _06371_);
  and (_18217_, _07914_, _08872_);
  nor (_18218_, _18217_, _18069_);
  nand (_18219_, _18218_, _06371_);
  and (_18220_, _18219_, _10905_);
  and (_18221_, _18220_, _18216_);
  or (_18222_, _10905_, _06292_);
  and (_18223_, _05888_, _06339_);
  not (_18224_, _18223_);
  and (_18225_, _06699_, _18224_);
  and (_18226_, _06352_, _05888_);
  and (_18227_, _05888_, _06347_);
  nor (_18228_, _18227_, _18226_);
  and (_18229_, _18228_, _18225_);
  nand (_18230_, _18229_, _18222_);
  or (_18231_, _18230_, _18221_);
  nand (_18232_, _10929_, _05932_);
  or (_18233_, _18229_, _18135_);
  and (_18234_, _18233_, _18232_);
  and (_18235_, _18234_, _18231_);
  and (_18236_, _07455_, _05888_);
  and (_18237_, _18236_, _18154_);
  nor (_18238_, _18237_, _18235_);
  nor (_18239_, _18238_, _18067_);
  and (_18240_, _18154_, _18067_);
  or (_18241_, _18240_, _06531_);
  or (_18242_, _18241_, _18239_);
  or (_18243_, _12523_, _06532_);
  and (_18244_, _18243_, _10534_);
  and (_18245_, _18244_, _18242_);
  and (_18246_, _12542_, _10533_);
  or (_18247_, _18246_, _06367_);
  or (_18248_, _18247_, _18245_);
  and (_18249_, _15018_, _07914_);
  or (_18250_, _18249_, _18069_);
  or (_18251_, _18250_, _07218_);
  and (_18252_, _18251_, _18248_);
  or (_18253_, _18252_, _06533_);
  or (_18254_, _18069_, _07216_);
  nor (_18255_, _12223_, _07033_);
  and (_18256_, _18255_, _18254_);
  and (_18257_, _18256_, _18253_);
  and (_18258_, _07129_, _06365_);
  not (_18259_, _18255_);
  and (_18260_, _18259_, _11127_);
  or (_18261_, _18260_, _18258_);
  or (_18262_, _18261_, _18257_);
  not (_18263_, _18258_);
  or (_18264_, _11127_, _18263_);
  and (_18265_, _18264_, _10962_);
  and (_18266_, _18265_, _18262_);
  and (_18267_, _10960_, _11171_);
  or (_18268_, _18267_, _06539_);
  or (_18269_, _18268_, _18266_);
  and (_18270_, _18269_, _18066_);
  or (_18271_, _18270_, _10966_);
  or (_18272_, _10972_, _11248_);
  and (_18273_, _18272_, _07213_);
  nand (_18274_, _18273_, _18271_);
  or (_18275_, _18218_, _07213_);
  or (_18276_, _18275_, _11211_);
  and (_18277_, _18276_, _18274_);
  or (_18278_, _18277_, _07032_);
  nand (_18279_, _11128_, _05730_);
  and (_18280_, _18279_, _06654_);
  nor (_18281_, _18280_, _07020_);
  nand (_18282_, _18281_, _18278_);
  or (_18283_, _07020_, _10980_);
  and (_18284_, _18283_, _11128_);
  nor (_18285_, _18284_, _17182_);
  and (_18286_, _18285_, _18282_);
  not (_18287_, _11128_);
  and (_18288_, _18287_, _17182_);
  or (_18289_, _18288_, _10998_);
  or (_18290_, _18289_, _18286_);
  nand (_18291_, _10998_, _11172_);
  and (_18292_, _18291_, _06527_);
  and (_18293_, _18292_, _18290_);
  nand (_18294_, _11007_, _11211_);
  and (_18295_, _18294_, _11006_);
  or (_18296_, _18295_, _18293_);
  nand (_18297_, _11004_, _11249_);
  and (_18298_, _18297_, _07231_);
  and (_18299_, _18298_, _18296_);
  and (_18300_, _15015_, _07914_);
  or (_18301_, _18300_, _18069_);
  and (_18302_, _18301_, _06383_);
  or (_18303_, _18302_, _11014_);
  or (_18304_, _18303_, _18299_);
  and (_18305_, _18304_, _18065_);
  or (_18306_, _18305_, _10452_);
  and (_18307_, _11035_, _10645_);
  nor (_18308_, _18307_, _11036_);
  or (_18309_, _18308_, _11022_);
  and (_18310_, _18309_, _06538_);
  and (_18311_, _18310_, _18306_);
  and (_18312_, _11065_, _10579_);
  nor (_18313_, _18312_, _11066_);
  or (_18314_, _18313_, _11050_);
  and (_18315_, _18314_, _11052_);
  or (_18316_, _18315_, _18311_);
  and (_18317_, _11095_, _10842_);
  nor (_18318_, _18317_, _11096_);
  or (_18319_, _18318_, _11082_);
  and (_18320_, _18319_, _11081_);
  and (_18321_, _18320_, _18316_);
  and (_18322_, _11080_, \oc8051_golden_model_1.ACC [2]);
  or (_18323_, _18322_, _12104_);
  or (_18324_, _18323_, _18321_);
  and (_18325_, _11140_, _18135_);
  nor (_18326_, _11140_, _18135_);
  or (_18327_, _18326_, _12103_);
  or (_18328_, _18327_, _18325_);
  and (_18329_, _18328_, _18324_);
  or (_18330_, _18329_, _11156_);
  and (_18331_, _11184_, _18154_);
  nor (_18332_, _11184_, _18154_);
  or (_18333_, _18332_, _18331_);
  or (_18334_, _18333_, _11160_);
  and (_18335_, _18334_, _06295_);
  and (_18336_, _18335_, _18330_);
  or (_18337_, _18336_, _18062_);
  and (_18338_, _18337_, _10451_);
  and (_18339_, _11261_, _12542_);
  nor (_18340_, _11261_, _12542_);
  or (_18341_, _18340_, _18339_);
  and (_18342_, _18341_, _10450_);
  or (_18343_, _18342_, _10448_);
  or (_18344_, _18343_, _18338_);
  and (_18345_, _18344_, _18058_);
  or (_18346_, _18345_, _06563_);
  or (_18347_, _18081_, _07241_);
  and (_18348_, _18347_, _11280_);
  and (_18349_, _18348_, _18346_);
  nor (_18350_, _11285_, _10218_);
  or (_18351_, _18350_, _11286_);
  nor (_18352_, _18351_, _11284_);
  nor (_18353_, _18352_, _12991_);
  or (_18354_, _18353_, _18349_);
  nand (_18355_, _11284_, _10087_);
  and (_18356_, _18355_, _06571_);
  and (_18357_, _18356_, _18354_);
  and (_18358_, _18122_, _06199_);
  or (_18359_, _18358_, _06188_);
  or (_18360_, _18359_, _18357_);
  and (_18361_, _15075_, _07914_);
  or (_18362_, _18361_, _18069_);
  or (_18363_, _18362_, _06189_);
  and (_18364_, _18363_, _11303_);
  and (_18365_, _18364_, _18360_);
  nor (_18366_, _11311_, \oc8051_golden_model_1.ACC [3]);
  nor (_18367_, _18366_, _11312_);
  and (_18368_, _18367_, _11302_);
  or (_18369_, _18368_, _11309_);
  or (_18370_, _18369_, _18365_);
  nand (_18371_, _11309_, _10087_);
  and (_18372_, _18371_, _01452_);
  and (_18373_, _18372_, _18370_);
  or (_18374_, _18373_, _18057_);
  and (_43773_, _18374_, _43223_);
  nor (_18375_, _01452_, _10087_);
  nand (_18376_, _10448_, _10218_);
  or (_18377_, _11225_, _11209_);
  and (_18378_, _18377_, _11226_);
  or (_18379_, _18378_, _06295_);
  and (_18380_, _18379_, _10451_);
  nand (_18381_, _11004_, _11246_);
  not (_18382_, _06654_);
  or (_18383_, _11124_, _18382_);
  or (_18384_, _11209_, _06532_);
  and (_18385_, _18384_, _10534_);
  and (_18386_, _05888_, _06817_);
  not (_18387_, _06698_);
  nor (_18388_, _11126_, _18387_);
  nor (_18389_, _18388_, _06697_);
  nand (_18390_, _06230_, _05935_);
  nor (_18391_, _07914_, _10087_);
  nor (_18392_, _08494_, _10538_);
  or (_18393_, _18392_, _18391_);
  or (_18394_, _18393_, _07188_);
  nor (_18395_, _12547_, _10854_);
  or (_18396_, _18180_, _14118_);
  and (_18397_, _18396_, _14119_);
  nor (_18398_, _11247_, _18397_);
  and (_18399_, _11247_, _18397_);
  nor (_18400_, _18399_, _18398_);
  and (_18401_, _18400_, \oc8051_golden_model_1.PSW [7]);
  nor (_18402_, _18400_, \oc8051_golden_model_1.PSW [7]);
  nor (_18403_, _18402_, _18401_);
  and (_18404_, _18403_, _18395_);
  nor (_18405_, _18403_, _18395_);
  nor (_18406_, _18405_, _18404_);
  or (_18407_, _18406_, _10543_);
  nor (_18408_, _12529_, _10854_);
  or (_18409_, _18169_, _14092_);
  and (_18410_, _18409_, _14091_);
  nor (_18411_, _11209_, _18410_);
  and (_18412_, _11209_, _18410_);
  nor (_18413_, _18412_, _18411_);
  and (_18414_, _18413_, \oc8051_golden_model_1.PSW [7]);
  nor (_18415_, _18413_, \oc8051_golden_model_1.PSW [7]);
  nor (_18416_, _18415_, _18414_);
  and (_18417_, _18416_, _18408_);
  nor (_18418_, _18416_, _18408_);
  nor (_18419_, _18418_, _18417_);
  or (_18420_, _18419_, _06516_);
  not (_18421_, _18158_);
  nand (_18422_, _18161_, _18421_);
  and (_18423_, _09205_, _10218_);
  or (_18424_, _09205_, _10218_);
  and (_18425_, _18424_, _18153_);
  or (_18426_, _18425_, _18423_);
  nor (_18427_, _11170_, _18426_);
  and (_18428_, _11170_, _18426_);
  nor (_18429_, _18428_, _18427_);
  and (_18430_, _18429_, \oc8051_golden_model_1.PSW [7]);
  nor (_18431_, _18429_, \oc8051_golden_model_1.PSW [7]);
  nor (_18432_, _18431_, _18430_);
  and (_18433_, _18432_, _18422_);
  nor (_18434_, _18432_, _18422_);
  nor (_18435_, _18434_, _18433_);
  or (_18436_, _18435_, _10611_);
  nand (_18437_, _10682_, _08494_);
  and (_18438_, _15108_, _07914_);
  or (_18439_, _18438_, _18391_);
  and (_18440_, _18439_, _06251_);
  or (_18441_, _10688_, _09159_);
  nor (_18442_, _10704_, _08494_);
  nor (_18443_, _06808_, _10087_);
  and (_18444_, _06808_, _10087_);
  or (_18445_, _18444_, _18443_);
  and (_18446_, _18445_, _10704_);
  or (_18447_, _18446_, _10687_);
  or (_18448_, _18447_, _18442_);
  and (_18449_, _18448_, _10714_);
  and (_18450_, _18449_, _18441_);
  or (_18451_, _18450_, _18440_);
  and (_18452_, _18451_, _10719_);
  nor (_18453_, _10722_, \oc8051_golden_model_1.ACC [4]);
  nor (_18454_, _18453_, _10723_);
  and (_18455_, _18454_, _10718_);
  or (_18456_, _18455_, _06475_);
  or (_18457_, _18456_, _18452_);
  nor (_18458_, _08545_, _10087_);
  and (_18459_, _15091_, _08545_);
  or (_18460_, _18459_, _18458_);
  or (_18461_, _18460_, _06476_);
  and (_18462_, _18461_, _07142_);
  and (_18463_, _18462_, _18457_);
  and (_18464_, _18393_, _06468_);
  or (_18465_, _18464_, _10682_);
  or (_18466_, _18465_, _18463_);
  and (_18467_, _18466_, _18437_);
  or (_18468_, _18467_, _07153_);
  or (_18469_, _09159_, _07353_);
  and (_18470_, _18469_, _06801_);
  and (_18471_, _18470_, _18468_);
  nor (_18472_, _08496_, _06801_);
  or (_18473_, _18472_, _10759_);
  or (_18474_, _18473_, _18471_);
  nand (_18475_, _10759_, _05997_);
  and (_18476_, _18475_, _18474_);
  or (_18477_, _18476_, _06483_);
  and (_18478_, _15089_, _08545_);
  or (_18479_, _18478_, _18458_);
  or (_18480_, _18479_, _06484_);
  and (_18481_, _18480_, _07164_);
  and (_18482_, _18481_, _18477_);
  or (_18483_, _18458_, _15125_);
  and (_18484_, _18483_, _06461_);
  and (_18485_, _18484_, _18460_);
  or (_18486_, _18485_, _09487_);
  or (_18487_, _18486_, _18482_);
  nor (_18488_, _09985_, _09983_);
  nor (_18489_, _18488_, _09986_);
  or (_18490_, _18489_, _09494_);
  and (_18491_, _18490_, _10779_);
  and (_18492_, _18491_, _18487_);
  or (_18493_, _18146_, _18139_);
  nor (_18494_, _07713_, \oc8051_golden_model_1.ACC [3]);
  nand (_18495_, _07713_, \oc8051_golden_model_1.ACC [3]);
  and (_18496_, _18495_, _18134_);
  or (_18497_, _18496_, _18494_);
  nor (_18498_, _11126_, _18497_);
  and (_18499_, _11126_, _18497_);
  nor (_18500_, _18499_, _18498_);
  and (_18501_, _18500_, \oc8051_golden_model_1.PSW [7]);
  nor (_18502_, _18500_, \oc8051_golden_model_1.PSW [7]);
  nor (_18503_, _18502_, _18501_);
  or (_18504_, _18503_, _18493_);
  and (_18505_, _18503_, _18493_);
  nor (_18506_, _18505_, _10779_);
  and (_18507_, _18506_, _18504_);
  or (_18508_, _18507_, _10610_);
  or (_18509_, _18508_, _18492_);
  and (_18510_, _18509_, _18436_);
  or (_18511_, _18510_, _06510_);
  and (_18512_, _18511_, _18420_);
  or (_18513_, _18512_, _10542_);
  and (_18514_, _18513_, _18407_);
  or (_18515_, _18514_, _05976_);
  nand (_18516_, _06230_, _05976_);
  and (_18517_, _18516_, _06242_);
  and (_18518_, _18517_, _18515_);
  or (_18519_, _18458_, _15141_);
  and (_18520_, _18519_, _06241_);
  and (_18521_, _18520_, _18460_);
  or (_18522_, _18521_, _07187_);
  or (_18523_, _18522_, _18518_);
  and (_18524_, _18523_, _18394_);
  or (_18525_, _18524_, _07182_);
  and (_18526_, _09159_, _07914_);
  or (_18527_, _18391_, _07183_);
  or (_18528_, _18527_, _18526_);
  and (_18529_, _18528_, _06336_);
  and (_18530_, _18529_, _18525_);
  and (_18531_, _15198_, _07914_);
  or (_18532_, _18531_, _18391_);
  and (_18533_, _18532_, _05968_);
  or (_18534_, _18533_, _10046_);
  or (_18535_, _18534_, _18530_);
  or (_18536_, _10133_, _10052_);
  and (_18537_, _18536_, _18535_);
  or (_18538_, _18537_, _05935_);
  and (_18539_, _18538_, _18390_);
  or (_18540_, _18539_, _06371_);
  and (_18541_, _08892_, _07914_);
  or (_18542_, _18541_, _18391_);
  or (_18543_, _18542_, _07198_);
  and (_18544_, _18543_, _10905_);
  and (_18545_, _18544_, _18540_);
  nor (_18546_, _10905_, _06230_);
  or (_18547_, _18546_, _18226_);
  or (_18548_, _18547_, _18545_);
  not (_18549_, _06683_);
  or (_18550_, _11126_, _18549_);
  and (_18551_, _18550_, _18224_);
  and (_18552_, _18551_, _18548_);
  and (_18553_, _11126_, _18223_);
  or (_18554_, _18553_, _06698_);
  or (_18555_, _18554_, _18552_);
  and (_18556_, _18555_, _18389_);
  and (_18557_, _11126_, _06697_);
  nor (_18558_, _18557_, _18556_);
  or (_18559_, _18558_, _17188_);
  nand (_18560_, _11126_, _17188_);
  and (_18561_, _18560_, _18559_);
  nor (_18562_, _18561_, _18386_);
  and (_18563_, _11126_, _18386_);
  or (_18564_, _18563_, _18562_);
  and (_18565_, _18564_, _17748_);
  and (_18566_, _17747_, _11126_);
  or (_18567_, _18566_, _17915_);
  or (_18568_, _18567_, _18565_);
  or (_18569_, _11126_, _17919_);
  and (_18570_, _18569_, _10930_);
  and (_18571_, _18570_, _18568_);
  and (_18572_, _10929_, _11170_);
  or (_18573_, _18572_, _06531_);
  or (_18574_, _18573_, _18571_);
  and (_18575_, _18574_, _18385_);
  and (_18576_, _11247_, _10533_);
  or (_18577_, _18576_, _06367_);
  or (_18578_, _18577_, _18575_);
  and (_18579_, _15214_, _07914_);
  or (_18580_, _18579_, _18391_);
  or (_18581_, _18580_, _07218_);
  and (_18582_, _18581_, _18578_);
  or (_18583_, _18582_, _06533_);
  or (_18584_, _18391_, _07216_);
  and (_18585_, _18584_, _12225_);
  and (_18586_, _18585_, _18583_);
  and (_18587_, _17938_, _11123_);
  or (_18588_, _18587_, _10960_);
  or (_18589_, _18588_, _18586_);
  or (_18590_, _10962_, _11167_);
  and (_18591_, _18590_, _18589_);
  or (_18592_, _18591_, _06539_);
  or (_18593_, _11206_, _06540_);
  and (_18594_, _18593_, _10972_);
  and (_18595_, _18594_, _18592_);
  and (_18596_, _10966_, _11244_);
  or (_18597_, _18596_, _18595_);
  and (_18598_, _18597_, _07213_);
  nand (_18599_, _18542_, _06366_);
  nor (_18600_, _18599_, _11208_);
  or (_18601_, _18600_, _06654_);
  or (_18602_, _18601_, _18598_);
  and (_18603_, _18602_, _18383_);
  and (_18604_, _12221_, _06382_);
  or (_18605_, _18604_, _18603_);
  not (_18606_, _18604_);
  or (_18607_, _18606_, _11124_);
  and (_18608_, _18607_, _10993_);
  and (_18609_, _18608_, _18605_);
  and (_18610_, _11124_, _10992_);
  or (_18611_, _18610_, _10998_);
  or (_18612_, _18611_, _18609_);
  not (_18613_, _10998_);
  or (_18614_, _18613_, _11169_);
  and (_18615_, _18614_, _06527_);
  and (_18616_, _18615_, _18612_);
  nand (_18617_, _11007_, _11208_);
  and (_18618_, _18617_, _11006_);
  or (_18619_, _18618_, _18616_);
  and (_18620_, _18619_, _18381_);
  or (_18621_, _18620_, _06383_);
  and (_18622_, _15211_, _07914_);
  or (_18623_, _18391_, _07231_);
  or (_18624_, _18623_, _18622_);
  and (_18625_, _18624_, _10526_);
  and (_18626_, _18625_, _18621_);
  or (_18627_, _10512_, _10484_);
  and (_18628_, _18627_, _10513_);
  and (_18629_, _18628_, _11014_);
  or (_18630_, _18629_, _10452_);
  or (_18631_, _18630_, _18626_);
  or (_18632_, _11037_, _10638_);
  and (_18633_, _18632_, _11038_);
  or (_18634_, _18633_, _11022_);
  and (_18635_, _18634_, _06538_);
  and (_18636_, _18635_, _18631_);
  or (_18637_, _11067_, _10573_);
  and (_18638_, _18637_, _11068_);
  or (_18639_, _18638_, _11050_);
  and (_18640_, _18639_, _11052_);
  or (_18641_, _18640_, _18636_);
  or (_18642_, _11097_, _10836_);
  and (_18643_, _18642_, _11098_);
  or (_18644_, _18643_, _11082_);
  and (_18645_, _18644_, _18641_);
  or (_18646_, _18645_, _11080_);
  nand (_18647_, _11080_, _10218_);
  and (_18648_, _18647_, _12103_);
  and (_18649_, _18648_, _18646_);
  or (_18650_, _11142_, _11126_);
  nor (_18651_, _12103_, _11143_);
  and (_18652_, _18651_, _18650_);
  or (_18653_, _18652_, _17443_);
  or (_18654_, _18653_, _18649_);
  or (_18655_, _11186_, _11170_);
  and (_18656_, _18655_, _11187_);
  or (_18657_, _18656_, _17444_);
  and (_18658_, _18657_, _18654_);
  and (_18659_, _18658_, _17700_);
  and (_18660_, _18656_, _17442_);
  or (_18661_, _18660_, _18659_);
  or (_18662_, _18661_, _06293_);
  and (_18663_, _18662_, _18380_);
  or (_18664_, _11263_, _11247_);
  and (_18665_, _18664_, _11264_);
  and (_18666_, _18665_, _10450_);
  or (_18667_, _18666_, _10448_);
  or (_18668_, _18667_, _18663_);
  and (_18669_, _18668_, _18376_);
  or (_18670_, _18669_, _06563_);
  or (_18671_, _18439_, _07241_);
  and (_18672_, _18671_, _11280_);
  and (_18673_, _18672_, _18670_);
  nor (_18674_, _11286_, _10087_);
  or (_18675_, _18674_, _11287_);
  and (_18676_, _18675_, _11279_);
  or (_18677_, _18676_, _11284_);
  or (_18678_, _18677_, _18673_);
  nand (_18679_, _11284_, _10122_);
  and (_18680_, _18679_, _06571_);
  and (_18681_, _18680_, _18678_);
  and (_18682_, _18479_, _06199_);
  or (_18683_, _18682_, _06188_);
  or (_18684_, _18683_, _18681_);
  and (_18685_, _15280_, _07914_);
  or (_18686_, _18685_, _18391_);
  or (_18687_, _18686_, _06189_);
  and (_18688_, _18687_, _11303_);
  and (_18689_, _18688_, _18684_);
  nor (_18690_, _11312_, \oc8051_golden_model_1.ACC [4]);
  nor (_18691_, _18690_, _11313_);
  and (_18692_, _18691_, _11302_);
  or (_18693_, _18692_, _11309_);
  or (_18694_, _18693_, _18689_);
  nand (_18695_, _11309_, _10122_);
  and (_18696_, _18695_, _01452_);
  and (_18697_, _18696_, _18694_);
  or (_18698_, _18697_, _18375_);
  and (_43774_, _18698_, _43223_);
  nor (_18699_, _01452_, _10122_);
  and (_18700_, _10514_, _10478_);
  nor (_18701_, _18700_, _10515_);
  or (_18702_, _18701_, _10526_);
  and (_18703_, _10919_, _11122_);
  nor (_18704_, _10905_, _06608_);
  nand (_18705_, _06608_, _05935_);
  nor (_18706_, _07914_, _10122_);
  nor (_18707_, _08209_, _10538_);
  or (_18708_, _18707_, _18706_);
  or (_18709_, _18708_, _07188_);
  and (_18710_, _06230_, \oc8051_golden_model_1.ACC [4]);
  nor (_18711_, _18398_, _18710_);
  and (_18712_, _12551_, _18711_);
  nor (_18713_, _12551_, _18711_);
  nor (_18714_, _18713_, _18712_);
  and (_18715_, _18714_, \oc8051_golden_model_1.PSW [7]);
  nor (_18716_, _18714_, \oc8051_golden_model_1.PSW [7]);
  nor (_18717_, _18716_, _18715_);
  nor (_18718_, _18404_, _18401_);
  not (_18719_, _18718_);
  and (_18720_, _18719_, _18717_);
  nor (_18721_, _18719_, _18717_);
  nor (_18722_, _18721_, _18720_);
  or (_18723_, _18722_, _10543_);
  nor (_18724_, _09159_, _10087_);
  nor (_18725_, _18427_, _18724_);
  nor (_18726_, _11166_, _18725_);
  and (_18727_, _11166_, _18725_);
  nor (_18728_, _18727_, _18726_);
  nor (_18729_, _18728_, _10854_);
  and (_18730_, _18728_, _10854_);
  nor (_18731_, _18730_, _18729_);
  nor (_18732_, _18433_, _18430_);
  not (_18733_, _18732_);
  nor (_18734_, _18733_, _18731_);
  and (_18735_, _18733_, _18731_);
  or (_18736_, _18735_, _10611_);
  nor (_18737_, _18736_, _18734_);
  nor (_18738_, _08545_, _10122_);
  and (_18739_, _15296_, _08545_);
  or (_18740_, _18739_, _18738_);
  or (_18741_, _18738_, _15328_);
  and (_18742_, _18741_, _06461_);
  and (_18743_, _18742_, _18740_);
  nand (_18744_, _10682_, _08209_);
  or (_18745_, _10688_, _09113_);
  nor (_18746_, _10704_, _08209_);
  or (_18747_, _06808_, \oc8051_golden_model_1.ACC [5]);
  nand (_18748_, _06808_, \oc8051_golden_model_1.ACC [5]);
  and (_18749_, _18748_, _18747_);
  and (_18750_, _18749_, _10704_);
  or (_18751_, _18750_, _10687_);
  or (_18752_, _18751_, _18746_);
  and (_18753_, _18752_, _10714_);
  and (_18754_, _18753_, _18745_);
  and (_18755_, _15311_, _07914_);
  or (_18756_, _18755_, _18706_);
  and (_18757_, _18756_, _06251_);
  or (_18758_, _18757_, _10718_);
  or (_18759_, _18758_, _18754_);
  nor (_18760_, _10738_, _10730_);
  and (_18761_, _10738_, _10730_);
  or (_18762_, _18761_, _18760_);
  or (_18763_, _18762_, _10719_);
  and (_18764_, _18763_, _18759_);
  or (_18765_, _18764_, _06475_);
  or (_18766_, _18740_, _06476_);
  and (_18767_, _18766_, _07142_);
  and (_18768_, _18767_, _18765_);
  and (_18769_, _18708_, _06468_);
  or (_18770_, _18769_, _10682_);
  or (_18771_, _18770_, _18768_);
  and (_18772_, _18771_, _18744_);
  or (_18773_, _18772_, _07153_);
  or (_18774_, _09113_, _07353_);
  and (_18775_, _18774_, _06801_);
  and (_18776_, _18775_, _18773_);
  nor (_18777_, _08211_, _06801_);
  or (_18779_, _18777_, _10759_);
  or (_18780_, _18779_, _18776_);
  nand (_18781_, _10759_, _05937_);
  and (_18782_, _18781_, _18780_);
  or (_18783_, _18782_, _06483_);
  and (_18784_, _15294_, _08545_);
  or (_18785_, _18784_, _18738_);
  or (_18786_, _18785_, _06484_);
  and (_18787_, _18786_, _07164_);
  and (_18788_, _18787_, _18783_);
  or (_18790_, _18788_, _18743_);
  and (_18791_, _18790_, _09494_);
  or (_18792_, _09988_, _09986_);
  nor (_18793_, _09989_, _09494_);
  and (_18794_, _18793_, _18792_);
  or (_18795_, _18794_, _12236_);
  or (_18796_, _18795_, _18791_);
  and (_18797_, _08494_, \oc8051_golden_model_1.ACC [4]);
  nor (_18798_, _18498_, _18797_);
  nor (_18799_, _11122_, _18798_);
  and (_18801_, _11122_, _18798_);
  nor (_18802_, _18801_, _18799_);
  and (_18803_, _18802_, \oc8051_golden_model_1.PSW [7]);
  nor (_18804_, _18802_, \oc8051_golden_model_1.PSW [7]);
  nor (_18805_, _18804_, _18803_);
  nor (_18806_, _18505_, _18501_);
  not (_18807_, _18806_);
  and (_18808_, _18807_, _18805_);
  nor (_18809_, _18807_, _18805_);
  nor (_18810_, _18809_, _18808_);
  or (_18812_, _18810_, _10779_);
  and (_18813_, _18812_, _10611_);
  and (_18814_, _18813_, _18796_);
  or (_18815_, _18814_, _18737_);
  and (_18816_, _18815_, _06516_);
  nor (_18817_, _18417_, _18414_);
  and (_18818_, _08496_, \oc8051_golden_model_1.ACC [4]);
  nor (_18819_, _18411_, _18818_);
  nor (_18820_, _11205_, _18819_);
  and (_18821_, _11205_, _18819_);
  nor (_18823_, _18821_, _18820_);
  and (_18824_, _18823_, \oc8051_golden_model_1.PSW [7]);
  nor (_18825_, _18823_, \oc8051_golden_model_1.PSW [7]);
  or (_18826_, _18825_, _18824_);
  nor (_18827_, _18826_, _18817_);
  and (_18828_, _18826_, _18817_);
  nor (_18829_, _18828_, _18827_);
  or (_18830_, _18829_, _10542_);
  and (_18831_, _18830_, _12589_);
  or (_18832_, _18831_, _18816_);
  and (_18834_, _18832_, _18723_);
  or (_18835_, _18834_, _05976_);
  nand (_18836_, _06608_, _05976_);
  and (_18837_, _18836_, _06242_);
  and (_18838_, _18837_, _18835_);
  or (_18839_, _18738_, _15344_);
  and (_18840_, _18839_, _06241_);
  and (_18841_, _18840_, _18740_);
  or (_18842_, _18841_, _07187_);
  or (_18843_, _18842_, _18838_);
  and (_18845_, _18843_, _18709_);
  or (_18846_, _18845_, _07182_);
  and (_18847_, _09113_, _07914_);
  or (_18848_, _18706_, _07183_);
  or (_18849_, _18848_, _18847_);
  and (_18850_, _18849_, _06336_);
  and (_18851_, _18850_, _18846_);
  and (_18852_, _15400_, _07914_);
  or (_18853_, _18852_, _18706_);
  and (_18854_, _18853_, _05968_);
  or (_18856_, _18854_, _10046_);
  or (_18857_, _18856_, _18851_);
  or (_18858_, _10105_, _10052_);
  and (_18859_, _18858_, _18857_);
  or (_18860_, _18859_, _05935_);
  and (_18861_, _18860_, _18705_);
  or (_18862_, _18861_, _06371_);
  and (_18863_, _08888_, _07914_);
  or (_18864_, _18863_, _18706_);
  or (_18865_, _18864_, _07198_);
  and (_18867_, _18865_, _10905_);
  and (_18868_, _18867_, _18862_);
  or (_18869_, _18868_, _18704_);
  and (_18870_, _18869_, _18549_);
  and (_18871_, _11122_, _06683_);
  or (_18872_, _18871_, _06698_);
  or (_18873_, _18872_, _18870_);
  or (_18874_, _11122_, _18387_);
  and (_18875_, _18874_, _10920_);
  and (_18876_, _18875_, _18873_);
  or (_18878_, _18876_, _18703_);
  and (_18879_, _18878_, _17748_);
  and (_18880_, _17747_, _11122_);
  or (_18881_, _18880_, _17915_);
  or (_18882_, _18881_, _18879_);
  or (_18883_, _11122_, _17919_);
  and (_18884_, _18883_, _10930_);
  and (_18885_, _18884_, _18882_);
  nor (_18886_, _10930_, _11166_);
  or (_18887_, _18886_, _06531_);
  or (_18889_, _18887_, _18885_);
  or (_18890_, _11205_, _06532_);
  and (_18891_, _18890_, _10534_);
  and (_18892_, _18891_, _18889_);
  nor (_18893_, _12550_, _10534_);
  or (_18894_, _18893_, _06367_);
  or (_18895_, _18894_, _18892_);
  and (_18896_, _15416_, _07914_);
  or (_18897_, _18896_, _18706_);
  or (_18898_, _18897_, _07218_);
  and (_18900_, _18898_, _18895_);
  or (_18901_, _18900_, _06533_);
  or (_18902_, _18706_, _07216_);
  and (_18903_, _18902_, _12225_);
  and (_18904_, _18903_, _18901_);
  and (_18905_, _17938_, _11120_);
  or (_18906_, _18905_, _10960_);
  or (_18907_, _18906_, _18904_);
  or (_18908_, _10962_, _11164_);
  and (_18909_, _18908_, _06540_);
  and (_18911_, _18909_, _18907_);
  or (_18912_, _10966_, _11203_);
  and (_18913_, _18912_, _10968_);
  or (_18914_, _18913_, _18911_);
  or (_18915_, _10972_, _11243_);
  and (_18916_, _18915_, _07213_);
  and (_18917_, _18916_, _18914_);
  nand (_18918_, _18864_, _06366_);
  nor (_18919_, _18918_, _11204_);
  or (_18920_, _18919_, _18917_);
  and (_18922_, _18920_, _17637_);
  nor (_18923_, _17637_, _11121_);
  or (_18924_, _18923_, _10988_);
  or (_18925_, _18924_, _18922_);
  nand (_18926_, _10988_, _11121_);
  and (_18927_, _18926_, _10993_);
  and (_18928_, _18927_, _18925_);
  nor (_18929_, _11121_, _10993_);
  or (_18930_, _18929_, _10998_);
  or (_18931_, _18930_, _18928_);
  nand (_18933_, _10998_, _10122_);
  or (_18934_, _18933_, _09113_);
  and (_18935_, _18934_, _18931_);
  or (_18936_, _18935_, _06526_);
  nand (_18937_, _11204_, _06526_);
  and (_18938_, _18937_, _11007_);
  and (_18939_, _18938_, _18936_);
  and (_18940_, _11004_, _11242_);
  or (_18941_, _18940_, _18939_);
  and (_18942_, _18941_, _07231_);
  and (_18944_, _15413_, _07914_);
  or (_18945_, _18944_, _18706_);
  and (_18946_, _18945_, _06383_);
  or (_18947_, _18946_, _11014_);
  or (_18948_, _18947_, _18942_);
  and (_18949_, _18948_, _18702_);
  or (_18950_, _18949_, _10452_);
  and (_18951_, _11039_, _10635_);
  nor (_18952_, _18951_, _11040_);
  or (_18953_, _18952_, _11022_);
  and (_18954_, _18953_, _06538_);
  and (_18955_, _18954_, _18950_);
  nand (_18956_, _11069_, _10570_);
  nor (_18957_, _11070_, _06538_);
  and (_18958_, _18957_, _18956_);
  or (_18959_, _18958_, _11050_);
  or (_18960_, _18959_, _18955_);
  and (_18961_, _11099_, _10833_);
  nor (_18962_, _18961_, _11100_);
  or (_18963_, _18962_, _11082_);
  and (_18965_, _18963_, _11081_);
  and (_18966_, _18965_, _18960_);
  and (_18967_, _11080_, \oc8051_golden_model_1.ACC [4]);
  or (_18968_, _18967_, _11111_);
  or (_18969_, _18968_, _18966_);
  nor (_18970_, _11145_, _11122_);
  nor (_18971_, _18970_, _11146_);
  or (_18972_, _18971_, _11116_);
  and (_18973_, _18972_, _11115_);
  and (_18974_, _18973_, _18969_);
  and (_18976_, _18971_, _11114_);
  or (_18977_, _18976_, _11156_);
  or (_18978_, _18977_, _18974_);
  and (_18979_, _11188_, _11166_);
  nor (_18980_, _18979_, _11189_);
  or (_18981_, _18980_, _11160_);
  and (_18982_, _18981_, _06295_);
  and (_18983_, _18982_, _18978_);
  nor (_18984_, _11228_, _11205_);
  nor (_18985_, _18984_, _11229_);
  and (_18987_, _18985_, _06293_);
  or (_18988_, _18987_, _10450_);
  or (_18989_, _18988_, _18983_);
  and (_18990_, _11265_, _12551_);
  nor (_18991_, _11265_, _12551_);
  or (_18992_, _18991_, _10451_);
  or (_18993_, _18992_, _18990_);
  and (_18994_, _18993_, _12966_);
  and (_18995_, _18994_, _18989_);
  and (_18996_, _10448_, \oc8051_golden_model_1.ACC [4]);
  or (_18998_, _18996_, _06563_);
  or (_18999_, _18998_, _18995_);
  or (_19000_, _18756_, _07241_);
  and (_19001_, _19000_, _11280_);
  and (_19002_, _19001_, _18999_);
  nor (_19003_, _11287_, _10122_);
  or (_19004_, _19003_, _11288_);
  nor (_19005_, _19004_, _11284_);
  nor (_19006_, _19005_, _12991_);
  or (_19007_, _19006_, _19002_);
  nand (_19009_, _11284_, _10068_);
  and (_19010_, _19009_, _06571_);
  and (_19011_, _19010_, _19007_);
  and (_19012_, _18785_, _06199_);
  or (_19013_, _19012_, _06188_);
  or (_19014_, _19013_, _19011_);
  and (_19015_, _15477_, _07914_);
  or (_19016_, _19015_, _18706_);
  or (_19017_, _19016_, _06189_);
  and (_19018_, _19017_, _11303_);
  and (_19020_, _19018_, _19014_);
  nor (_19021_, _11313_, \oc8051_golden_model_1.ACC [5]);
  nor (_19022_, _19021_, _11314_);
  nor (_19023_, _19022_, _11309_);
  nor (_19024_, _19023_, _13013_);
  or (_19025_, _19024_, _19020_);
  nand (_19026_, _11309_, _10068_);
  and (_19027_, _19026_, _01452_);
  and (_19028_, _19027_, _19025_);
  or (_19029_, _19028_, _18699_);
  and (_43775_, _19029_, _43223_);
  nor (_19031_, _01452_, _10068_);
  nand (_19032_, _10448_, _10122_);
  nor (_19033_, _11071_, _10603_);
  nor (_19034_, _19033_, _11072_);
  or (_19035_, _19034_, _06538_);
  and (_19036_, _19035_, _11082_);
  and (_19037_, _10998_, _11162_);
  not (_19038_, _18386_);
  or (_19039_, _11119_, _19038_);
  nor (_19041_, _07914_, _10068_);
  and (_19042_, _15601_, _07914_);
  or (_19043_, _19042_, _19041_);
  and (_19044_, _19043_, _05968_);
  nor (_19045_, _08106_, _10538_);
  or (_19046_, _19045_, _19041_);
  or (_19047_, _19046_, _07188_);
  or (_19048_, _09113_, _10122_);
  and (_19049_, _09113_, _10122_);
  or (_19050_, _18725_, _19049_);
  and (_19052_, _19050_, _19048_);
  nor (_19053_, _19052_, _11163_);
  and (_19054_, _19052_, _11163_);
  nor (_19055_, _19054_, _19053_);
  nor (_19056_, _18735_, _18729_);
  and (_19057_, _19056_, \oc8051_golden_model_1.PSW [7]);
  or (_19058_, _19057_, _19055_);
  nand (_19059_, _19057_, _19055_);
  and (_19060_, _19059_, _19058_);
  or (_19061_, _19060_, _10611_);
  nand (_19063_, _10682_, _08106_);
  not (_19064_, _10732_);
  nor (_19065_, _18760_, _19064_);
  or (_19066_, _10738_, _10734_);
  nand (_19067_, _19066_, _10718_);
  or (_19068_, _19067_, _19065_);
  or (_19069_, _10688_, _09067_);
  nor (_19070_, _10704_, _08106_);
  or (_19071_, _06808_, \oc8051_golden_model_1.ACC [6]);
  nand (_19072_, _06808_, \oc8051_golden_model_1.ACC [6]);
  and (_19074_, _19072_, _19071_);
  and (_19075_, _19074_, _10704_);
  or (_19076_, _19075_, _10687_);
  or (_19077_, _19076_, _19070_);
  and (_19078_, _19077_, _10714_);
  and (_19079_, _19078_, _19069_);
  and (_19080_, _15512_, _07914_);
  or (_19081_, _19080_, _19041_);
  and (_19082_, _19081_, _06251_);
  or (_19083_, _19082_, _10718_);
  or (_19085_, _19083_, _19079_);
  and (_19086_, _19085_, _19068_);
  or (_19087_, _19086_, _06475_);
  nor (_19088_, _08545_, _10068_);
  and (_19089_, _15499_, _08545_);
  or (_19090_, _19089_, _19088_);
  or (_19091_, _19090_, _06476_);
  and (_19092_, _19091_, _07142_);
  and (_19093_, _19092_, _19087_);
  and (_19094_, _19046_, _06468_);
  or (_19096_, _19094_, _10682_);
  or (_19097_, _19096_, _19093_);
  and (_19098_, _19097_, _19063_);
  or (_19099_, _19098_, _07153_);
  or (_19100_, _09067_, _07353_);
  and (_19101_, _19100_, _06801_);
  and (_19102_, _19101_, _19099_);
  nor (_19103_, _08108_, _06801_);
  or (_19104_, _19103_, _10759_);
  or (_19105_, _19104_, _19102_);
  nand (_19107_, _10759_, _10165_);
  and (_19108_, _19107_, _19105_);
  or (_19109_, _19108_, _06483_);
  and (_19110_, _15497_, _08545_);
  or (_19111_, _19110_, _19088_);
  or (_19112_, _19111_, _06484_);
  and (_19113_, _19112_, _07164_);
  and (_19114_, _19113_, _19109_);
  or (_19115_, _19088_, _15529_);
  and (_19116_, _19115_, _06461_);
  and (_19118_, _19116_, _19090_);
  or (_19119_, _19118_, _09487_);
  or (_19120_, _19119_, _19114_);
  nor (_19121_, _09991_, _09989_);
  nor (_19122_, _19121_, _09992_);
  or (_19123_, _19122_, _09494_);
  and (_19124_, _19123_, _10779_);
  and (_19125_, _19124_, _19120_);
  nand (_19126_, _08209_, \oc8051_golden_model_1.ACC [5]);
  nor (_19127_, _08209_, \oc8051_golden_model_1.ACC [5]);
  or (_19129_, _18798_, _19127_);
  and (_19130_, _19129_, _19126_);
  nor (_19131_, _19130_, _11119_);
  and (_19132_, _19130_, _11119_);
  nor (_19133_, _19132_, _19131_);
  nor (_19134_, _18808_, _18803_);
  and (_19135_, _19134_, \oc8051_golden_model_1.PSW [7]);
  or (_19136_, _19135_, _19133_);
  nand (_19137_, _19135_, _19133_);
  and (_19138_, _19137_, _19136_);
  and (_19140_, _19138_, _12236_);
  or (_19141_, _19140_, _10610_);
  or (_19142_, _19141_, _19125_);
  and (_19143_, _19142_, _12588_);
  and (_19144_, _19143_, _19061_);
  or (_19145_, _18711_, _12548_);
  and (_19146_, _19145_, _14112_);
  nor (_19147_, _19146_, _11241_);
  and (_19148_, _19146_, _11241_);
  nor (_19149_, _19148_, _19147_);
  nor (_19151_, _18720_, _18715_);
  and (_19152_, _19151_, \oc8051_golden_model_1.PSW [7]);
  or (_19153_, _19152_, _19149_);
  nand (_19154_, _19152_, _19149_);
  and (_19155_, _19154_, _10542_);
  and (_19156_, _19155_, _19153_);
  or (_19157_, _19156_, _05976_);
  or (_19158_, _18819_, _14081_);
  and (_19159_, _19158_, _14080_);
  nor (_19160_, _19159_, _11202_);
  and (_19162_, _19159_, _11202_);
  nor (_19163_, _19162_, _19160_);
  nor (_19164_, _18823_, _10854_);
  and (_19165_, _18817_, _19164_);
  nand (_19166_, _19165_, _19163_);
  or (_19167_, _19165_, _19163_);
  and (_19168_, _19167_, _06510_);
  and (_19169_, _19168_, _19166_);
  or (_19170_, _19169_, _19157_);
  or (_19171_, _19170_, _19144_);
  nand (_19173_, _06326_, _05976_);
  and (_19174_, _19173_, _06242_);
  and (_19175_, _19174_, _19171_);
  or (_19176_, _19088_, _15545_);
  and (_19177_, _19176_, _06241_);
  and (_19178_, _19177_, _19090_);
  or (_19179_, _19178_, _07187_);
  or (_19180_, _19179_, _19175_);
  and (_19181_, _19180_, _19047_);
  or (_19182_, _19181_, _07182_);
  and (_19184_, _09067_, _07914_);
  or (_19185_, _19041_, _07183_);
  or (_19186_, _19185_, _19184_);
  and (_19187_, _19186_, _06336_);
  and (_19188_, _19187_, _19182_);
  or (_19189_, _19188_, _19044_);
  and (_19190_, _19189_, _12611_);
  nor (_19191_, _06326_, _05975_);
  not (_19192_, _10074_);
  or (_19193_, _19192_, _10069_);
  nor (_19195_, _19193_, _05934_);
  and (_19196_, _19195_, _10046_);
  or (_19197_, _19196_, _19191_);
  or (_19198_, _19197_, _19190_);
  and (_19199_, _19198_, _07198_);
  and (_19200_, _15608_, _07914_);
  or (_19201_, _19200_, _19041_);
  and (_19202_, _19201_, _06371_);
  or (_19203_, _19202_, _10904_);
  or (_19204_, _19203_, _19199_);
  nand (_19206_, _10904_, _06326_);
  and (_19207_, _19206_, _18549_);
  and (_19208_, _19207_, _19204_);
  and (_19209_, _11119_, _06683_);
  or (_19210_, _19209_, _06698_);
  or (_19211_, _19210_, _19208_);
  or (_19212_, _11119_, _18387_);
  and (_19213_, _19212_, _17189_);
  and (_19214_, _19213_, _19211_);
  and (_19215_, _17190_, _11119_);
  or (_19217_, _19215_, _18386_);
  or (_19218_, _19217_, _19214_);
  and (_19219_, _19218_, _19039_);
  or (_19220_, _19219_, _17747_);
  or (_19221_, _17748_, _11119_);
  and (_19222_, _19221_, _17919_);
  and (_19223_, _19222_, _19220_);
  nand (_19224_, _11119_, _17915_);
  nand (_19225_, _19224_, _10930_);
  or (_19226_, _19225_, _19223_);
  or (_19228_, _10930_, _11163_);
  and (_19229_, _19228_, _19226_);
  or (_19230_, _19229_, _06531_);
  or (_19231_, _11202_, _06532_);
  and (_19232_, _19231_, _10534_);
  and (_19233_, _19232_, _19230_);
  and (_19234_, _11241_, _10533_);
  or (_19235_, _19234_, _06367_);
  or (_19236_, _19235_, _19233_);
  and (_19237_, _15618_, _07914_);
  or (_19239_, _19237_, _19041_);
  or (_19240_, _19239_, _07218_);
  and (_19241_, _19240_, _19236_);
  or (_19242_, _19241_, _06533_);
  or (_19243_, _19041_, _07216_);
  and (_19244_, _19243_, _12225_);
  and (_19245_, _19244_, _19242_);
  and (_19246_, _17938_, _11117_);
  or (_19247_, _19246_, _10960_);
  or (_19248_, _19247_, _19245_);
  or (_19250_, _10962_, _11161_);
  and (_19251_, _19250_, _06540_);
  and (_19252_, _19251_, _19248_);
  and (_19253_, _11199_, _06539_);
  or (_19254_, _19253_, _10966_);
  or (_19255_, _19254_, _19252_);
  or (_19256_, _10972_, _11239_);
  and (_19257_, _19256_, _07213_);
  and (_19258_, _19257_, _19255_);
  nand (_19259_, _19201_, _06366_);
  nor (_19261_, _19259_, _11201_);
  or (_19262_, _19261_, _19258_);
  and (_19263_, _19262_, _17637_);
  nor (_19264_, _17637_, _11118_);
  or (_19265_, _19264_, _10988_);
  or (_19266_, _19265_, _19263_);
  nand (_19267_, _10988_, _11118_);
  and (_19268_, _19267_, _10993_);
  nand (_19269_, _19268_, _19266_);
  or (_19270_, _11118_, _10993_);
  and (_19272_, _19270_, _18613_);
  and (_19273_, _19272_, _19269_);
  or (_19274_, _19273_, _19037_);
  and (_19275_, _19274_, _06527_);
  and (_19276_, _11201_, _06526_);
  or (_19277_, _19276_, _11004_);
  or (_19278_, _19277_, _19275_);
  or (_19279_, _11007_, _11240_);
  and (_19280_, _19279_, _07231_);
  and (_19281_, _19280_, _19278_);
  and (_19283_, _15615_, _07914_);
  or (_19284_, _19041_, _07231_);
  or (_19285_, _19284_, _19283_);
  nand (_19286_, _19285_, _10526_);
  or (_19287_, _19286_, _19281_);
  nor (_19288_, _10516_, _10472_);
  or (_19289_, _19288_, _10517_);
  or (_19290_, _19289_, _10526_);
  and (_19291_, _19290_, _17669_);
  and (_19292_, _19291_, _19287_);
  or (_19294_, _11041_, _10674_);
  and (_19295_, _19294_, _11042_);
  nand (_19296_, _19295_, _05932_);
  and (_19297_, _19296_, _10452_);
  nor (_19298_, _19297_, _19292_);
  nand (_19299_, _19295_, _17673_);
  nand (_19300_, _19299_, _06538_);
  or (_19301_, _19300_, _19298_);
  and (_19302_, _19301_, _19036_);
  or (_19303_, _11101_, _10869_);
  and (_19305_, _11102_, _11050_);
  and (_19306_, _19305_, _19303_);
  or (_19307_, _19306_, _11080_);
  or (_19308_, _19307_, _19302_);
  nand (_19309_, _11080_, _10122_);
  and (_19310_, _19309_, _12103_);
  and (_19311_, _19310_, _19308_);
  nor (_19312_, _11147_, _11119_);
  nor (_19313_, _19312_, _11148_);
  and (_19314_, _19313_, _12104_);
  or (_19316_, _19314_, _17443_);
  or (_19317_, _19316_, _19311_);
  nor (_19318_, _11190_, _11163_);
  nor (_19319_, _19318_, _11191_);
  or (_19320_, _19319_, _17444_);
  and (_19321_, _19320_, _19317_);
  or (_19322_, _19321_, _17442_);
  or (_19323_, _19319_, _17700_);
  and (_19324_, _19323_, _06295_);
  and (_19325_, _19324_, _19322_);
  or (_19327_, _11230_, _11202_);
  and (_19328_, _11231_, _06293_);
  and (_19329_, _19328_, _19327_);
  or (_19330_, _19329_, _19325_);
  and (_19331_, _19330_, _10451_);
  or (_19332_, _11268_, _11241_);
  nor (_19333_, _11269_, _10451_);
  and (_19334_, _19333_, _19332_);
  or (_19335_, _19334_, _10448_);
  or (_19336_, _19335_, _19331_);
  and (_19338_, _19336_, _19032_);
  or (_19339_, _19338_, _06563_);
  or (_19340_, _19081_, _07241_);
  and (_19341_, _19340_, _11280_);
  and (_19342_, _19341_, _19339_);
  nor (_19343_, _11288_, _10068_);
  or (_19344_, _19343_, _11289_);
  and (_19345_, _19344_, _11279_);
  or (_19346_, _19345_, _11284_);
  or (_19347_, _19346_, _19342_);
  nand (_19349_, _11284_, _08506_);
  and (_19350_, _19349_, _06571_);
  and (_19351_, _19350_, _19347_);
  and (_19352_, _19111_, _06199_);
  or (_19353_, _19352_, _06188_);
  or (_19354_, _19353_, _19351_);
  and (_19355_, _15676_, _07914_);
  or (_19356_, _19355_, _19041_);
  or (_19357_, _19356_, _06189_);
  and (_19358_, _19357_, _11303_);
  and (_19360_, _19358_, _19354_);
  nor (_19361_, _11314_, \oc8051_golden_model_1.ACC [6]);
  nor (_19362_, _19361_, _11315_);
  and (_19363_, _19362_, _11302_);
  or (_19364_, _19363_, _11309_);
  or (_19365_, _19364_, _19360_);
  nand (_19366_, _11309_, _08506_);
  and (_19367_, _19366_, _01452_);
  and (_19368_, _19367_, _19365_);
  or (_19369_, _19368_, _19031_);
  and (_43776_, _19369_, _43223_);
  not (_19371_, \oc8051_golden_model_1.PCON [0]);
  nor (_19372_, _01452_, _19371_);
  nand (_19373_, _11218_, _07923_);
  nor (_19374_, _07923_, _19371_);
  nor (_19375_, _19374_, _07210_);
  nand (_19376_, _19375_, _19373_);
  nor (_19377_, _08351_, _11326_);
  or (_19378_, _19377_, _19374_);
  or (_19379_, _19378_, _06252_);
  and (_19381_, _07923_, \oc8051_golden_model_1.ACC [0]);
  or (_19382_, _19381_, _19374_);
  and (_19383_, _19382_, _07123_);
  nor (_19384_, _07123_, _19371_);
  or (_19385_, _19384_, _06251_);
  or (_19386_, _19385_, _19383_);
  and (_19387_, _19386_, _07142_);
  and (_19388_, _19387_, _19379_);
  and (_19389_, _07923_, _07325_);
  or (_19390_, _19389_, _19374_);
  and (_19392_, _19390_, _06468_);
  or (_19393_, _19392_, _19388_);
  and (_19394_, _19393_, _06801_);
  and (_19395_, _19382_, _06466_);
  or (_19396_, _19395_, _07187_);
  or (_19397_, _19396_, _19394_);
  or (_19398_, _19390_, _07188_);
  and (_19399_, _19398_, _19397_);
  or (_19400_, _19399_, _07182_);
  and (_19401_, _09342_, _07923_);
  or (_19403_, _19374_, _07183_);
  or (_19404_, _19403_, _19401_);
  and (_19405_, _19404_, _19400_);
  or (_19406_, _19405_, _05968_);
  and (_19407_, _14427_, _07923_);
  or (_19408_, _19374_, _06336_);
  or (_19409_, _19408_, _19407_);
  and (_19410_, _19409_, _07198_);
  and (_19411_, _19410_, _19406_);
  and (_19412_, _07923_, _08908_);
  or (_19414_, _19412_, _19374_);
  and (_19415_, _19414_, _06371_);
  or (_19416_, _19415_, _06367_);
  or (_19417_, _19416_, _19411_);
  and (_19418_, _14442_, _07923_);
  or (_19419_, _19418_, _19374_);
  or (_19420_, _19419_, _07218_);
  and (_19421_, _19420_, _07216_);
  and (_19422_, _19421_, _19417_);
  nor (_19423_, _12526_, _11326_);
  or (_19425_, _19423_, _19374_);
  and (_19426_, _19373_, _06533_);
  and (_19427_, _19426_, _19425_);
  or (_19428_, _19427_, _19422_);
  and (_19429_, _19428_, _07213_);
  nand (_19430_, _19414_, _06366_);
  nor (_19431_, _19430_, _19377_);
  or (_19432_, _19431_, _06541_);
  or (_19433_, _19432_, _19429_);
  and (_19434_, _19433_, _19376_);
  or (_19436_, _19434_, _06383_);
  and (_19437_, _14325_, _07923_);
  or (_19438_, _19437_, _19374_);
  or (_19439_, _19438_, _07231_);
  and (_19440_, _19439_, _07229_);
  and (_19441_, _19440_, _19436_);
  not (_19442_, _06756_);
  and (_19443_, _19425_, _06528_);
  or (_19444_, _19443_, _19442_);
  or (_19445_, _19444_, _19441_);
  or (_19447_, _19378_, _06756_);
  and (_19448_, _19447_, _01452_);
  and (_19449_, _19448_, _19445_);
  or (_19450_, _19449_, _19372_);
  and (_43778_, _19450_, _43223_);
  not (_19451_, \oc8051_golden_model_1.PCON [1]);
  nor (_19452_, _01452_, _19451_);
  nand (_19453_, _07923_, _07018_);
  or (_19454_, _07923_, \oc8051_golden_model_1.PCON [1]);
  and (_19455_, _19454_, _06371_);
  and (_19457_, _19455_, _19453_);
  and (_19458_, _09297_, _07923_);
  nor (_19459_, _07923_, _19451_);
  or (_19460_, _19459_, _07183_);
  or (_19461_, _19460_, _19458_);
  nor (_19462_, _11326_, _07120_);
  nor (_19463_, _07187_, _06468_);
  or (_19464_, _19463_, _19459_);
  or (_19465_, _19464_, _19462_);
  and (_19466_, _07923_, \oc8051_golden_model_1.ACC [1]);
  or (_19468_, _19466_, _19459_);
  and (_19469_, _19468_, _06466_);
  or (_19470_, _19469_, _07187_);
  and (_19471_, _14503_, _07923_);
  not (_19472_, _19471_);
  and (_19473_, _19472_, _19454_);
  and (_19474_, _19473_, _06251_);
  nor (_19475_, _07123_, _19451_);
  and (_19476_, _19468_, _07123_);
  or (_19477_, _19476_, _19475_);
  and (_19479_, _19477_, _06252_);
  or (_19480_, _19479_, _06468_);
  or (_19481_, _19480_, _19474_);
  and (_19482_, _19481_, _06801_);
  or (_19483_, _19482_, _19470_);
  and (_19484_, _19483_, _19465_);
  or (_19485_, _19484_, _07182_);
  and (_19486_, _19485_, _06336_);
  and (_19487_, _19486_, _19461_);
  or (_19488_, _14609_, _11326_);
  and (_19490_, _19454_, _05968_);
  and (_19491_, _19490_, _19488_);
  or (_19492_, _19491_, _19487_);
  and (_19493_, _19492_, _07198_);
  or (_19494_, _19493_, _19457_);
  and (_19495_, _19494_, _07218_);
  or (_19496_, _14625_, _11326_);
  and (_19497_, _19454_, _06367_);
  and (_19498_, _19497_, _19496_);
  or (_19499_, _19498_, _06533_);
  or (_19501_, _19499_, _19495_);
  nor (_19502_, _11216_, _11326_);
  or (_19503_, _19502_, _19459_);
  nand (_19504_, _11215_, _07923_);
  and (_19505_, _19504_, _19503_);
  or (_19506_, _19505_, _07216_);
  and (_19507_, _19506_, _07213_);
  and (_19508_, _19507_, _19501_);
  or (_19509_, _14623_, _11326_);
  and (_19510_, _19454_, _06366_);
  and (_19512_, _19510_, _19509_);
  or (_19513_, _19512_, _06541_);
  or (_19514_, _19513_, _19508_);
  nor (_19515_, _19459_, _07210_);
  nand (_19516_, _19515_, _19504_);
  and (_19517_, _19516_, _07231_);
  and (_19518_, _19517_, _19514_);
  or (_19519_, _19453_, _08302_);
  and (_19520_, _19454_, _06383_);
  and (_19521_, _19520_, _19519_);
  or (_19523_, _19521_, _06528_);
  or (_19524_, _19523_, _19518_);
  or (_19525_, _19503_, _07229_);
  and (_19526_, _19525_, _07241_);
  and (_19527_, _19526_, _19524_);
  and (_19528_, _19473_, _06563_);
  or (_19529_, _19528_, _06188_);
  or (_19530_, _19529_, _19527_);
  or (_19531_, _19459_, _06189_);
  or (_19532_, _19531_, _19471_);
  and (_19534_, _19532_, _01452_);
  and (_19535_, _19534_, _19530_);
  or (_19536_, _19535_, _19452_);
  and (_43779_, _19536_, _43223_);
  not (_19537_, \oc8051_golden_model_1.PCON [2]);
  nor (_19538_, _01452_, _19537_);
  nor (_19539_, _07923_, _19537_);
  and (_19540_, _09251_, _07923_);
  or (_19541_, _19540_, _19539_);
  and (_19542_, _19541_, _07182_);
  and (_19544_, _14712_, _07923_);
  or (_19545_, _19544_, _19539_);
  or (_19546_, _19545_, _06252_);
  and (_19547_, _07923_, \oc8051_golden_model_1.ACC [2]);
  or (_19548_, _19547_, _19539_);
  and (_19549_, _19548_, _07123_);
  nor (_19550_, _07123_, _19537_);
  or (_19551_, _19550_, _06251_);
  or (_19552_, _19551_, _19549_);
  and (_19553_, _19552_, _07142_);
  and (_19555_, _19553_, _19546_);
  nor (_19556_, _11326_, _07578_);
  or (_19557_, _19556_, _19539_);
  and (_19558_, _19557_, _06468_);
  or (_19559_, _19558_, _19555_);
  and (_19560_, _19559_, _06801_);
  and (_19561_, _19548_, _06466_);
  or (_19562_, _19561_, _07187_);
  or (_19563_, _19562_, _19560_);
  or (_19564_, _19557_, _07188_);
  and (_19566_, _19564_, _07183_);
  and (_19567_, _19566_, _19563_);
  or (_19568_, _19567_, _05968_);
  or (_19569_, _19568_, _19542_);
  and (_19570_, _14808_, _07923_);
  or (_19571_, _19539_, _06336_);
  or (_19572_, _19571_, _19570_);
  and (_19573_, _19572_, _07198_);
  and (_19574_, _19573_, _19569_);
  and (_19575_, _07923_, _08945_);
  or (_19577_, _19575_, _19539_);
  and (_19578_, _19577_, _06371_);
  or (_19579_, _19578_, _06367_);
  or (_19580_, _19579_, _19574_);
  and (_19581_, _14824_, _07923_);
  or (_19582_, _19581_, _19539_);
  or (_19583_, _19582_, _07218_);
  and (_19584_, _19583_, _07216_);
  and (_19585_, _19584_, _19580_);
  and (_19586_, _11214_, _07923_);
  or (_19588_, _19586_, _19539_);
  and (_19589_, _19588_, _06533_);
  or (_19590_, _19589_, _19585_);
  and (_19591_, _19590_, _07213_);
  or (_19592_, _19539_, _08397_);
  and (_19593_, _19577_, _06366_);
  and (_19594_, _19593_, _19592_);
  or (_19595_, _19594_, _19591_);
  and (_19596_, _19595_, _07210_);
  and (_19597_, _19548_, _06541_);
  and (_19599_, _19597_, _19592_);
  or (_19600_, _19599_, _06383_);
  or (_19601_, _19600_, _19596_);
  and (_19602_, _14821_, _07923_);
  or (_19603_, _19539_, _07231_);
  or (_19604_, _19603_, _19602_);
  and (_19605_, _19604_, _07229_);
  and (_19606_, _19605_, _19601_);
  nor (_19607_, _11213_, _11326_);
  or (_19608_, _19607_, _19539_);
  and (_19610_, _19608_, _06528_);
  or (_19611_, _19610_, _19606_);
  and (_19612_, _19611_, _07241_);
  and (_19613_, _19545_, _06563_);
  or (_19614_, _19613_, _06188_);
  or (_19615_, _19614_, _19612_);
  and (_19616_, _14884_, _07923_);
  or (_19617_, _19539_, _06189_);
  or (_19618_, _19617_, _19616_);
  and (_19619_, _19618_, _01452_);
  and (_19621_, _19619_, _19615_);
  or (_19622_, _19621_, _19538_);
  and (_43780_, _19622_, _43223_);
  and (_19623_, _11326_, \oc8051_golden_model_1.PCON [3]);
  and (_19624_, _14898_, _07923_);
  or (_19625_, _19624_, _19623_);
  or (_19626_, _19625_, _06252_);
  and (_19627_, _07923_, \oc8051_golden_model_1.ACC [3]);
  or (_19628_, _19627_, _19623_);
  and (_19629_, _19628_, _07123_);
  and (_19631_, _07124_, \oc8051_golden_model_1.PCON [3]);
  or (_19632_, _19631_, _06251_);
  or (_19633_, _19632_, _19629_);
  and (_19634_, _19633_, _07142_);
  and (_19635_, _19634_, _19626_);
  nor (_19636_, _11326_, _07713_);
  or (_19637_, _19636_, _19623_);
  and (_19638_, _19637_, _06468_);
  or (_19639_, _19638_, _19635_);
  and (_19640_, _19639_, _06801_);
  and (_19642_, _19628_, _06466_);
  or (_19643_, _19642_, _07187_);
  or (_19644_, _19643_, _19640_);
  or (_19645_, _19637_, _07188_);
  and (_19646_, _19645_, _07183_);
  and (_19647_, _19646_, _19644_);
  and (_19648_, _09205_, _07923_);
  or (_19649_, _19648_, _19623_);
  and (_19650_, _19649_, _07182_);
  or (_19651_, _19650_, _05968_);
  or (_19653_, _19651_, _19647_);
  and (_19654_, _15003_, _07923_);
  or (_19655_, _19623_, _06336_);
  or (_19656_, _19655_, _19654_);
  and (_19657_, _19656_, _07198_);
  and (_19658_, _19657_, _19653_);
  and (_19659_, _07923_, _08872_);
  or (_19660_, _19659_, _19623_);
  and (_19661_, _19660_, _06371_);
  or (_19662_, _19661_, _06367_);
  or (_19664_, _19662_, _19658_);
  and (_19665_, _15018_, _07923_);
  or (_19666_, _19665_, _19623_);
  or (_19667_, _19666_, _07218_);
  and (_19668_, _19667_, _07216_);
  and (_19669_, _19668_, _19664_);
  and (_19670_, _12523_, _07923_);
  or (_19671_, _19670_, _19623_);
  and (_19672_, _19671_, _06533_);
  or (_19673_, _19672_, _19669_);
  and (_19675_, _19673_, _07213_);
  or (_19676_, _19623_, _08257_);
  and (_19677_, _19660_, _06366_);
  and (_19678_, _19677_, _19676_);
  or (_19679_, _19678_, _19675_);
  and (_19680_, _19679_, _07210_);
  and (_19681_, _19628_, _06541_);
  and (_19682_, _19681_, _19676_);
  or (_19683_, _19682_, _06383_);
  or (_19684_, _19683_, _19680_);
  and (_19686_, _15015_, _07923_);
  or (_19687_, _19623_, _07231_);
  or (_19688_, _19687_, _19686_);
  and (_19689_, _19688_, _07229_);
  and (_19690_, _19689_, _19684_);
  nor (_19691_, _11211_, _11326_);
  or (_19692_, _19691_, _19623_);
  and (_19693_, _19692_, _06528_);
  or (_19694_, _19693_, _06563_);
  or (_19695_, _19694_, _19690_);
  or (_19697_, _19625_, _07241_);
  and (_19698_, _19697_, _06189_);
  and (_19699_, _19698_, _19695_);
  and (_19700_, _15075_, _07923_);
  or (_19701_, _19700_, _19623_);
  and (_19702_, _19701_, _06188_);
  or (_19703_, _19702_, _01456_);
  or (_19704_, _19703_, _19699_);
  or (_19705_, _01452_, \oc8051_golden_model_1.PCON [3]);
  and (_19706_, _19705_, _43223_);
  and (_43781_, _19706_, _19704_);
  and (_19708_, _11326_, \oc8051_golden_model_1.PCON [4]);
  and (_19709_, _15108_, _07923_);
  or (_19710_, _19709_, _19708_);
  or (_19711_, _19710_, _06252_);
  and (_19712_, _07923_, \oc8051_golden_model_1.ACC [4]);
  or (_19713_, _19712_, _19708_);
  and (_19714_, _19713_, _07123_);
  and (_19715_, _07124_, \oc8051_golden_model_1.PCON [4]);
  or (_19716_, _19715_, _06251_);
  or (_19718_, _19716_, _19714_);
  and (_19719_, _19718_, _07142_);
  and (_19720_, _19719_, _19711_);
  nor (_19721_, _08494_, _11326_);
  or (_19722_, _19721_, _19708_);
  and (_19723_, _19722_, _06468_);
  or (_19724_, _19723_, _19720_);
  and (_19725_, _19724_, _06801_);
  and (_19726_, _19713_, _06466_);
  or (_19727_, _19726_, _07187_);
  or (_19729_, _19727_, _19725_);
  or (_19730_, _19722_, _07188_);
  and (_19731_, _19730_, _19729_);
  or (_19732_, _19731_, _07182_);
  and (_19733_, _09159_, _07923_);
  or (_19734_, _19708_, _07183_);
  or (_19735_, _19734_, _19733_);
  and (_19736_, _19735_, _19732_);
  or (_19737_, _19736_, _05968_);
  and (_19738_, _15198_, _07923_);
  or (_19740_, _19708_, _06336_);
  or (_19741_, _19740_, _19738_);
  and (_19742_, _19741_, _07198_);
  and (_19743_, _19742_, _19737_);
  and (_19744_, _08892_, _07923_);
  or (_19745_, _19744_, _19708_);
  and (_19746_, _19745_, _06371_);
  or (_19747_, _19746_, _06367_);
  or (_19748_, _19747_, _19743_);
  and (_19749_, _15214_, _07923_);
  or (_19752_, _19749_, _19708_);
  or (_19753_, _19752_, _07218_);
  and (_19754_, _19753_, _07216_);
  and (_19755_, _19754_, _19748_);
  and (_19756_, _11209_, _07923_);
  or (_19757_, _19756_, _19708_);
  and (_19758_, _19757_, _06533_);
  or (_19759_, _19758_, _19755_);
  and (_19760_, _19759_, _07213_);
  or (_19761_, _19708_, _08497_);
  and (_19764_, _19745_, _06366_);
  and (_19765_, _19764_, _19761_);
  or (_19766_, _19765_, _19760_);
  and (_19767_, _19766_, _07210_);
  and (_19768_, _19713_, _06541_);
  and (_19769_, _19768_, _19761_);
  or (_19770_, _19769_, _06383_);
  or (_19771_, _19770_, _19767_);
  and (_19772_, _15211_, _07923_);
  or (_19773_, _19708_, _07231_);
  or (_19776_, _19773_, _19772_);
  and (_19777_, _19776_, _07229_);
  and (_19778_, _19777_, _19771_);
  nor (_19779_, _11208_, _11326_);
  or (_19780_, _19779_, _19708_);
  and (_19781_, _19780_, _06528_);
  or (_19782_, _19781_, _06563_);
  or (_19783_, _19782_, _19778_);
  or (_19784_, _19710_, _07241_);
  and (_19785_, _19784_, _06189_);
  and (_19788_, _19785_, _19783_);
  and (_19789_, _15280_, _07923_);
  or (_19790_, _19789_, _19708_);
  and (_19791_, _19790_, _06188_);
  or (_19792_, _19791_, _01456_);
  or (_19793_, _19792_, _19788_);
  or (_19794_, _01452_, \oc8051_golden_model_1.PCON [4]);
  and (_19795_, _19794_, _43223_);
  and (_43782_, _19795_, _19793_);
  and (_19796_, _11326_, \oc8051_golden_model_1.PCON [5]);
  nor (_19799_, _08209_, _11326_);
  or (_19800_, _19799_, _19796_);
  or (_19801_, _19800_, _07188_);
  and (_19802_, _15311_, _07923_);
  or (_19803_, _19802_, _19796_);
  or (_19804_, _19803_, _06252_);
  and (_19805_, _07923_, \oc8051_golden_model_1.ACC [5]);
  or (_19806_, _19805_, _19796_);
  and (_19807_, _19806_, _07123_);
  and (_19808_, _07124_, \oc8051_golden_model_1.PCON [5]);
  or (_19811_, _19808_, _06251_);
  or (_19812_, _19811_, _19807_);
  and (_19813_, _19812_, _07142_);
  and (_19814_, _19813_, _19804_);
  and (_19815_, _19800_, _06468_);
  or (_19816_, _19815_, _19814_);
  and (_19817_, _19816_, _06801_);
  and (_19818_, _19806_, _06466_);
  or (_19819_, _19818_, _07187_);
  or (_19820_, _19819_, _19817_);
  and (_19823_, _19820_, _19801_);
  or (_19824_, _19823_, _07182_);
  and (_19825_, _09113_, _07923_);
  or (_19826_, _19796_, _07183_);
  or (_19827_, _19826_, _19825_);
  and (_19828_, _19827_, _06336_);
  and (_19829_, _19828_, _19824_);
  and (_19830_, _15400_, _07923_);
  or (_19831_, _19830_, _19796_);
  and (_19832_, _19831_, _05968_);
  or (_19834_, _19832_, _06371_);
  or (_19835_, _19834_, _19829_);
  and (_19836_, _08888_, _07923_);
  or (_19837_, _19836_, _19796_);
  or (_19838_, _19837_, _07198_);
  and (_19839_, _19838_, _19835_);
  or (_19840_, _19839_, _06367_);
  and (_19841_, _15416_, _07923_);
  or (_19842_, _19841_, _19796_);
  or (_19843_, _19842_, _07218_);
  and (_19845_, _19843_, _07216_);
  and (_19846_, _19845_, _19840_);
  and (_19847_, _11205_, _07923_);
  or (_19848_, _19847_, _19796_);
  and (_19849_, _19848_, _06533_);
  or (_19850_, _19849_, _19846_);
  and (_19851_, _19850_, _07213_);
  or (_19852_, _19796_, _08212_);
  and (_19853_, _19837_, _06366_);
  and (_19854_, _19853_, _19852_);
  or (_19856_, _19854_, _19851_);
  and (_19857_, _19856_, _07210_);
  and (_19858_, _19806_, _06541_);
  and (_19859_, _19858_, _19852_);
  or (_19860_, _19859_, _06383_);
  or (_19861_, _19860_, _19857_);
  and (_19862_, _15413_, _07923_);
  or (_19863_, _19796_, _07231_);
  or (_19864_, _19863_, _19862_);
  and (_19865_, _19864_, _07229_);
  and (_19867_, _19865_, _19861_);
  nor (_19868_, _11204_, _11326_);
  or (_19869_, _19868_, _19796_);
  and (_19870_, _19869_, _06528_);
  or (_19871_, _19870_, _06563_);
  or (_19872_, _19871_, _19867_);
  or (_19873_, _19803_, _07241_);
  and (_19874_, _19873_, _06189_);
  and (_19875_, _19874_, _19872_);
  and (_19876_, _15477_, _07923_);
  or (_19878_, _19876_, _19796_);
  and (_19879_, _19878_, _06188_);
  or (_19880_, _19879_, _01456_);
  or (_19881_, _19880_, _19875_);
  or (_19882_, _01452_, \oc8051_golden_model_1.PCON [5]);
  and (_19883_, _19882_, _43223_);
  and (_43783_, _19883_, _19881_);
  and (_19884_, _11326_, \oc8051_golden_model_1.PCON [6]);
  and (_19885_, _15512_, _07923_);
  or (_19886_, _19885_, _19884_);
  or (_19888_, _19886_, _06252_);
  and (_19889_, _07923_, \oc8051_golden_model_1.ACC [6]);
  or (_19890_, _19889_, _19884_);
  and (_19891_, _19890_, _07123_);
  and (_19892_, _07124_, \oc8051_golden_model_1.PCON [6]);
  or (_19893_, _19892_, _06251_);
  or (_19894_, _19893_, _19891_);
  and (_19895_, _19894_, _07142_);
  and (_19896_, _19895_, _19888_);
  nor (_19897_, _08106_, _11326_);
  or (_19899_, _19897_, _19884_);
  and (_19900_, _19899_, _06468_);
  or (_19901_, _19900_, _19896_);
  and (_19902_, _19901_, _06801_);
  and (_19903_, _19890_, _06466_);
  or (_19904_, _19903_, _07187_);
  or (_19905_, _19904_, _19902_);
  or (_19906_, _19899_, _07188_);
  and (_19907_, _19906_, _19905_);
  or (_19908_, _19907_, _07182_);
  and (_19910_, _09067_, _07923_);
  or (_19911_, _19884_, _07183_);
  or (_19912_, _19911_, _19910_);
  and (_19913_, _19912_, _06336_);
  and (_19914_, _19913_, _19908_);
  and (_19915_, _15601_, _07923_);
  or (_19916_, _19915_, _19884_);
  and (_19917_, _19916_, _05968_);
  or (_19918_, _19917_, _06371_);
  or (_19919_, _19918_, _19914_);
  and (_19921_, _15608_, _07923_);
  or (_19922_, _19921_, _19884_);
  or (_19923_, _19922_, _07198_);
  and (_19924_, _19923_, _19919_);
  or (_19925_, _19924_, _06367_);
  and (_19926_, _15618_, _07923_);
  or (_19927_, _19926_, _19884_);
  or (_19928_, _19927_, _07218_);
  and (_19929_, _19928_, _07216_);
  and (_19930_, _19929_, _19925_);
  and (_19932_, _11202_, _07923_);
  or (_19933_, _19932_, _19884_);
  and (_19934_, _19933_, _06533_);
  or (_19935_, _19934_, _19930_);
  and (_19936_, _19935_, _07213_);
  or (_19937_, _19884_, _08109_);
  and (_19938_, _19922_, _06366_);
  and (_19939_, _19938_, _19937_);
  or (_19940_, _19939_, _19936_);
  and (_19941_, _19940_, _07210_);
  and (_19943_, _19890_, _06541_);
  and (_19944_, _19943_, _19937_);
  or (_19945_, _19944_, _06383_);
  or (_19946_, _19945_, _19941_);
  and (_19947_, _15615_, _07923_);
  or (_19948_, _19884_, _07231_);
  or (_19949_, _19948_, _19947_);
  and (_19950_, _19949_, _07229_);
  and (_19951_, _19950_, _19946_);
  nor (_19952_, _11201_, _11326_);
  or (_19954_, _19952_, _19884_);
  and (_19955_, _19954_, _06528_);
  or (_19956_, _19955_, _06563_);
  or (_19957_, _19956_, _19951_);
  or (_19958_, _19886_, _07241_);
  and (_19959_, _19958_, _06189_);
  and (_19960_, _19959_, _19957_);
  and (_19961_, _15676_, _07923_);
  or (_19962_, _19961_, _19884_);
  and (_19963_, _19962_, _06188_);
  or (_19965_, _19963_, _01456_);
  or (_19966_, _19965_, _19960_);
  or (_19967_, _01452_, \oc8051_golden_model_1.PCON [6]);
  and (_19968_, _19967_, _43223_);
  and (_43784_, _19968_, _19966_);
  not (_19969_, \oc8051_golden_model_1.TMOD [0]);
  nor (_19970_, _01452_, _19969_);
  nand (_19971_, _11218_, _07885_);
  nor (_19972_, _07885_, _19969_);
  nor (_19973_, _19972_, _07210_);
  nand (_19975_, _19973_, _19971_);
  nor (_19976_, _08351_, _11404_);
  or (_19977_, _19976_, _19972_);
  or (_19978_, _19977_, _06252_);
  and (_19979_, _07885_, \oc8051_golden_model_1.ACC [0]);
  or (_19980_, _19979_, _19972_);
  and (_19981_, _19980_, _07123_);
  nor (_19982_, _07123_, _19969_);
  or (_19983_, _19982_, _06251_);
  or (_19984_, _19983_, _19981_);
  and (_19986_, _19984_, _07142_);
  and (_19987_, _19986_, _19978_);
  and (_19988_, _07885_, _07325_);
  or (_19989_, _19988_, _19972_);
  and (_19990_, _19989_, _06468_);
  or (_19991_, _19990_, _19987_);
  and (_19992_, _19991_, _06801_);
  and (_19993_, _19980_, _06466_);
  or (_19994_, _19993_, _07187_);
  or (_19995_, _19994_, _19992_);
  or (_19997_, _19989_, _07188_);
  and (_19998_, _19997_, _19995_);
  or (_19999_, _19998_, _07182_);
  and (_20000_, _09342_, _07885_);
  or (_20001_, _19972_, _07183_);
  or (_20002_, _20001_, _20000_);
  and (_20003_, _20002_, _19999_);
  or (_20004_, _20003_, _05968_);
  and (_20005_, _14427_, _07885_);
  or (_20006_, _19972_, _06336_);
  or (_20008_, _20006_, _20005_);
  and (_20009_, _20008_, _07198_);
  and (_20010_, _20009_, _20004_);
  and (_20011_, _07885_, _08908_);
  or (_20012_, _20011_, _19972_);
  and (_20013_, _20012_, _06371_);
  or (_20014_, _20013_, _06367_);
  or (_20015_, _20014_, _20010_);
  and (_20016_, _14442_, _07885_);
  or (_20017_, _20016_, _19972_);
  or (_20019_, _20017_, _07218_);
  and (_20020_, _20019_, _07216_);
  and (_20021_, _20020_, _20015_);
  nor (_20022_, _12526_, _11404_);
  or (_20023_, _20022_, _19972_);
  and (_20024_, _19971_, _06533_);
  and (_20025_, _20024_, _20023_);
  or (_20026_, _20025_, _20021_);
  and (_20027_, _20026_, _07213_);
  nand (_20028_, _20012_, _06366_);
  nor (_20030_, _20028_, _19976_);
  or (_20031_, _20030_, _06541_);
  or (_20032_, _20031_, _20027_);
  and (_20033_, _20032_, _19975_);
  or (_20034_, _20033_, _06383_);
  and (_20035_, _14325_, _07885_);
  or (_20036_, _19972_, _07231_);
  or (_20037_, _20036_, _20035_);
  and (_20038_, _20037_, _07229_);
  and (_20039_, _20038_, _20034_);
  and (_20041_, _20023_, _06528_);
  or (_20042_, _20041_, _19442_);
  or (_20043_, _20042_, _20039_);
  or (_20044_, _19977_, _06756_);
  and (_20045_, _20044_, _01452_);
  and (_20046_, _20045_, _20043_);
  or (_20047_, _20046_, _19970_);
  and (_43786_, _20047_, _43223_);
  and (_20048_, _11404_, \oc8051_golden_model_1.TMOD [1]);
  nor (_20049_, _11216_, _11404_);
  or (_20051_, _20049_, _20048_);
  or (_20052_, _20051_, _07229_);
  or (_20053_, _07885_, \oc8051_golden_model_1.TMOD [1]);
  and (_20054_, _14503_, _07885_);
  not (_20055_, _20054_);
  and (_20056_, _20055_, _20053_);
  or (_20057_, _20056_, _06252_);
  and (_20058_, _07885_, \oc8051_golden_model_1.ACC [1]);
  or (_20059_, _20058_, _20048_);
  and (_20060_, _20059_, _07123_);
  and (_20062_, _07124_, \oc8051_golden_model_1.TMOD [1]);
  or (_20063_, _20062_, _06251_);
  or (_20064_, _20063_, _20060_);
  and (_20065_, _20064_, _07142_);
  and (_20066_, _20065_, _20057_);
  nor (_20067_, _11404_, _07120_);
  or (_20068_, _20067_, _20048_);
  and (_20069_, _20068_, _06468_);
  or (_20070_, _20069_, _20066_);
  and (_20071_, _20070_, _06801_);
  and (_20073_, _20059_, _06466_);
  or (_20074_, _20073_, _07187_);
  or (_20075_, _20074_, _20071_);
  or (_20076_, _20068_, _07188_);
  and (_20077_, _20076_, _07183_);
  and (_20078_, _20077_, _20075_);
  or (_20079_, _09297_, _11404_);
  and (_20080_, _20053_, _07182_);
  and (_20081_, _20080_, _20079_);
  or (_20082_, _20081_, _20078_);
  and (_20084_, _20082_, _06336_);
  or (_20085_, _14609_, _11404_);
  and (_20086_, _20053_, _05968_);
  and (_20087_, _20086_, _20085_);
  or (_20088_, _20087_, _20084_);
  and (_20089_, _20088_, _07198_);
  nand (_20090_, _07885_, _07018_);
  and (_20091_, _20053_, _06371_);
  and (_20092_, _20091_, _20090_);
  or (_20093_, _20092_, _20089_);
  and (_20095_, _20093_, _07218_);
  or (_20096_, _14625_, _11404_);
  and (_20097_, _20053_, _06367_);
  and (_20098_, _20097_, _20096_);
  or (_20099_, _20098_, _06533_);
  or (_20100_, _20099_, _20095_);
  and (_20101_, _11217_, _07885_);
  or (_20102_, _20101_, _20048_);
  or (_20103_, _20102_, _07216_);
  and (_20104_, _20103_, _07213_);
  and (_20106_, _20104_, _20100_);
  or (_20107_, _14623_, _11404_);
  and (_20108_, _20053_, _06366_);
  and (_20109_, _20108_, _20107_);
  or (_20110_, _20109_, _06541_);
  or (_20111_, _20110_, _20106_);
  and (_20112_, _20058_, _08302_);
  or (_20113_, _20048_, _07210_);
  or (_20114_, _20113_, _20112_);
  and (_20115_, _20114_, _07231_);
  and (_20117_, _20115_, _20111_);
  or (_20118_, _20090_, _08302_);
  and (_20119_, _20053_, _06383_);
  and (_20120_, _20119_, _20118_);
  or (_20121_, _20120_, _06528_);
  or (_20122_, _20121_, _20117_);
  and (_20123_, _20122_, _20052_);
  or (_20124_, _20123_, _06563_);
  or (_20125_, _20056_, _07241_);
  and (_20126_, _20125_, _06189_);
  and (_20128_, _20126_, _20124_);
  or (_20129_, _20054_, _20048_);
  and (_20130_, _20129_, _06188_);
  or (_20131_, _20130_, _01456_);
  or (_20132_, _20131_, _20128_);
  or (_20133_, _01452_, \oc8051_golden_model_1.TMOD [1]);
  and (_20134_, _20133_, _43223_);
  and (_43787_, _20134_, _20132_);
  and (_20135_, _01456_, \oc8051_golden_model_1.TMOD [2]);
  and (_20136_, _11404_, \oc8051_golden_model_1.TMOD [2]);
  and (_20138_, _09251_, _07885_);
  or (_20139_, _20138_, _20136_);
  and (_20140_, _20139_, _07182_);
  and (_20141_, _14712_, _07885_);
  or (_20142_, _20141_, _20136_);
  or (_20143_, _20142_, _06252_);
  and (_20144_, _07885_, \oc8051_golden_model_1.ACC [2]);
  or (_20145_, _20144_, _20136_);
  and (_20146_, _20145_, _07123_);
  and (_20147_, _07124_, \oc8051_golden_model_1.TMOD [2]);
  or (_20149_, _20147_, _06251_);
  or (_20150_, _20149_, _20146_);
  and (_20151_, _20150_, _07142_);
  and (_20152_, _20151_, _20143_);
  nor (_20153_, _11404_, _07578_);
  or (_20154_, _20153_, _20136_);
  and (_20155_, _20154_, _06468_);
  or (_20156_, _20155_, _20152_);
  and (_20157_, _20156_, _06801_);
  and (_20158_, _20145_, _06466_);
  or (_20160_, _20158_, _07187_);
  or (_20161_, _20160_, _20157_);
  or (_20162_, _20154_, _07188_);
  and (_20163_, _20162_, _07183_);
  and (_20164_, _20163_, _20161_);
  or (_20165_, _20164_, _05968_);
  or (_20166_, _20165_, _20140_);
  and (_20167_, _14808_, _07885_);
  or (_20168_, _20136_, _06336_);
  or (_20169_, _20168_, _20167_);
  and (_20171_, _20169_, _07198_);
  and (_20172_, _20171_, _20166_);
  and (_20173_, _07885_, _08945_);
  or (_20174_, _20173_, _20136_);
  and (_20175_, _20174_, _06371_);
  or (_20176_, _20175_, _06367_);
  or (_20177_, _20176_, _20172_);
  and (_20178_, _14824_, _07885_);
  or (_20179_, _20178_, _20136_);
  or (_20180_, _20179_, _07218_);
  and (_20182_, _20180_, _07216_);
  and (_20183_, _20182_, _20177_);
  and (_20184_, _11214_, _07885_);
  or (_20185_, _20184_, _20136_);
  and (_20186_, _20185_, _06533_);
  or (_20187_, _20186_, _20183_);
  and (_20188_, _20187_, _07213_);
  or (_20189_, _20136_, _08397_);
  and (_20190_, _20174_, _06366_);
  and (_20191_, _20190_, _20189_);
  or (_20193_, _20191_, _20188_);
  and (_20194_, _20193_, _07210_);
  and (_20195_, _20145_, _06541_);
  and (_20196_, _20195_, _20189_);
  or (_20197_, _20196_, _06383_);
  or (_20198_, _20197_, _20194_);
  and (_20199_, _14821_, _07885_);
  or (_20200_, _20136_, _07231_);
  or (_20201_, _20200_, _20199_);
  and (_20202_, _20201_, _07229_);
  and (_20204_, _20202_, _20198_);
  nor (_20205_, _11213_, _11404_);
  or (_20206_, _20205_, _20136_);
  and (_20207_, _20206_, _06528_);
  or (_20208_, _20207_, _20204_);
  and (_20209_, _20208_, _07241_);
  and (_20210_, _20142_, _06563_);
  or (_20211_, _20210_, _06188_);
  or (_20212_, _20211_, _20209_);
  and (_20213_, _14884_, _07885_);
  or (_20215_, _20136_, _06189_);
  or (_20216_, _20215_, _20213_);
  and (_20217_, _20216_, _01452_);
  and (_20218_, _20217_, _20212_);
  or (_20219_, _20218_, _20135_);
  and (_43788_, _20219_, _43223_);
  and (_20220_, _11404_, \oc8051_golden_model_1.TMOD [3]);
  and (_20221_, _14898_, _07885_);
  or (_20222_, _20221_, _20220_);
  or (_20223_, _20222_, _06252_);
  and (_20225_, _07885_, \oc8051_golden_model_1.ACC [3]);
  or (_20226_, _20225_, _20220_);
  and (_20227_, _20226_, _07123_);
  and (_20228_, _07124_, \oc8051_golden_model_1.TMOD [3]);
  or (_20229_, _20228_, _06251_);
  or (_20230_, _20229_, _20227_);
  and (_20231_, _20230_, _07142_);
  and (_20232_, _20231_, _20223_);
  nor (_20233_, _11404_, _07713_);
  or (_20234_, _20233_, _20220_);
  and (_20236_, _20234_, _06468_);
  or (_20237_, _20236_, _20232_);
  and (_20238_, _20237_, _06801_);
  and (_20239_, _20226_, _06466_);
  or (_20240_, _20239_, _07187_);
  or (_20241_, _20240_, _20238_);
  or (_20242_, _20234_, _07188_);
  and (_20243_, _20242_, _07183_);
  and (_20244_, _20243_, _20241_);
  and (_20245_, _09205_, _07885_);
  or (_20247_, _20245_, _20220_);
  and (_20248_, _20247_, _07182_);
  or (_20249_, _20248_, _05968_);
  or (_20250_, _20249_, _20244_);
  and (_20251_, _15003_, _07885_);
  or (_20252_, _20220_, _06336_);
  or (_20253_, _20252_, _20251_);
  and (_20254_, _20253_, _07198_);
  and (_20255_, _20254_, _20250_);
  and (_20256_, _07885_, _08872_);
  or (_20258_, _20256_, _20220_);
  and (_20259_, _20258_, _06371_);
  or (_20260_, _20259_, _06367_);
  or (_20261_, _20260_, _20255_);
  and (_20262_, _15018_, _07885_);
  or (_20263_, _20262_, _20220_);
  or (_20264_, _20263_, _07218_);
  and (_20265_, _20264_, _07216_);
  and (_20266_, _20265_, _20261_);
  and (_20267_, _12523_, _07885_);
  or (_20269_, _20267_, _20220_);
  and (_20270_, _20269_, _06533_);
  or (_20271_, _20270_, _20266_);
  and (_20272_, _20271_, _07213_);
  or (_20273_, _20220_, _08257_);
  and (_20274_, _20258_, _06366_);
  and (_20275_, _20274_, _20273_);
  or (_20276_, _20275_, _20272_);
  and (_20277_, _20276_, _07210_);
  and (_20278_, _20226_, _06541_);
  and (_20280_, _20278_, _20273_);
  or (_20281_, _20280_, _06383_);
  or (_20282_, _20281_, _20277_);
  and (_20283_, _15015_, _07885_);
  or (_20284_, _20220_, _07231_);
  or (_20285_, _20284_, _20283_);
  and (_20286_, _20285_, _07229_);
  and (_20287_, _20286_, _20282_);
  nor (_20288_, _11211_, _11404_);
  or (_20289_, _20288_, _20220_);
  and (_20291_, _20289_, _06528_);
  or (_20292_, _20291_, _06563_);
  or (_20293_, _20292_, _20287_);
  or (_20294_, _20222_, _07241_);
  and (_20295_, _20294_, _06189_);
  and (_20296_, _20295_, _20293_);
  and (_20297_, _15075_, _07885_);
  or (_20298_, _20297_, _20220_);
  and (_20299_, _20298_, _06188_);
  or (_20300_, _20299_, _01456_);
  or (_20302_, _20300_, _20296_);
  or (_20303_, _01452_, \oc8051_golden_model_1.TMOD [3]);
  and (_20304_, _20303_, _43223_);
  and (_43790_, _20304_, _20302_);
  and (_20305_, _11404_, \oc8051_golden_model_1.TMOD [4]);
  and (_20306_, _15108_, _07885_);
  or (_20307_, _20306_, _20305_);
  or (_20308_, _20307_, _06252_);
  and (_20309_, _07885_, \oc8051_golden_model_1.ACC [4]);
  or (_20310_, _20309_, _20305_);
  and (_20312_, _20310_, _07123_);
  and (_20313_, _07124_, \oc8051_golden_model_1.TMOD [4]);
  or (_20314_, _20313_, _06251_);
  or (_20315_, _20314_, _20312_);
  and (_20316_, _20315_, _07142_);
  and (_20317_, _20316_, _20308_);
  nor (_20318_, _08494_, _11404_);
  or (_20319_, _20318_, _20305_);
  and (_20320_, _20319_, _06468_);
  or (_20321_, _20320_, _20317_);
  and (_20323_, _20321_, _06801_);
  and (_20324_, _20310_, _06466_);
  or (_20325_, _20324_, _07187_);
  or (_20326_, _20325_, _20323_);
  or (_20327_, _20319_, _07188_);
  and (_20328_, _20327_, _20326_);
  or (_20329_, _20328_, _07182_);
  and (_20330_, _09159_, _07885_);
  or (_20331_, _20305_, _07183_);
  or (_20332_, _20331_, _20330_);
  and (_20334_, _20332_, _20329_);
  or (_20335_, _20334_, _05968_);
  and (_20336_, _15198_, _07885_);
  or (_20337_, _20305_, _06336_);
  or (_20338_, _20337_, _20336_);
  and (_20339_, _20338_, _07198_);
  and (_20340_, _20339_, _20335_);
  and (_20341_, _08892_, _07885_);
  or (_20342_, _20341_, _20305_);
  and (_20343_, _20342_, _06371_);
  or (_20345_, _20343_, _06367_);
  or (_20346_, _20345_, _20340_);
  and (_20347_, _15214_, _07885_);
  or (_20348_, _20347_, _20305_);
  or (_20349_, _20348_, _07218_);
  and (_20350_, _20349_, _07216_);
  and (_20351_, _20350_, _20346_);
  and (_20352_, _11209_, _07885_);
  or (_20353_, _20352_, _20305_);
  and (_20354_, _20353_, _06533_);
  or (_20356_, _20354_, _20351_);
  and (_20357_, _20356_, _07213_);
  or (_20358_, _20305_, _08497_);
  and (_20359_, _20342_, _06366_);
  and (_20360_, _20359_, _20358_);
  or (_20361_, _20360_, _20357_);
  and (_20362_, _20361_, _07210_);
  and (_20363_, _20310_, _06541_);
  and (_20364_, _20363_, _20358_);
  or (_20365_, _20364_, _06383_);
  or (_20367_, _20365_, _20362_);
  and (_20368_, _15211_, _07885_);
  or (_20369_, _20305_, _07231_);
  or (_20370_, _20369_, _20368_);
  and (_20371_, _20370_, _07229_);
  and (_20372_, _20371_, _20367_);
  nor (_20373_, _11208_, _11404_);
  or (_20374_, _20373_, _20305_);
  and (_20375_, _20374_, _06528_);
  or (_20376_, _20375_, _06563_);
  or (_20378_, _20376_, _20372_);
  or (_20379_, _20307_, _07241_);
  and (_20380_, _20379_, _06189_);
  and (_20381_, _20380_, _20378_);
  and (_20382_, _15280_, _07885_);
  or (_20383_, _20382_, _20305_);
  and (_20384_, _20383_, _06188_);
  or (_20385_, _20384_, _01456_);
  or (_20386_, _20385_, _20381_);
  or (_20387_, _01452_, \oc8051_golden_model_1.TMOD [4]);
  and (_20389_, _20387_, _43223_);
  and (_43791_, _20389_, _20386_);
  and (_20390_, _11404_, \oc8051_golden_model_1.TMOD [5]);
  nor (_20391_, _08209_, _11404_);
  or (_20392_, _20391_, _20390_);
  or (_20393_, _20392_, _07188_);
  and (_20394_, _15311_, _07885_);
  or (_20395_, _20394_, _20390_);
  or (_20396_, _20395_, _06252_);
  and (_20397_, _07885_, \oc8051_golden_model_1.ACC [5]);
  or (_20399_, _20397_, _20390_);
  and (_20400_, _20399_, _07123_);
  and (_20401_, _07124_, \oc8051_golden_model_1.TMOD [5]);
  or (_20402_, _20401_, _06251_);
  or (_20403_, _20402_, _20400_);
  and (_20404_, _20403_, _07142_);
  and (_20405_, _20404_, _20396_);
  and (_20406_, _20392_, _06468_);
  or (_20407_, _20406_, _20405_);
  and (_20408_, _20407_, _06801_);
  and (_20410_, _20399_, _06466_);
  or (_20411_, _20410_, _07187_);
  or (_20412_, _20411_, _20408_);
  and (_20413_, _20412_, _20393_);
  or (_20414_, _20413_, _07182_);
  and (_20415_, _09113_, _07885_);
  or (_20416_, _20390_, _07183_);
  or (_20417_, _20416_, _20415_);
  and (_20418_, _20417_, _06336_);
  and (_20419_, _20418_, _20414_);
  and (_20421_, _15400_, _07885_);
  or (_20422_, _20421_, _20390_);
  and (_20423_, _20422_, _05968_);
  or (_20424_, _20423_, _06371_);
  or (_20425_, _20424_, _20419_);
  and (_20426_, _08888_, _07885_);
  or (_20427_, _20426_, _20390_);
  or (_20428_, _20427_, _07198_);
  and (_20429_, _20428_, _20425_);
  or (_20430_, _20429_, _06367_);
  and (_20432_, _15416_, _07885_);
  or (_20433_, _20432_, _20390_);
  or (_20434_, _20433_, _07218_);
  and (_20435_, _20434_, _07216_);
  and (_20436_, _20435_, _20430_);
  and (_20437_, _11205_, _07885_);
  or (_20438_, _20437_, _20390_);
  and (_20439_, _20438_, _06533_);
  or (_20440_, _20439_, _20436_);
  and (_20441_, _20440_, _07213_);
  or (_20443_, _20390_, _08212_);
  and (_20444_, _20427_, _06366_);
  and (_20445_, _20444_, _20443_);
  or (_20446_, _20445_, _20441_);
  and (_20447_, _20446_, _07210_);
  and (_20448_, _20399_, _06541_);
  and (_20449_, _20448_, _20443_);
  or (_20450_, _20449_, _06383_);
  or (_20451_, _20450_, _20447_);
  and (_20452_, _15413_, _07885_);
  or (_20454_, _20390_, _07231_);
  or (_20455_, _20454_, _20452_);
  and (_20456_, _20455_, _07229_);
  and (_20457_, _20456_, _20451_);
  nor (_20458_, _11204_, _11404_);
  or (_20459_, _20458_, _20390_);
  and (_20460_, _20459_, _06528_);
  or (_20461_, _20460_, _06563_);
  or (_20462_, _20461_, _20457_);
  or (_20463_, _20395_, _07241_);
  and (_20465_, _20463_, _06189_);
  and (_20466_, _20465_, _20462_);
  and (_20467_, _15477_, _07885_);
  or (_20468_, _20467_, _20390_);
  and (_20469_, _20468_, _06188_);
  or (_20470_, _20469_, _01456_);
  or (_20471_, _20470_, _20466_);
  or (_20472_, _01452_, \oc8051_golden_model_1.TMOD [5]);
  and (_20473_, _20472_, _43223_);
  and (_43792_, _20473_, _20471_);
  and (_20475_, _11404_, \oc8051_golden_model_1.TMOD [6]);
  nor (_20476_, _08106_, _11404_);
  or (_20477_, _20476_, _20475_);
  or (_20478_, _20477_, _07188_);
  and (_20479_, _15512_, _07885_);
  or (_20480_, _20479_, _20475_);
  or (_20481_, _20480_, _06252_);
  and (_20482_, _07885_, \oc8051_golden_model_1.ACC [6]);
  or (_20483_, _20482_, _20475_);
  and (_20484_, _20483_, _07123_);
  and (_20486_, _07124_, \oc8051_golden_model_1.TMOD [6]);
  or (_20487_, _20486_, _06251_);
  or (_20488_, _20487_, _20484_);
  and (_20489_, _20488_, _07142_);
  and (_20490_, _20489_, _20481_);
  and (_20491_, _20477_, _06468_);
  or (_20492_, _20491_, _20490_);
  and (_20493_, _20492_, _06801_);
  and (_20494_, _20483_, _06466_);
  or (_20495_, _20494_, _07187_);
  or (_20497_, _20495_, _20493_);
  and (_20498_, _20497_, _20478_);
  or (_20499_, _20498_, _07182_);
  and (_20500_, _09067_, _07885_);
  or (_20501_, _20475_, _07183_);
  or (_20502_, _20501_, _20500_);
  and (_20503_, _20502_, _06336_);
  and (_20504_, _20503_, _20499_);
  and (_20505_, _15601_, _07885_);
  or (_20506_, _20505_, _20475_);
  and (_20508_, _20506_, _05968_);
  or (_20509_, _20508_, _06371_);
  or (_20510_, _20509_, _20504_);
  and (_20511_, _15608_, _07885_);
  or (_20512_, _20511_, _20475_);
  or (_20513_, _20512_, _07198_);
  and (_20514_, _20513_, _20510_);
  or (_20515_, _20514_, _06367_);
  and (_20516_, _15618_, _07885_);
  or (_20517_, _20516_, _20475_);
  or (_20519_, _20517_, _07218_);
  and (_20520_, _20519_, _07216_);
  and (_20521_, _20520_, _20515_);
  and (_20522_, _11202_, _07885_);
  or (_20523_, _20522_, _20475_);
  and (_20524_, _20523_, _06533_);
  or (_20525_, _20524_, _20521_);
  and (_20526_, _20525_, _07213_);
  or (_20527_, _20475_, _08109_);
  and (_20528_, _20512_, _06366_);
  and (_20530_, _20528_, _20527_);
  or (_20531_, _20530_, _20526_);
  and (_20532_, _20531_, _07210_);
  and (_20533_, _20483_, _06541_);
  and (_20534_, _20533_, _20527_);
  or (_20535_, _20534_, _06383_);
  or (_20536_, _20535_, _20532_);
  and (_20537_, _15615_, _07885_);
  or (_20538_, _20475_, _07231_);
  or (_20539_, _20538_, _20537_);
  and (_20541_, _20539_, _07229_);
  and (_20542_, _20541_, _20536_);
  nor (_20543_, _11201_, _11404_);
  or (_20544_, _20543_, _20475_);
  and (_20545_, _20544_, _06528_);
  or (_20546_, _20545_, _06563_);
  or (_20547_, _20546_, _20542_);
  or (_20548_, _20480_, _07241_);
  and (_20549_, _20548_, _06189_);
  and (_20550_, _20549_, _20547_);
  and (_20552_, _15676_, _07885_);
  or (_20553_, _20552_, _20475_);
  and (_20554_, _20553_, _06188_);
  or (_20555_, _20554_, _01456_);
  or (_20556_, _20555_, _20550_);
  or (_20557_, _01452_, \oc8051_golden_model_1.TMOD [6]);
  and (_20558_, _20557_, _43223_);
  and (_43793_, _20558_, _20556_);
  not (_20559_, \oc8051_golden_model_1.DPL [0]);
  nor (_20560_, _01452_, _20559_);
  and (_20562_, _07932_, \oc8051_golden_model_1.ACC [0]);
  and (_20563_, _20562_, _08351_);
  nor (_20564_, _07932_, _20559_);
  or (_20565_, _20564_, _07210_);
  or (_20566_, _20565_, _20563_);
  and (_20567_, _07932_, _07325_);
  or (_20568_, _20567_, _20564_);
  or (_20569_, _20568_, _07188_);
  or (_20570_, _20564_, _20562_);
  or (_20571_, _20570_, _06801_);
  nor (_20573_, _08351_, _11487_);
  or (_20574_, _20573_, _20564_);
  or (_20575_, _20574_, _06252_);
  and (_20576_, _20570_, _07123_);
  nor (_20577_, _07123_, _20559_);
  or (_20578_, _20577_, _06251_);
  or (_20579_, _20578_, _20576_);
  and (_20580_, _20579_, _07142_);
  and (_20581_, _20580_, _20575_);
  and (_20582_, _20568_, _06468_);
  or (_20584_, _20582_, _06466_);
  or (_20585_, _20584_, _20581_);
  and (_20586_, _20585_, _20571_);
  or (_20587_, _20586_, _11505_);
  nand (_20588_, _11505_, \oc8051_golden_model_1.DPL [0]);
  and (_20589_, _20588_, _06370_);
  and (_20590_, _20589_, _20587_);
  nor (_20591_, _06912_, _06370_);
  or (_20592_, _20591_, _07187_);
  or (_20593_, _20592_, _20590_);
  and (_20595_, _20593_, _20569_);
  or (_20596_, _20595_, _07182_);
  and (_20597_, _09342_, _07932_);
  or (_20598_, _20564_, _07183_);
  or (_20599_, _20598_, _20597_);
  and (_20600_, _20599_, _20596_);
  or (_20601_, _20600_, _05968_);
  and (_20602_, _14427_, _07932_);
  or (_20603_, _20564_, _06336_);
  or (_20604_, _20603_, _20602_);
  and (_20606_, _20604_, _07198_);
  and (_20607_, _20606_, _20601_);
  and (_20608_, _07932_, _08908_);
  or (_20609_, _20608_, _20564_);
  and (_20610_, _20609_, _06371_);
  or (_20611_, _20610_, _06367_);
  or (_20612_, _20611_, _20607_);
  and (_20613_, _14442_, _07932_);
  or (_20614_, _20613_, _20564_);
  or (_20615_, _20614_, _07218_);
  and (_20617_, _20615_, _07216_);
  and (_20618_, _20617_, _20612_);
  nor (_20619_, _12526_, _11487_);
  or (_20620_, _20619_, _20564_);
  nor (_20621_, _20563_, _07216_);
  and (_20622_, _20621_, _20620_);
  or (_20623_, _20622_, _20618_);
  and (_20624_, _20623_, _07213_);
  nand (_20625_, _20609_, _06366_);
  nor (_20626_, _20625_, _20573_);
  or (_20628_, _20626_, _06541_);
  or (_20629_, _20628_, _20624_);
  and (_20630_, _20629_, _20566_);
  or (_20631_, _20630_, _06383_);
  and (_20632_, _14325_, _07932_);
  or (_20633_, _20632_, _20564_);
  or (_20634_, _20633_, _07231_);
  and (_20635_, _20634_, _07229_);
  and (_20636_, _20635_, _20631_);
  and (_20637_, _20620_, _06528_);
  or (_20639_, _20637_, _19442_);
  or (_20640_, _20639_, _20636_);
  or (_20641_, _20574_, _06756_);
  and (_20642_, _20641_, _01452_);
  and (_20643_, _20642_, _20640_);
  or (_20644_, _20643_, _20560_);
  and (_43795_, _20644_, _43223_);
  not (_20645_, \oc8051_golden_model_1.DPL [1]);
  nor (_20646_, _01452_, _20645_);
  or (_20647_, _09297_, _11487_);
  or (_20648_, _07932_, \oc8051_golden_model_1.DPL [1]);
  and (_20649_, _20648_, _07182_);
  and (_20650_, _20649_, _20647_);
  and (_20651_, _14503_, _07932_);
  not (_20652_, _20651_);
  and (_20653_, _20652_, _20648_);
  or (_20654_, _20653_, _06252_);
  nor (_20655_, _07932_, _20645_);
  and (_20656_, _07932_, \oc8051_golden_model_1.ACC [1]);
  or (_20657_, _20656_, _20655_);
  and (_20659_, _20657_, _07123_);
  nor (_20660_, _07123_, _20645_);
  or (_20661_, _20660_, _06251_);
  or (_20662_, _20661_, _20659_);
  and (_20663_, _20662_, _07142_);
  and (_20664_, _20663_, _20654_);
  nor (_20665_, _11487_, _07120_);
  or (_20666_, _20665_, _20655_);
  and (_20667_, _20666_, _06468_);
  or (_20668_, _20667_, _06466_);
  or (_20671_, _20668_, _20664_);
  or (_20672_, _20657_, _06801_);
  and (_20673_, _20672_, _11506_);
  and (_20674_, _20673_, _20671_);
  nor (_20675_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_20676_, _20675_, _11510_);
  and (_20677_, _20676_, _11505_);
  or (_20678_, _20677_, _20674_);
  and (_20679_, _20678_, _06370_);
  nor (_20680_, _07018_, _06370_);
  or (_20682_, _20680_, _07187_);
  or (_20683_, _20682_, _20679_);
  or (_20684_, _20666_, _07188_);
  and (_20685_, _20684_, _07183_);
  and (_20686_, _20685_, _20683_);
  or (_20687_, _20686_, _20650_);
  and (_20688_, _20687_, _06336_);
  or (_20689_, _14609_, _11487_);
  and (_20690_, _20648_, _05968_);
  and (_20691_, _20690_, _20689_);
  or (_20692_, _20691_, _20688_);
  and (_20693_, _20692_, _07198_);
  nand (_20694_, _07932_, _07018_);
  and (_20695_, _20648_, _06371_);
  and (_20696_, _20695_, _20694_);
  or (_20697_, _20696_, _20693_);
  and (_20698_, _20697_, _07218_);
  or (_20699_, _14625_, _11487_);
  and (_20700_, _20648_, _06367_);
  and (_20701_, _20700_, _20699_);
  or (_20703_, _20701_, _06533_);
  or (_20704_, _20703_, _20698_);
  nor (_20705_, _11216_, _11487_);
  or (_20706_, _20705_, _20655_);
  nand (_20707_, _11215_, _07932_);
  and (_20708_, _20707_, _20706_);
  or (_20709_, _20708_, _07216_);
  and (_20710_, _20709_, _07213_);
  and (_20711_, _20710_, _20704_);
  or (_20712_, _14623_, _11487_);
  and (_20715_, _20648_, _06366_);
  and (_20716_, _20715_, _20712_);
  or (_20717_, _20716_, _06541_);
  or (_20718_, _20717_, _20711_);
  nor (_20719_, _20655_, _07210_);
  nand (_20720_, _20719_, _20707_);
  and (_20721_, _20720_, _07231_);
  and (_20722_, _20721_, _20718_);
  or (_20723_, _20694_, _08302_);
  and (_20724_, _20648_, _06383_);
  and (_20725_, _20724_, _20723_);
  or (_20726_, _20725_, _06528_);
  or (_20727_, _20726_, _20722_);
  or (_20728_, _20706_, _07229_);
  and (_20729_, _20728_, _07241_);
  and (_20730_, _20729_, _20727_);
  and (_20731_, _20653_, _06563_);
  or (_20732_, _20731_, _06188_);
  or (_20733_, _20732_, _20730_);
  or (_20734_, _20655_, _06189_);
  or (_20736_, _20734_, _20651_);
  and (_20737_, _20736_, _01452_);
  and (_20738_, _20737_, _20733_);
  or (_20739_, _20738_, _20646_);
  and (_43796_, _20739_, _43223_);
  not (_20740_, \oc8051_golden_model_1.DPL [2]);
  nor (_20741_, _01452_, _20740_);
  nor (_20742_, _07932_, _20740_);
  nor (_20743_, _11487_, _07578_);
  or (_20744_, _20743_, _20742_);
  or (_20747_, _20744_, _07188_);
  and (_20748_, _14712_, _07932_);
  or (_20749_, _20748_, _20742_);
  or (_20750_, _20749_, _06252_);
  and (_20751_, _07932_, \oc8051_golden_model_1.ACC [2]);
  or (_20752_, _20751_, _20742_);
  and (_20753_, _20752_, _07123_);
  nor (_20754_, _07123_, _20740_);
  or (_20755_, _20754_, _06251_);
  or (_20756_, _20755_, _20753_);
  and (_20758_, _20756_, _07142_);
  and (_20759_, _20758_, _20750_);
  and (_20760_, _20744_, _06468_);
  or (_20761_, _20760_, _06466_);
  or (_20762_, _20761_, _20759_);
  or (_20763_, _20752_, _06801_);
  and (_20764_, _20763_, _11506_);
  and (_20765_, _20764_, _20762_);
  nor (_20766_, _11510_, \oc8051_golden_model_1.DPL [2]);
  nor (_20767_, _20766_, _11511_);
  and (_20769_, _20767_, _11505_);
  or (_20770_, _20769_, _20765_);
  and (_20771_, _20770_, _06370_);
  nor (_20772_, _06651_, _06370_);
  or (_20773_, _20772_, _07187_);
  or (_20774_, _20773_, _20771_);
  and (_20775_, _20774_, _20747_);
  or (_20776_, _20775_, _07182_);
  and (_20777_, _09251_, _07932_);
  or (_20778_, _20742_, _07183_);
  or (_20780_, _20778_, _20777_);
  and (_20781_, _20780_, _06336_);
  and (_20782_, _20781_, _20776_);
  and (_20783_, _14808_, _07932_);
  or (_20784_, _20783_, _20742_);
  and (_20785_, _20784_, _05968_);
  or (_20786_, _20785_, _06371_);
  or (_20787_, _20786_, _20782_);
  and (_20788_, _07932_, _08945_);
  or (_20789_, _20788_, _20742_);
  or (_20790_, _20789_, _07198_);
  and (_20791_, _20790_, _20787_);
  or (_20792_, _20791_, _06367_);
  and (_20793_, _14824_, _07932_);
  or (_20794_, _20793_, _20742_);
  or (_20795_, _20794_, _07218_);
  and (_20796_, _20795_, _07216_);
  and (_20797_, _20796_, _20792_);
  and (_20798_, _11214_, _07932_);
  or (_20799_, _20798_, _20742_);
  and (_20802_, _20799_, _06533_);
  or (_20803_, _20802_, _20797_);
  and (_20804_, _20803_, _07213_);
  or (_20805_, _20742_, _08397_);
  and (_20806_, _20789_, _06366_);
  and (_20807_, _20806_, _20805_);
  or (_20808_, _20807_, _20804_);
  and (_20809_, _20808_, _07210_);
  and (_20810_, _20752_, _06541_);
  and (_20811_, _20810_, _20805_);
  or (_20813_, _20811_, _06383_);
  or (_20814_, _20813_, _20809_);
  and (_20815_, _14821_, _07932_);
  or (_20816_, _20742_, _07231_);
  or (_20817_, _20816_, _20815_);
  and (_20818_, _20817_, _07229_);
  and (_20819_, _20818_, _20814_);
  nor (_20820_, _11213_, _11487_);
  or (_20821_, _20820_, _20742_);
  and (_20822_, _20821_, _06528_);
  or (_20824_, _20822_, _20819_);
  and (_20825_, _20824_, _07241_);
  and (_20826_, _20749_, _06563_);
  or (_20827_, _20826_, _06188_);
  or (_20828_, _20827_, _20825_);
  and (_20829_, _14884_, _07932_);
  or (_20830_, _20742_, _06189_);
  or (_20831_, _20830_, _20829_);
  and (_20832_, _20831_, _01452_);
  and (_20833_, _20832_, _20828_);
  or (_20835_, _20833_, _20741_);
  and (_43797_, _20835_, _43223_);
  and (_20836_, _11487_, \oc8051_golden_model_1.DPL [3]);
  nor (_20837_, _11487_, _07713_);
  or (_20838_, _20837_, _20836_);
  or (_20839_, _20838_, _07188_);
  and (_20840_, _14898_, _07932_);
  or (_20841_, _20840_, _20836_);
  or (_20842_, _20841_, _06252_);
  and (_20843_, _07932_, \oc8051_golden_model_1.ACC [3]);
  or (_20845_, _20843_, _20836_);
  and (_20846_, _20845_, _07123_);
  and (_20847_, _07124_, \oc8051_golden_model_1.DPL [3]);
  or (_20848_, _20847_, _06251_);
  or (_20849_, _20848_, _20846_);
  and (_20850_, _20849_, _07142_);
  and (_20851_, _20850_, _20842_);
  and (_20852_, _20838_, _06468_);
  or (_20853_, _20852_, _06466_);
  or (_20854_, _20853_, _20851_);
  or (_20856_, _20845_, _06801_);
  and (_20857_, _20856_, _11506_);
  and (_20858_, _20857_, _20854_);
  nor (_20859_, _11511_, \oc8051_golden_model_1.DPL [3]);
  nor (_20860_, _20859_, _11512_);
  and (_20861_, _20860_, _11505_);
  or (_20862_, _20861_, _20858_);
  and (_20863_, _20862_, _06370_);
  nor (_20864_, _06458_, _06370_);
  or (_20865_, _20864_, _07187_);
  or (_20867_, _20865_, _20863_);
  and (_20868_, _20867_, _20839_);
  or (_20869_, _20868_, _07182_);
  and (_20870_, _09205_, _07932_);
  or (_20871_, _20836_, _07183_);
  or (_20872_, _20871_, _20870_);
  and (_20873_, _20872_, _06336_);
  and (_20874_, _20873_, _20869_);
  and (_20875_, _15003_, _07932_);
  or (_20876_, _20875_, _20836_);
  and (_20878_, _20876_, _05968_);
  or (_20879_, _20878_, _06371_);
  or (_20880_, _20879_, _20874_);
  and (_20881_, _07932_, _08872_);
  or (_20882_, _20881_, _20836_);
  or (_20883_, _20882_, _07198_);
  and (_20884_, _20883_, _20880_);
  or (_20885_, _20884_, _06367_);
  and (_20886_, _15018_, _07932_);
  or (_20887_, _20886_, _20836_);
  or (_20889_, _20887_, _07218_);
  and (_20890_, _20889_, _07216_);
  and (_20891_, _20890_, _20885_);
  and (_20892_, _12523_, _07932_);
  or (_20893_, _20892_, _20836_);
  and (_20894_, _20893_, _06533_);
  or (_20895_, _20894_, _20891_);
  and (_20896_, _20895_, _07213_);
  or (_20897_, _20836_, _08257_);
  and (_20898_, _20882_, _06366_);
  and (_20900_, _20898_, _20897_);
  or (_20901_, _20900_, _20896_);
  and (_20902_, _20901_, _07210_);
  and (_20903_, _20845_, _06541_);
  and (_20904_, _20903_, _20897_);
  or (_20905_, _20904_, _06383_);
  or (_20906_, _20905_, _20902_);
  and (_20907_, _15015_, _07932_);
  or (_20908_, _20836_, _07231_);
  or (_20909_, _20908_, _20907_);
  and (_20911_, _20909_, _07229_);
  and (_20912_, _20911_, _20906_);
  nor (_20913_, _11211_, _11487_);
  or (_20914_, _20913_, _20836_);
  and (_20915_, _20914_, _06528_);
  or (_20916_, _20915_, _06563_);
  or (_20917_, _20916_, _20912_);
  or (_20918_, _20841_, _07241_);
  and (_20919_, _20918_, _06189_);
  and (_20920_, _20919_, _20917_);
  and (_20921_, _15075_, _07932_);
  or (_20922_, _20921_, _20836_);
  and (_20923_, _20922_, _06188_);
  or (_20924_, _20923_, _01456_);
  or (_20925_, _20924_, _20920_);
  or (_20926_, _01452_, \oc8051_golden_model_1.DPL [3]);
  and (_20927_, _20926_, _43223_);
  and (_43798_, _20927_, _20925_);
  and (_20928_, _11487_, \oc8051_golden_model_1.DPL [4]);
  nor (_20929_, _08494_, _11487_);
  or (_20932_, _20929_, _20928_);
  or (_20933_, _20932_, _07188_);
  and (_20934_, _15108_, _07932_);
  or (_20935_, _20934_, _20928_);
  or (_20936_, _20935_, _06252_);
  and (_20937_, _07932_, \oc8051_golden_model_1.ACC [4]);
  or (_20938_, _20937_, _20928_);
  and (_20939_, _20938_, _07123_);
  and (_20940_, _07124_, \oc8051_golden_model_1.DPL [4]);
  or (_20941_, _20940_, _06251_);
  or (_20943_, _20941_, _20939_);
  and (_20944_, _20943_, _07142_);
  and (_20945_, _20944_, _20936_);
  and (_20946_, _20932_, _06468_);
  or (_20947_, _20946_, _06466_);
  or (_20948_, _20947_, _20945_);
  or (_20949_, _20938_, _06801_);
  and (_20950_, _20949_, _11506_);
  and (_20951_, _20950_, _20948_);
  nor (_20952_, _11512_, \oc8051_golden_model_1.DPL [4]);
  nor (_20954_, _20952_, _11513_);
  and (_20955_, _20954_, _11505_);
  or (_20956_, _20955_, _20951_);
  and (_20957_, _20956_, _06370_);
  nor (_20958_, _08834_, _06370_);
  or (_20959_, _20958_, _07187_);
  or (_20960_, _20959_, _20957_);
  and (_20961_, _20960_, _20933_);
  or (_20962_, _20961_, _07182_);
  and (_20963_, _09159_, _07932_);
  or (_20965_, _20928_, _07183_);
  or (_20966_, _20965_, _20963_);
  and (_20967_, _20966_, _06336_);
  and (_20968_, _20967_, _20962_);
  and (_20969_, _15198_, _07932_);
  or (_20970_, _20969_, _20928_);
  and (_20971_, _20970_, _05968_);
  or (_20972_, _20971_, _06371_);
  or (_20973_, _20972_, _20968_);
  and (_20974_, _08892_, _07932_);
  or (_20976_, _20974_, _20928_);
  or (_20977_, _20976_, _07198_);
  and (_20978_, _20977_, _20973_);
  or (_20979_, _20978_, _06367_);
  and (_20980_, _15214_, _07932_);
  or (_20981_, _20980_, _20928_);
  or (_20982_, _20981_, _07218_);
  and (_20983_, _20982_, _07216_);
  and (_20984_, _20983_, _20979_);
  and (_20985_, _11209_, _07932_);
  or (_20987_, _20985_, _20928_);
  and (_20988_, _20987_, _06533_);
  or (_20989_, _20988_, _20984_);
  and (_20990_, _20989_, _07213_);
  or (_20991_, _20928_, _08497_);
  and (_20992_, _20976_, _06366_);
  and (_20993_, _20992_, _20991_);
  or (_20994_, _20993_, _20990_);
  and (_20995_, _20994_, _07210_);
  and (_20996_, _20938_, _06541_);
  and (_20998_, _20996_, _20991_);
  or (_20999_, _20998_, _06383_);
  or (_21000_, _20999_, _20995_);
  and (_21001_, _15211_, _07932_);
  or (_21002_, _20928_, _07231_);
  or (_21003_, _21002_, _21001_);
  and (_21004_, _21003_, _07229_);
  and (_21005_, _21004_, _21000_);
  nor (_21006_, _11208_, _11487_);
  or (_21007_, _21006_, _20928_);
  and (_21009_, _21007_, _06528_);
  or (_21010_, _21009_, _06563_);
  or (_21011_, _21010_, _21005_);
  or (_21012_, _20935_, _07241_);
  and (_21013_, _21012_, _06189_);
  and (_21014_, _21013_, _21011_);
  and (_21015_, _15280_, _07932_);
  or (_21016_, _21015_, _20928_);
  and (_21017_, _21016_, _06188_);
  or (_21018_, _21017_, _01456_);
  or (_21020_, _21018_, _21014_);
  or (_21021_, _01452_, \oc8051_golden_model_1.DPL [4]);
  and (_21022_, _21021_, _43223_);
  and (_43799_, _21022_, _21020_);
  and (_21023_, _11487_, \oc8051_golden_model_1.DPL [5]);
  nor (_21024_, _08209_, _11487_);
  or (_21025_, _21024_, _21023_);
  or (_21026_, _21025_, _07188_);
  and (_21027_, _15311_, _07932_);
  or (_21028_, _21027_, _21023_);
  or (_21030_, _21028_, _06252_);
  and (_21031_, _07932_, \oc8051_golden_model_1.ACC [5]);
  or (_21032_, _21031_, _21023_);
  and (_21033_, _21032_, _07123_);
  and (_21034_, _07124_, \oc8051_golden_model_1.DPL [5]);
  or (_21035_, _21034_, _06251_);
  or (_21036_, _21035_, _21033_);
  and (_21037_, _21036_, _07142_);
  and (_21038_, _21037_, _21030_);
  and (_21039_, _21025_, _06468_);
  or (_21041_, _21039_, _06466_);
  or (_21042_, _21041_, _21038_);
  or (_21043_, _21032_, _06801_);
  and (_21044_, _21043_, _11506_);
  and (_21045_, _21044_, _21042_);
  nor (_21046_, _11513_, \oc8051_golden_model_1.DPL [5]);
  nor (_21047_, _21046_, _11514_);
  and (_21048_, _21047_, _11505_);
  or (_21049_, _21048_, _21045_);
  and (_21050_, _21049_, _06370_);
  nor (_21052_, _08867_, _06370_);
  or (_21053_, _21052_, _07187_);
  or (_21054_, _21053_, _21050_);
  and (_21055_, _21054_, _21026_);
  or (_21056_, _21055_, _07182_);
  and (_21057_, _09113_, _07932_);
  or (_21058_, _21023_, _07183_);
  or (_21059_, _21058_, _21057_);
  and (_21060_, _21059_, _06336_);
  and (_21061_, _21060_, _21056_);
  and (_21063_, _15400_, _07932_);
  or (_21064_, _21063_, _21023_);
  and (_21065_, _21064_, _05968_);
  or (_21066_, _21065_, _06371_);
  or (_21067_, _21066_, _21061_);
  and (_21068_, _08888_, _07932_);
  or (_21069_, _21068_, _21023_);
  or (_21070_, _21069_, _07198_);
  and (_21071_, _21070_, _21067_);
  or (_21072_, _21071_, _06367_);
  and (_21074_, _15416_, _07932_);
  or (_21075_, _21074_, _21023_);
  or (_21076_, _21075_, _07218_);
  and (_21077_, _21076_, _07216_);
  and (_21078_, _21077_, _21072_);
  and (_21079_, _11205_, _07932_);
  or (_21080_, _21079_, _21023_);
  and (_21081_, _21080_, _06533_);
  or (_21082_, _21081_, _21078_);
  and (_21083_, _21082_, _07213_);
  or (_21085_, _21023_, _08212_);
  and (_21086_, _21069_, _06366_);
  and (_21087_, _21086_, _21085_);
  or (_21088_, _21087_, _21083_);
  and (_21089_, _21088_, _07210_);
  and (_21090_, _21032_, _06541_);
  and (_21091_, _21090_, _21085_);
  or (_21092_, _21091_, _06383_);
  or (_21093_, _21092_, _21089_);
  and (_21094_, _15413_, _07932_);
  or (_21095_, _21023_, _07231_);
  or (_21096_, _21095_, _21094_);
  and (_21097_, _21096_, _07229_);
  and (_21098_, _21097_, _21093_);
  nor (_21099_, _11204_, _11487_);
  or (_21100_, _21099_, _21023_);
  and (_21101_, _21100_, _06528_);
  or (_21102_, _21101_, _06563_);
  or (_21103_, _21102_, _21098_);
  or (_21104_, _21028_, _07241_);
  and (_21107_, _21104_, _06189_);
  and (_21108_, _21107_, _21103_);
  and (_21109_, _15477_, _07932_);
  or (_21110_, _21109_, _21023_);
  and (_21111_, _21110_, _06188_);
  or (_21112_, _21111_, _01456_);
  or (_21113_, _21112_, _21108_);
  or (_21114_, _01452_, \oc8051_golden_model_1.DPL [5]);
  and (_21115_, _21114_, _43223_);
  and (_43800_, _21115_, _21113_);
  and (_21117_, _11487_, \oc8051_golden_model_1.DPL [6]);
  nor (_21118_, _08106_, _11487_);
  or (_21119_, _21118_, _21117_);
  or (_21120_, _21119_, _07188_);
  and (_21121_, _15512_, _07932_);
  or (_21122_, _21121_, _21117_);
  or (_21123_, _21122_, _06252_);
  and (_21124_, _07932_, \oc8051_golden_model_1.ACC [6]);
  or (_21125_, _21124_, _21117_);
  and (_21126_, _21125_, _07123_);
  and (_21128_, _07124_, \oc8051_golden_model_1.DPL [6]);
  or (_21129_, _21128_, _06251_);
  or (_21130_, _21129_, _21126_);
  and (_21131_, _21130_, _07142_);
  and (_21132_, _21131_, _21123_);
  and (_21133_, _21119_, _06468_);
  or (_21134_, _21133_, _06466_);
  or (_21135_, _21134_, _21132_);
  or (_21136_, _21125_, _06801_);
  and (_21137_, _21136_, _11506_);
  and (_21139_, _21137_, _21135_);
  nor (_21140_, _11514_, \oc8051_golden_model_1.DPL [6]);
  nor (_21141_, _21140_, _11515_);
  and (_21142_, _21141_, _11505_);
  or (_21143_, _21142_, _21139_);
  and (_21144_, _21143_, _06370_);
  nor (_21145_, _08802_, _06370_);
  or (_21146_, _21145_, _07187_);
  or (_21147_, _21146_, _21144_);
  and (_21148_, _21147_, _21120_);
  or (_21150_, _21148_, _07182_);
  and (_21151_, _09067_, _07932_);
  or (_21152_, _21117_, _07183_);
  or (_21153_, _21152_, _21151_);
  and (_21154_, _21153_, _06336_);
  and (_21155_, _21154_, _21150_);
  and (_21156_, _15601_, _07932_);
  or (_21157_, _21156_, _21117_);
  and (_21158_, _21157_, _05968_);
  or (_21159_, _21158_, _06371_);
  or (_21161_, _21159_, _21155_);
  and (_21162_, _15608_, _07932_);
  or (_21163_, _21162_, _21117_);
  or (_21164_, _21163_, _07198_);
  and (_21165_, _21164_, _21161_);
  or (_21166_, _21165_, _06367_);
  and (_21167_, _15618_, _07932_);
  or (_21168_, _21167_, _21117_);
  or (_21169_, _21168_, _07218_);
  and (_21170_, _21169_, _07216_);
  and (_21172_, _21170_, _21166_);
  and (_21173_, _11202_, _07932_);
  or (_21174_, _21173_, _21117_);
  and (_21175_, _21174_, _06533_);
  or (_21176_, _21175_, _21172_);
  and (_21177_, _21176_, _07213_);
  or (_21178_, _21117_, _08109_);
  and (_21179_, _21163_, _06366_);
  and (_21180_, _21179_, _21178_);
  or (_21181_, _21180_, _21177_);
  and (_21183_, _21181_, _07210_);
  and (_21184_, _21125_, _06541_);
  and (_21185_, _21184_, _21178_);
  or (_21186_, _21185_, _06383_);
  or (_21187_, _21186_, _21183_);
  and (_21188_, _15615_, _07932_);
  or (_21189_, _21117_, _07231_);
  or (_21190_, _21189_, _21188_);
  and (_21191_, _21190_, _07229_);
  and (_21192_, _21191_, _21187_);
  nor (_21194_, _11201_, _11487_);
  or (_21195_, _21194_, _21117_);
  and (_21196_, _21195_, _06528_);
  or (_21197_, _21196_, _06563_);
  or (_21198_, _21197_, _21192_);
  or (_21199_, _21122_, _07241_);
  and (_21200_, _21199_, _06189_);
  and (_21201_, _21200_, _21198_);
  and (_21202_, _15676_, _07932_);
  or (_21203_, _21202_, _21117_);
  and (_21205_, _21203_, _06188_);
  or (_21206_, _21205_, _01456_);
  or (_21207_, _21206_, _21201_);
  or (_21208_, _01452_, \oc8051_golden_model_1.DPL [6]);
  and (_21209_, _21208_, _43223_);
  and (_43801_, _21209_, _21207_);
  nor (_21210_, _01452_, _12637_);
  nor (_21211_, _07935_, _12637_);
  and (_21212_, _07935_, \oc8051_golden_model_1.ACC [0]);
  and (_21213_, _21212_, _08351_);
  or (_21215_, _21213_, _21211_);
  or (_21216_, _21215_, _07210_);
  and (_21217_, _09342_, _07935_);
  or (_21218_, _21217_, _21211_);
  and (_21219_, _21218_, _07182_);
  nor (_21220_, _11517_, \oc8051_golden_model_1.DPH [0]);
  nor (_21221_, _21220_, _11604_);
  and (_21222_, _21221_, _11505_);
  and (_21223_, _08151_, _07325_);
  or (_21224_, _21223_, _21211_);
  or (_21226_, _21224_, _07142_);
  nor (_21227_, _08351_, _11583_);
  or (_21228_, _21227_, _21211_);
  and (_21229_, _21228_, _06251_);
  nor (_21230_, _07123_, _12637_);
  or (_21231_, _21212_, _21211_);
  and (_21232_, _21231_, _07123_);
  or (_21233_, _21232_, _21230_);
  and (_21234_, _21233_, _06252_);
  or (_21235_, _21234_, _06468_);
  or (_21237_, _21235_, _21229_);
  and (_21238_, _21237_, _21226_);
  or (_21239_, _21238_, _06466_);
  or (_21240_, _21231_, _06801_);
  and (_21241_, _21240_, _11506_);
  and (_21242_, _21241_, _21239_);
  or (_21243_, _21242_, _21222_);
  and (_21244_, _21243_, _06370_);
  and (_21245_, _06799_, _06369_);
  or (_21246_, _21245_, _07187_);
  or (_21248_, _21246_, _21244_);
  or (_21249_, _21224_, _07188_);
  and (_21250_, _21249_, _07183_);
  and (_21251_, _21250_, _21248_);
  or (_21252_, _21251_, _05968_);
  or (_21253_, _21252_, _21219_);
  and (_21254_, _14427_, _08151_);
  or (_21255_, _21211_, _06336_);
  or (_21256_, _21255_, _21254_);
  and (_21257_, _21256_, _07198_);
  and (_21259_, _21257_, _21253_);
  and (_21260_, _07935_, _08908_);
  or (_21261_, _21260_, _21211_);
  and (_21262_, _21261_, _06371_);
  or (_21263_, _21262_, _06367_);
  or (_21264_, _21263_, _21259_);
  and (_21265_, _14442_, _07935_);
  or (_21266_, _21265_, _21211_);
  or (_21267_, _21266_, _07218_);
  and (_21268_, _21267_, _07216_);
  and (_21270_, _21268_, _21264_);
  nor (_21271_, _12526_, _11583_);
  or (_21272_, _21271_, _21211_);
  nor (_21273_, _21213_, _07216_);
  and (_21274_, _21273_, _21272_);
  or (_21275_, _21274_, _21270_);
  and (_21276_, _21275_, _07213_);
  nand (_21277_, _21261_, _06366_);
  nor (_21278_, _21277_, _21227_);
  or (_21279_, _21278_, _06541_);
  or (_21281_, _21279_, _21276_);
  and (_21282_, _21281_, _21216_);
  or (_21283_, _21282_, _06383_);
  and (_21284_, _14325_, _07935_);
  or (_21285_, _21284_, _21211_);
  or (_21286_, _21285_, _07231_);
  and (_21287_, _21286_, _07229_);
  and (_21288_, _21287_, _21283_);
  and (_21289_, _21272_, _06528_);
  or (_21290_, _21289_, _19442_);
  or (_21291_, _21290_, _21288_);
  or (_21292_, _21228_, _06756_);
  and (_21293_, _21292_, _01452_);
  and (_21294_, _21293_, _21291_);
  or (_21295_, _21294_, _21210_);
  and (_43803_, _21295_, _43223_);
  not (_21296_, \oc8051_golden_model_1.DPH [1]);
  nor (_21297_, _07935_, _21296_);
  nor (_21298_, _11216_, _11583_);
  or (_21299_, _21298_, _21297_);
  or (_21302_, _21299_, _07229_);
  or (_21303_, _07935_, \oc8051_golden_model_1.DPH [1]);
  and (_21304_, _21303_, _06371_);
  nand (_21305_, _08151_, _07018_);
  and (_21306_, _21305_, _21304_);
  or (_21307_, _09297_, _11583_);
  and (_21308_, _21303_, _07182_);
  and (_21309_, _21308_, _21307_);
  nor (_21310_, _11604_, \oc8051_golden_model_1.DPH [1]);
  nor (_21311_, _21310_, _11605_);
  and (_21313_, _21311_, _11505_);
  and (_21314_, _14503_, _08151_);
  not (_21315_, _21314_);
  and (_21316_, _21315_, _21303_);
  or (_21317_, _21316_, _06252_);
  and (_21318_, _07935_, \oc8051_golden_model_1.ACC [1]);
  or (_21319_, _21318_, _21297_);
  and (_21320_, _21319_, _07123_);
  nor (_21321_, _07123_, _21296_);
  or (_21322_, _21321_, _06251_);
  or (_21324_, _21322_, _21320_);
  and (_21325_, _21324_, _07142_);
  and (_21326_, _21325_, _21317_);
  nor (_21327_, _11583_, _07120_);
  or (_21328_, _21327_, _21297_);
  and (_21329_, _21328_, _06468_);
  or (_21330_, _21329_, _06466_);
  or (_21331_, _21330_, _21326_);
  or (_21332_, _21319_, _06801_);
  and (_21333_, _21332_, _11506_);
  and (_21335_, _21333_, _21331_);
  or (_21336_, _21335_, _21313_);
  and (_21337_, _21336_, _06370_);
  nor (_21338_, _06155_, _06370_);
  or (_21339_, _21338_, _07187_);
  or (_21340_, _21339_, _21337_);
  or (_21341_, _21328_, _07188_);
  and (_21342_, _21341_, _07183_);
  and (_21343_, _21342_, _21340_);
  or (_21344_, _21343_, _21309_);
  and (_21346_, _21344_, _06336_);
  and (_21347_, _14609_, _07935_);
  or (_21348_, _21347_, _21297_);
  and (_21349_, _21348_, _05968_);
  or (_21350_, _21349_, _21346_);
  and (_21351_, _21350_, _07198_);
  or (_21352_, _21351_, _21306_);
  and (_21353_, _21352_, _07218_);
  or (_21354_, _14625_, _11583_);
  and (_21355_, _21303_, _06367_);
  and (_21357_, _21355_, _21354_);
  or (_21358_, _21357_, _06533_);
  or (_21359_, _21358_, _21353_);
  nand (_21360_, _11215_, _08151_);
  and (_21361_, _21360_, _21299_);
  or (_21362_, _21361_, _07216_);
  and (_21363_, _21362_, _07213_);
  and (_21364_, _21363_, _21359_);
  or (_21365_, _14623_, _11583_);
  and (_21366_, _21303_, _06366_);
  and (_21368_, _21366_, _21365_);
  or (_21369_, _21368_, _06541_);
  or (_21370_, _21369_, _21364_);
  nor (_21371_, _21297_, _07210_);
  nand (_21372_, _21371_, _21360_);
  and (_21373_, _21372_, _07231_);
  and (_21374_, _21373_, _21370_);
  or (_21375_, _21305_, _08302_);
  and (_21376_, _21303_, _06383_);
  and (_21377_, _21376_, _21375_);
  or (_21379_, _21377_, _06528_);
  or (_21380_, _21379_, _21374_);
  and (_21381_, _21380_, _21302_);
  or (_21382_, _21381_, _06563_);
  or (_21383_, _21316_, _07241_);
  and (_21384_, _21383_, _06189_);
  and (_21385_, _21384_, _21382_);
  or (_21386_, _21314_, _21297_);
  and (_21387_, _21386_, _06188_);
  or (_21388_, _21387_, _01456_);
  or (_21390_, _21388_, _21385_);
  or (_21391_, _01452_, \oc8051_golden_model_1.DPH [1]);
  and (_21392_, _21391_, _43223_);
  and (_43804_, _21392_, _21390_);
  and (_21393_, _01456_, \oc8051_golden_model_1.DPH [2]);
  and (_21394_, _11583_, \oc8051_golden_model_1.DPH [2]);
  nor (_21395_, _11583_, _07578_);
  or (_21396_, _21395_, _21394_);
  or (_21397_, _21396_, _07188_);
  or (_21398_, _11605_, \oc8051_golden_model_1.DPH [2]);
  nor (_21400_, _11606_, _11506_);
  and (_21401_, _21400_, _21398_);
  and (_21402_, _14712_, _08151_);
  or (_21403_, _21402_, _21394_);
  or (_21404_, _21403_, _06252_);
  and (_21405_, _07935_, \oc8051_golden_model_1.ACC [2]);
  or (_21406_, _21405_, _21394_);
  and (_21407_, _21406_, _07123_);
  and (_21408_, _07124_, \oc8051_golden_model_1.DPH [2]);
  or (_21409_, _21408_, _06251_);
  or (_21411_, _21409_, _21407_);
  and (_21412_, _21411_, _07142_);
  and (_21413_, _21412_, _21404_);
  and (_21414_, _21396_, _06468_);
  or (_21415_, _21414_, _06466_);
  or (_21416_, _21415_, _21413_);
  or (_21417_, _21406_, _06801_);
  and (_21418_, _21417_, _11506_);
  and (_21419_, _21418_, _21416_);
  or (_21420_, _21419_, _21401_);
  and (_21422_, _21420_, _06370_);
  nor (_21423_, _06750_, _06370_);
  or (_21424_, _21423_, _07187_);
  or (_21425_, _21424_, _21422_);
  and (_21426_, _21425_, _21397_);
  or (_21427_, _21426_, _07182_);
  or (_21428_, _21394_, _07183_);
  and (_21429_, _09251_, _07935_);
  or (_21430_, _21429_, _21428_);
  and (_21431_, _21430_, _06336_);
  and (_21433_, _21431_, _21427_);
  and (_21434_, _14808_, _07935_);
  or (_21435_, _21434_, _21394_);
  and (_21436_, _21435_, _05968_);
  or (_21437_, _21436_, _06371_);
  or (_21438_, _21437_, _21433_);
  and (_21439_, _07935_, _08945_);
  or (_21440_, _21439_, _21394_);
  or (_21441_, _21440_, _07198_);
  and (_21442_, _21441_, _21438_);
  or (_21444_, _21442_, _06367_);
  and (_21445_, _14824_, _07935_);
  or (_21446_, _21445_, _21394_);
  or (_21447_, _21446_, _07218_);
  and (_21448_, _21447_, _07216_);
  and (_21449_, _21448_, _21444_);
  and (_21450_, _11214_, _07935_);
  or (_21451_, _21450_, _21394_);
  and (_21452_, _21451_, _06533_);
  or (_21453_, _21452_, _21449_);
  and (_21455_, _21453_, _07213_);
  or (_21456_, _21394_, _08397_);
  and (_21457_, _21440_, _06366_);
  and (_21458_, _21457_, _21456_);
  or (_21459_, _21458_, _21455_);
  and (_21460_, _21459_, _07210_);
  and (_21461_, _21406_, _06541_);
  and (_21462_, _21461_, _21456_);
  or (_21463_, _21462_, _06383_);
  or (_21464_, _21463_, _21460_);
  and (_21466_, _14821_, _08151_);
  or (_21467_, _21394_, _07231_);
  or (_21468_, _21467_, _21466_);
  and (_21469_, _21468_, _07229_);
  and (_21470_, _21469_, _21464_);
  nor (_21471_, _11213_, _11583_);
  or (_21472_, _21471_, _21394_);
  and (_21473_, _21472_, _06528_);
  or (_21474_, _21473_, _21470_);
  and (_21475_, _21474_, _07241_);
  and (_21477_, _21403_, _06563_);
  or (_21478_, _21477_, _06188_);
  or (_21479_, _21478_, _21475_);
  and (_21480_, _14884_, _08151_);
  or (_21481_, _21394_, _06189_);
  or (_21482_, _21481_, _21480_);
  and (_21483_, _21482_, _01452_);
  and (_21484_, _21483_, _21479_);
  or (_21485_, _21484_, _21393_);
  and (_43805_, _21485_, _43223_);
  not (_21487_, \oc8051_golden_model_1.DPH [3]);
  nor (_21488_, _07935_, _21487_);
  nor (_21489_, _11583_, _07713_);
  or (_21490_, _21489_, _21488_);
  or (_21491_, _21490_, _07188_);
  or (_21492_, _11606_, \oc8051_golden_model_1.DPH [3]);
  nand (_21493_, _21492_, _11505_);
  nor (_21494_, _21493_, _11607_);
  and (_21495_, _14898_, _08151_);
  or (_21496_, _21495_, _21488_);
  or (_21498_, _21496_, _06252_);
  and (_21499_, _07935_, \oc8051_golden_model_1.ACC [3]);
  or (_21500_, _21499_, _21488_);
  and (_21501_, _21500_, _07123_);
  nor (_21502_, _07123_, _21487_);
  or (_21503_, _21502_, _06251_);
  or (_21504_, _21503_, _21501_);
  and (_21505_, _21504_, _07142_);
  and (_21506_, _21505_, _21498_);
  and (_21507_, _21490_, _06468_);
  or (_21509_, _21507_, _06466_);
  or (_21510_, _21509_, _21506_);
  or (_21511_, _21500_, _06801_);
  and (_21512_, _21511_, _11506_);
  and (_21513_, _21512_, _21510_);
  or (_21514_, _21513_, _21494_);
  and (_21515_, _21514_, _06370_);
  nor (_21516_, _06370_, _06292_);
  or (_21517_, _21516_, _07187_);
  or (_21518_, _21517_, _21515_);
  and (_21520_, _21518_, _21491_);
  or (_21521_, _21520_, _07182_);
  or (_21522_, _21488_, _07183_);
  and (_21523_, _09205_, _07935_);
  or (_21524_, _21523_, _21522_);
  and (_21525_, _21524_, _06336_);
  and (_21526_, _21525_, _21521_);
  and (_21527_, _15003_, _07935_);
  or (_21528_, _21527_, _21488_);
  and (_21529_, _21528_, _05968_);
  or (_21531_, _21529_, _06371_);
  or (_21532_, _21531_, _21526_);
  and (_21533_, _07935_, _08872_);
  or (_21534_, _21533_, _21488_);
  or (_21535_, _21534_, _07198_);
  and (_21536_, _21535_, _21532_);
  or (_21537_, _21536_, _06367_);
  and (_21538_, _15018_, _07935_);
  or (_21539_, _21538_, _21488_);
  or (_21540_, _21539_, _07218_);
  and (_21542_, _21540_, _07216_);
  and (_21543_, _21542_, _21537_);
  and (_21544_, _12523_, _07935_);
  or (_21545_, _21544_, _21488_);
  and (_21546_, _21545_, _06533_);
  or (_21547_, _21546_, _21543_);
  and (_21548_, _21547_, _07213_);
  or (_21549_, _21488_, _08257_);
  and (_21550_, _21534_, _06366_);
  and (_21551_, _21550_, _21549_);
  or (_21553_, _21551_, _21548_);
  and (_21554_, _21553_, _07210_);
  and (_21555_, _21500_, _06541_);
  and (_21556_, _21555_, _21549_);
  or (_21557_, _21556_, _06383_);
  or (_21558_, _21557_, _21554_);
  and (_21559_, _15015_, _08151_);
  or (_21560_, _21488_, _07231_);
  or (_21561_, _21560_, _21559_);
  and (_21562_, _21561_, _07229_);
  and (_21564_, _21562_, _21558_);
  nor (_21565_, _11211_, _11583_);
  or (_21566_, _21565_, _21488_);
  and (_21567_, _21566_, _06528_);
  or (_21568_, _21567_, _06563_);
  or (_21569_, _21568_, _21564_);
  or (_21570_, _21496_, _07241_);
  and (_21571_, _21570_, _06189_);
  and (_21572_, _21571_, _21569_);
  and (_21573_, _15075_, _08151_);
  or (_21575_, _21573_, _21488_);
  and (_21576_, _21575_, _06188_);
  or (_21577_, _21576_, _01456_);
  or (_21578_, _21577_, _21572_);
  or (_21579_, _01452_, \oc8051_golden_model_1.DPH [3]);
  and (_21580_, _21579_, _43223_);
  and (_43806_, _21580_, _21578_);
  not (_21581_, \oc8051_golden_model_1.DPH [4]);
  nor (_21582_, _07935_, _21581_);
  nor (_21583_, _08494_, _11583_);
  or (_21585_, _21583_, _21582_);
  or (_21586_, _21585_, _07188_);
  and (_21587_, _15108_, _08151_);
  or (_21588_, _21587_, _21582_);
  or (_21589_, _21588_, _06252_);
  and (_21590_, _07935_, \oc8051_golden_model_1.ACC [4]);
  or (_21591_, _21590_, _21582_);
  and (_21592_, _21591_, _07123_);
  nor (_21593_, _07123_, _21581_);
  or (_21594_, _21593_, _06251_);
  or (_21596_, _21594_, _21592_);
  and (_21597_, _21596_, _07142_);
  and (_21598_, _21597_, _21589_);
  and (_21599_, _21585_, _06468_);
  or (_21600_, _21599_, _06466_);
  or (_21601_, _21600_, _21598_);
  or (_21602_, _21591_, _06801_);
  and (_21603_, _21602_, _11506_);
  and (_21604_, _21603_, _21601_);
  or (_21605_, _11607_, \oc8051_golden_model_1.DPH [4]);
  nor (_21607_, _11608_, _11506_);
  and (_21608_, _21607_, _21605_);
  or (_21609_, _21608_, _21604_);
  and (_21610_, _21609_, _06370_);
  nor (_21611_, _06230_, _06370_);
  or (_21612_, _21611_, _07187_);
  or (_21613_, _21612_, _21610_);
  and (_21614_, _21613_, _21586_);
  or (_21615_, _21614_, _07182_);
  or (_21616_, _21582_, _07183_);
  and (_21618_, _09159_, _07935_);
  or (_21619_, _21618_, _21616_);
  and (_21620_, _21619_, _06336_);
  and (_21621_, _21620_, _21615_);
  and (_21622_, _15198_, _07935_);
  or (_21623_, _21622_, _21582_);
  and (_21624_, _21623_, _05968_);
  or (_21625_, _21624_, _06371_);
  or (_21626_, _21625_, _21621_);
  and (_21627_, _08892_, _07935_);
  or (_21629_, _21627_, _21582_);
  or (_21630_, _21629_, _07198_);
  and (_21631_, _21630_, _21626_);
  or (_21632_, _21631_, _06367_);
  and (_21633_, _15214_, _07935_);
  or (_21634_, _21633_, _21582_);
  or (_21635_, _21634_, _07218_);
  and (_21636_, _21635_, _07216_);
  and (_21637_, _21636_, _21632_);
  and (_21638_, _11209_, _07935_);
  or (_21639_, _21638_, _21582_);
  and (_21640_, _21639_, _06533_);
  or (_21641_, _21640_, _21637_);
  and (_21642_, _21641_, _07213_);
  or (_21643_, _21582_, _08497_);
  and (_21644_, _21629_, _06366_);
  and (_21645_, _21644_, _21643_);
  or (_21646_, _21645_, _21642_);
  and (_21647_, _21646_, _07210_);
  and (_21648_, _21591_, _06541_);
  and (_21651_, _21648_, _21643_);
  or (_21652_, _21651_, _06383_);
  or (_21653_, _21652_, _21647_);
  and (_21654_, _15211_, _08151_);
  or (_21655_, _21582_, _07231_);
  or (_21656_, _21655_, _21654_);
  and (_21657_, _21656_, _07229_);
  and (_21658_, _21657_, _21653_);
  nor (_21659_, _11208_, _11583_);
  or (_21660_, _21659_, _21582_);
  and (_21662_, _21660_, _06528_);
  or (_21663_, _21662_, _06563_);
  or (_21664_, _21663_, _21658_);
  or (_21665_, _21588_, _07241_);
  and (_21666_, _21665_, _06189_);
  and (_21667_, _21666_, _21664_);
  and (_21668_, _15280_, _08151_);
  or (_21669_, _21668_, _21582_);
  and (_21670_, _21669_, _06188_);
  or (_21671_, _21670_, _01456_);
  or (_21673_, _21671_, _21667_);
  or (_21674_, _01452_, \oc8051_golden_model_1.DPH [4]);
  and (_21675_, _21674_, _43223_);
  and (_43807_, _21675_, _21673_);
  and (_21676_, _11583_, \oc8051_golden_model_1.DPH [5]);
  nor (_21677_, _08209_, _11583_);
  or (_21678_, _21677_, _21676_);
  or (_21679_, _21678_, _07188_);
  and (_21680_, _15311_, _08151_);
  or (_21681_, _21680_, _21676_);
  or (_21683_, _21681_, _06252_);
  and (_21684_, _07935_, \oc8051_golden_model_1.ACC [5]);
  or (_21685_, _21684_, _21676_);
  and (_21686_, _21685_, _07123_);
  and (_21687_, _07124_, \oc8051_golden_model_1.DPH [5]);
  or (_21688_, _21687_, _06251_);
  or (_21689_, _21688_, _21686_);
  and (_21690_, _21689_, _07142_);
  and (_21691_, _21690_, _21683_);
  and (_21692_, _21678_, _06468_);
  or (_21694_, _21692_, _06466_);
  or (_21695_, _21694_, _21691_);
  or (_21696_, _21685_, _06801_);
  and (_21697_, _21696_, _11506_);
  and (_21698_, _21697_, _21695_);
  or (_21699_, _11608_, \oc8051_golden_model_1.DPH [5]);
  nor (_21700_, _11609_, _11506_);
  and (_21701_, _21700_, _21699_);
  or (_21702_, _21701_, _21698_);
  and (_21703_, _21702_, _06370_);
  nor (_21705_, _06608_, _06370_);
  or (_21706_, _21705_, _07187_);
  or (_21707_, _21706_, _21703_);
  and (_21708_, _21707_, _21679_);
  or (_21709_, _21708_, _07182_);
  or (_21710_, _21676_, _07183_);
  and (_21711_, _09113_, _07935_);
  or (_21712_, _21711_, _21710_);
  and (_21713_, _21712_, _06336_);
  and (_21714_, _21713_, _21709_);
  and (_21716_, _15400_, _07935_);
  or (_21717_, _21716_, _21676_);
  and (_21718_, _21717_, _05968_);
  or (_21719_, _21718_, _06371_);
  or (_21720_, _21719_, _21714_);
  and (_21721_, _08888_, _07935_);
  or (_21722_, _21721_, _21676_);
  or (_21723_, _21722_, _07198_);
  and (_21724_, _21723_, _21720_);
  or (_21725_, _21724_, _06367_);
  and (_21727_, _15416_, _07935_);
  or (_21728_, _21727_, _21676_);
  or (_21729_, _21728_, _07218_);
  and (_21730_, _21729_, _07216_);
  and (_21731_, _21730_, _21725_);
  and (_21732_, _11205_, _07935_);
  or (_21733_, _21732_, _21676_);
  and (_21734_, _21733_, _06533_);
  or (_21735_, _21734_, _21731_);
  and (_21736_, _21735_, _07213_);
  or (_21738_, _21676_, _08212_);
  and (_21739_, _21722_, _06366_);
  and (_21740_, _21739_, _21738_);
  or (_21741_, _21740_, _21736_);
  and (_21742_, _21741_, _07210_);
  and (_21743_, _21685_, _06541_);
  and (_21744_, _21743_, _21738_);
  or (_21745_, _21744_, _06383_);
  or (_21746_, _21745_, _21742_);
  and (_21747_, _15413_, _08151_);
  or (_21748_, _21676_, _07231_);
  or (_21749_, _21748_, _21747_);
  and (_21750_, _21749_, _07229_);
  and (_21751_, _21750_, _21746_);
  nor (_21752_, _11204_, _11583_);
  or (_21753_, _21752_, _21676_);
  and (_21754_, _21753_, _06528_);
  or (_21755_, _21754_, _06563_);
  or (_21756_, _21755_, _21751_);
  or (_21757_, _21681_, _07241_);
  and (_21760_, _21757_, _06189_);
  and (_21761_, _21760_, _21756_);
  and (_21762_, _15477_, _08151_);
  or (_21763_, _21762_, _21676_);
  and (_21764_, _21763_, _06188_);
  or (_21765_, _21764_, _01456_);
  or (_21766_, _21765_, _21761_);
  or (_21767_, _01452_, \oc8051_golden_model_1.DPH [5]);
  and (_21768_, _21767_, _43223_);
  and (_43809_, _21768_, _21766_);
  and (_21770_, _11583_, \oc8051_golden_model_1.DPH [6]);
  nor (_21771_, _08106_, _11583_);
  or (_21772_, _21771_, _21770_);
  or (_21773_, _21772_, _07188_);
  and (_21774_, _15512_, _08151_);
  or (_21775_, _21774_, _21770_);
  or (_21776_, _21775_, _06252_);
  and (_21777_, _07935_, \oc8051_golden_model_1.ACC [6]);
  or (_21778_, _21777_, _21770_);
  and (_21779_, _21778_, _07123_);
  and (_21781_, _07124_, \oc8051_golden_model_1.DPH [6]);
  or (_21782_, _21781_, _06251_);
  or (_21783_, _21782_, _21779_);
  and (_21784_, _21783_, _07142_);
  and (_21785_, _21784_, _21776_);
  and (_21786_, _21772_, _06468_);
  or (_21787_, _21786_, _06466_);
  or (_21788_, _21787_, _21785_);
  or (_21789_, _21778_, _06801_);
  and (_21790_, _21789_, _11506_);
  and (_21792_, _21790_, _21788_);
  or (_21793_, _11609_, \oc8051_golden_model_1.DPH [6]);
  nor (_21794_, _11610_, _11506_);
  and (_21795_, _21794_, _21793_);
  or (_21796_, _21795_, _21792_);
  and (_21797_, _21796_, _06370_);
  nor (_21798_, _06370_, _06326_);
  or (_21799_, _21798_, _07187_);
  or (_21800_, _21799_, _21797_);
  and (_21801_, _21800_, _21773_);
  or (_21803_, _21801_, _07182_);
  or (_21804_, _21770_, _07183_);
  and (_21805_, _09067_, _07935_);
  or (_21806_, _21805_, _21804_);
  and (_21807_, _21806_, _06336_);
  and (_21808_, _21807_, _21803_);
  and (_21809_, _15601_, _07935_);
  or (_21810_, _21809_, _21770_);
  and (_21811_, _21810_, _05968_);
  or (_21812_, _21811_, _06371_);
  or (_21814_, _21812_, _21808_);
  and (_21815_, _15608_, _07935_);
  or (_21816_, _21815_, _21770_);
  or (_21817_, _21816_, _07198_);
  and (_21818_, _21817_, _21814_);
  or (_21819_, _21818_, _06367_);
  and (_21820_, _15618_, _07935_);
  or (_21821_, _21820_, _21770_);
  or (_21822_, _21821_, _07218_);
  and (_21823_, _21822_, _07216_);
  and (_21825_, _21823_, _21819_);
  and (_21826_, _11202_, _07935_);
  or (_21827_, _21826_, _21770_);
  and (_21828_, _21827_, _06533_);
  or (_21829_, _21828_, _21825_);
  and (_21830_, _21829_, _07213_);
  or (_21831_, _21770_, _08109_);
  and (_21832_, _21816_, _06366_);
  and (_21833_, _21832_, _21831_);
  or (_21834_, _21833_, _21830_);
  and (_21836_, _21834_, _07210_);
  and (_21837_, _21778_, _06541_);
  and (_21838_, _21837_, _21831_);
  or (_21839_, _21838_, _06383_);
  or (_21840_, _21839_, _21836_);
  and (_21841_, _15615_, _08151_);
  or (_21842_, _21770_, _07231_);
  or (_21843_, _21842_, _21841_);
  and (_21844_, _21843_, _07229_);
  and (_21845_, _21844_, _21840_);
  nor (_21847_, _11201_, _11583_);
  or (_21848_, _21847_, _21770_);
  and (_21849_, _21848_, _06528_);
  or (_21850_, _21849_, _06563_);
  or (_21851_, _21850_, _21845_);
  or (_21852_, _21775_, _07241_);
  and (_21853_, _21852_, _06189_);
  and (_21854_, _21853_, _21851_);
  and (_21855_, _15676_, _08151_);
  or (_21856_, _21855_, _21770_);
  and (_21858_, _21856_, _06188_);
  or (_21859_, _21858_, _01456_);
  or (_21860_, _21859_, _21854_);
  or (_21861_, _01452_, \oc8051_golden_model_1.DPH [6]);
  and (_21862_, _21861_, _43223_);
  and (_43810_, _21862_, _21860_);
  not (_21863_, \oc8051_golden_model_1.TL1 [0]);
  nor (_21864_, _01452_, _21863_);
  nand (_21865_, _11218_, _07940_);
  nor (_21866_, _07940_, _21863_);
  nor (_21868_, _21866_, _07210_);
  nand (_21869_, _21868_, _21865_);
  and (_21870_, _07940_, _07325_);
  or (_21871_, _21870_, _21866_);
  or (_21872_, _21871_, _07188_);
  nor (_21873_, _08351_, _11673_);
  or (_21874_, _21873_, _21866_);
  or (_21875_, _21874_, _06252_);
  and (_21876_, _07940_, \oc8051_golden_model_1.ACC [0]);
  or (_21877_, _21876_, _21866_);
  and (_21879_, _21877_, _07123_);
  nor (_21880_, _07123_, _21863_);
  or (_21881_, _21880_, _06251_);
  or (_21882_, _21881_, _21879_);
  and (_21883_, _21882_, _07142_);
  and (_21884_, _21883_, _21875_);
  and (_21885_, _21871_, _06468_);
  or (_21886_, _21885_, _21884_);
  and (_21887_, _21886_, _06801_);
  and (_21888_, _21877_, _06466_);
  or (_21890_, _21888_, _07187_);
  or (_21891_, _21890_, _21887_);
  and (_21892_, _21891_, _21872_);
  or (_21893_, _21892_, _07182_);
  and (_21894_, _09342_, _07940_);
  or (_21895_, _21866_, _07183_);
  or (_21896_, _21895_, _21894_);
  and (_21897_, _21896_, _21893_);
  or (_21898_, _21897_, _05968_);
  and (_21899_, _14427_, _07940_);
  or (_21901_, _21866_, _06336_);
  or (_21902_, _21901_, _21899_);
  and (_21903_, _21902_, _07198_);
  and (_21904_, _21903_, _21898_);
  and (_21905_, _07940_, _08908_);
  or (_21906_, _21905_, _21866_);
  and (_21907_, _21906_, _06371_);
  or (_21908_, _21907_, _06367_);
  or (_21909_, _21908_, _21904_);
  and (_21910_, _14442_, _07940_);
  or (_21912_, _21910_, _21866_);
  or (_21913_, _21912_, _07218_);
  and (_21914_, _21913_, _07216_);
  and (_21915_, _21914_, _21909_);
  nor (_21916_, _12526_, _11673_);
  or (_21917_, _21916_, _21866_);
  and (_21918_, _21865_, _06533_);
  and (_21919_, _21918_, _21917_);
  or (_21920_, _21919_, _21915_);
  and (_21921_, _21920_, _07213_);
  nand (_21923_, _21906_, _06366_);
  nor (_21924_, _21923_, _21873_);
  or (_21925_, _21924_, _06541_);
  or (_21926_, _21925_, _21921_);
  and (_21927_, _21926_, _21869_);
  or (_21928_, _21927_, _06383_);
  and (_21929_, _14325_, _07940_);
  or (_21930_, _21929_, _21866_);
  or (_21931_, _21930_, _07231_);
  and (_21932_, _21931_, _07229_);
  and (_21934_, _21932_, _21928_);
  and (_21935_, _21917_, _06528_);
  or (_21936_, _21935_, _19442_);
  or (_21937_, _21936_, _21934_);
  or (_21938_, _21874_, _06756_);
  and (_21939_, _21938_, _01452_);
  and (_21940_, _21939_, _21937_);
  or (_21941_, _21940_, _21864_);
  and (_43811_, _21941_, _43223_);
  not (_21942_, \oc8051_golden_model_1.TL1 [1]);
  nor (_21944_, _07940_, _21942_);
  nor (_21945_, _11216_, _11673_);
  or (_21946_, _21945_, _21944_);
  or (_21947_, _21946_, _07229_);
  or (_21948_, _07940_, \oc8051_golden_model_1.TL1 [1]);
  and (_21949_, _14503_, _07940_);
  not (_21950_, _21949_);
  and (_21951_, _21950_, _21948_);
  or (_21952_, _21951_, _06252_);
  and (_21953_, _07940_, \oc8051_golden_model_1.ACC [1]);
  or (_21955_, _21953_, _21944_);
  and (_21956_, _21955_, _07123_);
  nor (_21957_, _07123_, _21942_);
  or (_21958_, _21957_, _06251_);
  or (_21959_, _21958_, _21956_);
  and (_21960_, _21959_, _07142_);
  and (_21961_, _21960_, _21952_);
  nor (_21962_, _11673_, _07120_);
  or (_21963_, _21962_, _21944_);
  and (_21964_, _21963_, _06468_);
  or (_21966_, _21964_, _21961_);
  and (_21967_, _21966_, _06801_);
  and (_21968_, _21955_, _06466_);
  or (_21969_, _21968_, _07187_);
  or (_21970_, _21969_, _21967_);
  or (_21971_, _21963_, _07188_);
  and (_21972_, _21971_, _07183_);
  and (_21973_, _21972_, _21970_);
  or (_21974_, _09297_, _11673_);
  and (_21975_, _21948_, _07182_);
  and (_21977_, _21975_, _21974_);
  or (_21978_, _21977_, _21973_);
  and (_21979_, _21978_, _06336_);
  or (_21980_, _14609_, _11673_);
  and (_21981_, _21948_, _05968_);
  and (_21982_, _21981_, _21980_);
  or (_21983_, _21982_, _21979_);
  and (_21984_, _21983_, _07198_);
  nand (_21985_, _07940_, _07018_);
  and (_21986_, _21948_, _06371_);
  and (_21988_, _21986_, _21985_);
  or (_21989_, _21988_, _21984_);
  and (_21990_, _21989_, _07218_);
  or (_21991_, _14625_, _11673_);
  and (_21992_, _21948_, _06367_);
  and (_21993_, _21992_, _21991_);
  or (_21994_, _21993_, _06533_);
  or (_21995_, _21994_, _21990_);
  nand (_21996_, _11215_, _07940_);
  and (_21997_, _21996_, _21946_);
  or (_21999_, _21997_, _07216_);
  and (_22000_, _21999_, _07213_);
  and (_22001_, _22000_, _21995_);
  or (_22002_, _14623_, _11673_);
  and (_22003_, _21948_, _06366_);
  and (_22004_, _22003_, _22002_);
  or (_22005_, _22004_, _06541_);
  or (_22006_, _22005_, _22001_);
  nor (_22007_, _21944_, _07210_);
  nand (_22008_, _22007_, _21996_);
  and (_22010_, _22008_, _07231_);
  and (_22011_, _22010_, _22006_);
  or (_22012_, _21985_, _08302_);
  and (_22013_, _21948_, _06383_);
  and (_22014_, _22013_, _22012_);
  or (_22015_, _22014_, _06528_);
  or (_22016_, _22015_, _22011_);
  and (_22017_, _22016_, _21947_);
  or (_22018_, _22017_, _06563_);
  or (_22019_, _21951_, _07241_);
  and (_22021_, _22019_, _06189_);
  and (_22022_, _22021_, _22018_);
  or (_22023_, _21949_, _21944_);
  and (_22024_, _22023_, _06188_);
  or (_22025_, _22024_, _01456_);
  or (_22026_, _22025_, _22022_);
  or (_22027_, _01452_, \oc8051_golden_model_1.TL1 [1]);
  and (_22028_, _22027_, _43223_);
  and (_43813_, _22028_, _22026_);
  not (_22029_, \oc8051_golden_model_1.TL1 [2]);
  nor (_22031_, _01452_, _22029_);
  nor (_22032_, _07940_, _22029_);
  and (_22033_, _09251_, _07940_);
  or (_22034_, _22033_, _22032_);
  and (_22035_, _22034_, _07182_);
  and (_22036_, _14712_, _07940_);
  or (_22037_, _22036_, _22032_);
  or (_22038_, _22037_, _06252_);
  and (_22039_, _07940_, \oc8051_golden_model_1.ACC [2]);
  or (_22040_, _22039_, _22032_);
  and (_22042_, _22040_, _07123_);
  nor (_22043_, _07123_, _22029_);
  or (_22044_, _22043_, _06251_);
  or (_22045_, _22044_, _22042_);
  and (_22046_, _22045_, _07142_);
  and (_22047_, _22046_, _22038_);
  nor (_22048_, _11673_, _07578_);
  or (_22049_, _22048_, _22032_);
  and (_22050_, _22049_, _06468_);
  or (_22051_, _22050_, _22047_);
  and (_22053_, _22051_, _06801_);
  and (_22054_, _22040_, _06466_);
  or (_22055_, _22054_, _07187_);
  or (_22056_, _22055_, _22053_);
  or (_22057_, _22049_, _07188_);
  and (_22058_, _22057_, _07183_);
  and (_22059_, _22058_, _22056_);
  or (_22060_, _22059_, _05968_);
  or (_22061_, _22060_, _22035_);
  and (_22062_, _14808_, _07940_);
  or (_22064_, _22032_, _06336_);
  or (_22065_, _22064_, _22062_);
  and (_22066_, _22065_, _07198_);
  and (_22067_, _22066_, _22061_);
  and (_22068_, _07940_, _08945_);
  or (_22069_, _22068_, _22032_);
  and (_22070_, _22069_, _06371_);
  or (_22071_, _22070_, _06367_);
  or (_22072_, _22071_, _22067_);
  and (_22073_, _14824_, _07940_);
  or (_22075_, _22073_, _22032_);
  or (_22076_, _22075_, _07218_);
  and (_22077_, _22076_, _07216_);
  and (_22078_, _22077_, _22072_);
  and (_22079_, _11214_, _07940_);
  or (_22080_, _22079_, _22032_);
  and (_22081_, _22080_, _06533_);
  or (_22082_, _22081_, _22078_);
  and (_22083_, _22082_, _07213_);
  or (_22084_, _22032_, _08397_);
  and (_22086_, _22069_, _06366_);
  and (_22087_, _22086_, _22084_);
  or (_22088_, _22087_, _22083_);
  and (_22089_, _22088_, _07210_);
  and (_22090_, _22040_, _06541_);
  and (_22091_, _22090_, _22084_);
  or (_22092_, _22091_, _06383_);
  or (_22093_, _22092_, _22089_);
  and (_22094_, _14821_, _07940_);
  or (_22095_, _22032_, _07231_);
  or (_22097_, _22095_, _22094_);
  and (_22098_, _22097_, _07229_);
  and (_22099_, _22098_, _22093_);
  nor (_22100_, _11213_, _11673_);
  or (_22101_, _22100_, _22032_);
  and (_22102_, _22101_, _06528_);
  or (_22103_, _22102_, _22099_);
  and (_22104_, _22103_, _07241_);
  and (_22105_, _22037_, _06563_);
  or (_22106_, _22105_, _06188_);
  or (_22109_, _22106_, _22104_);
  and (_22110_, _14884_, _07940_);
  or (_22111_, _22032_, _06189_);
  or (_22112_, _22111_, _22110_);
  and (_22113_, _22112_, _01452_);
  and (_22114_, _22113_, _22109_);
  or (_22115_, _22114_, _22031_);
  and (_43814_, _22115_, _43223_);
  and (_22116_, _11673_, \oc8051_golden_model_1.TL1 [3]);
  and (_22117_, _14898_, _07940_);
  or (_22119_, _22117_, _22116_);
  or (_22120_, _22119_, _06252_);
  and (_22121_, _07940_, \oc8051_golden_model_1.ACC [3]);
  or (_22122_, _22121_, _22116_);
  and (_22123_, _22122_, _07123_);
  and (_22124_, _07124_, \oc8051_golden_model_1.TL1 [3]);
  or (_22125_, _22124_, _06251_);
  or (_22126_, _22125_, _22123_);
  and (_22127_, _22126_, _07142_);
  and (_22128_, _22127_, _22120_);
  nor (_22130_, _11673_, _07713_);
  or (_22131_, _22130_, _22116_);
  and (_22132_, _22131_, _06468_);
  or (_22133_, _22132_, _22128_);
  and (_22134_, _22133_, _06801_);
  and (_22135_, _22122_, _06466_);
  or (_22136_, _22135_, _07187_);
  or (_22137_, _22136_, _22134_);
  or (_22138_, _22131_, _07188_);
  and (_22139_, _22138_, _07183_);
  and (_22141_, _22139_, _22137_);
  and (_22142_, _09205_, _07940_);
  or (_22143_, _22142_, _22116_);
  and (_22144_, _22143_, _07182_);
  or (_22145_, _22144_, _05968_);
  or (_22146_, _22145_, _22141_);
  and (_22147_, _15003_, _07940_);
  or (_22148_, _22116_, _06336_);
  or (_22149_, _22148_, _22147_);
  and (_22150_, _22149_, _07198_);
  and (_22152_, _22150_, _22146_);
  and (_22153_, _07940_, _08872_);
  or (_22154_, _22153_, _22116_);
  and (_22155_, _22154_, _06371_);
  or (_22156_, _22155_, _06367_);
  or (_22157_, _22156_, _22152_);
  and (_22158_, _15018_, _07940_);
  or (_22159_, _22158_, _22116_);
  or (_22160_, _22159_, _07218_);
  and (_22161_, _22160_, _07216_);
  and (_22163_, _22161_, _22157_);
  and (_22164_, _12523_, _07940_);
  or (_22165_, _22164_, _22116_);
  and (_22166_, _22165_, _06533_);
  or (_22167_, _22166_, _22163_);
  and (_22168_, _22167_, _07213_);
  or (_22169_, _22116_, _08257_);
  and (_22170_, _22154_, _06366_);
  and (_22171_, _22170_, _22169_);
  or (_22172_, _22171_, _22168_);
  and (_22174_, _22172_, _07210_);
  and (_22175_, _22122_, _06541_);
  and (_22176_, _22175_, _22169_);
  or (_22177_, _22176_, _06383_);
  or (_22178_, _22177_, _22174_);
  and (_22179_, _15015_, _07940_);
  or (_22180_, _22116_, _07231_);
  or (_22181_, _22180_, _22179_);
  and (_22182_, _22181_, _07229_);
  and (_22183_, _22182_, _22178_);
  nor (_22185_, _11211_, _11673_);
  or (_22186_, _22185_, _22116_);
  and (_22187_, _22186_, _06528_);
  or (_22188_, _22187_, _06563_);
  or (_22189_, _22188_, _22183_);
  or (_22190_, _22119_, _07241_);
  and (_22191_, _22190_, _06189_);
  and (_22192_, _22191_, _22189_);
  and (_22193_, _15075_, _07940_);
  or (_22194_, _22193_, _22116_);
  and (_22195_, _22194_, _06188_);
  or (_22196_, _22195_, _01456_);
  or (_22197_, _22196_, _22192_);
  or (_22198_, _01452_, \oc8051_golden_model_1.TL1 [3]);
  and (_22199_, _22198_, _43223_);
  and (_43815_, _22199_, _22197_);
  and (_22200_, _11673_, \oc8051_golden_model_1.TL1 [4]);
  nor (_22201_, _08494_, _11673_);
  or (_22202_, _22201_, _22200_);
  or (_22203_, _22202_, _07188_);
  and (_22206_, _15108_, _07940_);
  or (_22207_, _22206_, _22200_);
  or (_22208_, _22207_, _06252_);
  and (_22209_, _07940_, \oc8051_golden_model_1.ACC [4]);
  or (_22210_, _22209_, _22200_);
  and (_22211_, _22210_, _07123_);
  and (_22212_, _07124_, \oc8051_golden_model_1.TL1 [4]);
  or (_22213_, _22212_, _06251_);
  or (_22214_, _22213_, _22211_);
  and (_22215_, _22214_, _07142_);
  and (_22217_, _22215_, _22208_);
  and (_22218_, _22202_, _06468_);
  or (_22219_, _22218_, _22217_);
  and (_22220_, _22219_, _06801_);
  and (_22221_, _22210_, _06466_);
  or (_22222_, _22221_, _07187_);
  or (_22223_, _22222_, _22220_);
  and (_22224_, _22223_, _22203_);
  or (_22225_, _22224_, _07182_);
  and (_22226_, _09159_, _07940_);
  or (_22228_, _22200_, _07183_);
  or (_22229_, _22228_, _22226_);
  and (_22230_, _22229_, _22225_);
  or (_22231_, _22230_, _05968_);
  and (_22232_, _15198_, _07940_);
  or (_22233_, _22200_, _06336_);
  or (_22234_, _22233_, _22232_);
  and (_22235_, _22234_, _07198_);
  and (_22236_, _22235_, _22231_);
  and (_22237_, _08892_, _07940_);
  or (_22239_, _22237_, _22200_);
  and (_22240_, _22239_, _06371_);
  or (_22241_, _22240_, _06367_);
  or (_22242_, _22241_, _22236_);
  and (_22243_, _15214_, _07940_);
  or (_22244_, _22243_, _22200_);
  or (_22245_, _22244_, _07218_);
  and (_22246_, _22245_, _07216_);
  and (_22247_, _22246_, _22242_);
  and (_22248_, _11209_, _07940_);
  or (_22250_, _22248_, _22200_);
  and (_22251_, _22250_, _06533_);
  or (_22252_, _22251_, _22247_);
  and (_22253_, _22252_, _07213_);
  or (_22254_, _22200_, _08497_);
  and (_22255_, _22239_, _06366_);
  and (_22256_, _22255_, _22254_);
  or (_22257_, _22256_, _22253_);
  and (_22258_, _22257_, _07210_);
  and (_22259_, _22210_, _06541_);
  and (_22261_, _22259_, _22254_);
  or (_22262_, _22261_, _06383_);
  or (_22263_, _22262_, _22258_);
  and (_22264_, _15211_, _07940_);
  or (_22265_, _22200_, _07231_);
  or (_22266_, _22265_, _22264_);
  and (_22267_, _22266_, _07229_);
  and (_22268_, _22267_, _22263_);
  nor (_22269_, _11208_, _11673_);
  or (_22270_, _22269_, _22200_);
  and (_22272_, _22270_, _06528_);
  or (_22273_, _22272_, _06563_);
  or (_22274_, _22273_, _22268_);
  or (_22275_, _22207_, _07241_);
  and (_22276_, _22275_, _06189_);
  and (_22277_, _22276_, _22274_);
  and (_22278_, _15280_, _07940_);
  or (_22279_, _22278_, _22200_);
  and (_22280_, _22279_, _06188_);
  or (_22281_, _22280_, _01456_);
  or (_22283_, _22281_, _22277_);
  or (_22284_, _01452_, \oc8051_golden_model_1.TL1 [4]);
  and (_22285_, _22284_, _43223_);
  and (_43816_, _22285_, _22283_);
  and (_22286_, _11673_, \oc8051_golden_model_1.TL1 [5]);
  nor (_22287_, _08209_, _11673_);
  or (_22288_, _22287_, _22286_);
  or (_22289_, _22288_, _07188_);
  and (_22290_, _15311_, _07940_);
  or (_22291_, _22290_, _22286_);
  or (_22293_, _22291_, _06252_);
  and (_22294_, _07940_, \oc8051_golden_model_1.ACC [5]);
  or (_22295_, _22294_, _22286_);
  and (_22296_, _22295_, _07123_);
  and (_22297_, _07124_, \oc8051_golden_model_1.TL1 [5]);
  or (_22298_, _22297_, _06251_);
  or (_22299_, _22298_, _22296_);
  and (_22300_, _22299_, _07142_);
  and (_22301_, _22300_, _22293_);
  and (_22302_, _22288_, _06468_);
  or (_22304_, _22302_, _22301_);
  and (_22305_, _22304_, _06801_);
  and (_22306_, _22295_, _06466_);
  or (_22307_, _22306_, _07187_);
  or (_22308_, _22307_, _22305_);
  and (_22309_, _22308_, _22289_);
  or (_22310_, _22309_, _07182_);
  and (_22311_, _09113_, _07940_);
  or (_22312_, _22286_, _07183_);
  or (_22313_, _22312_, _22311_);
  and (_22315_, _22313_, _06336_);
  and (_22316_, _22315_, _22310_);
  and (_22317_, _15400_, _07940_);
  or (_22318_, _22317_, _22286_);
  and (_22319_, _22318_, _05968_);
  or (_22320_, _22319_, _06371_);
  or (_22321_, _22320_, _22316_);
  and (_22322_, _08888_, _07940_);
  or (_22323_, _22322_, _22286_);
  or (_22324_, _22323_, _07198_);
  and (_22326_, _22324_, _22321_);
  or (_22327_, _22326_, _06367_);
  and (_22328_, _15416_, _07940_);
  or (_22329_, _22328_, _22286_);
  or (_22330_, _22329_, _07218_);
  and (_22331_, _22330_, _07216_);
  and (_22332_, _22331_, _22327_);
  and (_22333_, _11205_, _07940_);
  or (_22334_, _22333_, _22286_);
  and (_22335_, _22334_, _06533_);
  or (_22337_, _22335_, _22332_);
  and (_22338_, _22337_, _07213_);
  or (_22339_, _22286_, _08212_);
  and (_22340_, _22323_, _06366_);
  and (_22341_, _22340_, _22339_);
  or (_22342_, _22341_, _22338_);
  and (_22343_, _22342_, _07210_);
  and (_22344_, _22295_, _06541_);
  and (_22345_, _22344_, _22339_);
  or (_22346_, _22345_, _06383_);
  or (_22348_, _22346_, _22343_);
  and (_22349_, _15413_, _07940_);
  or (_22350_, _22286_, _07231_);
  or (_22351_, _22350_, _22349_);
  and (_22352_, _22351_, _07229_);
  and (_22353_, _22352_, _22348_);
  nor (_22354_, _11204_, _11673_);
  or (_22355_, _22354_, _22286_);
  and (_22356_, _22355_, _06528_);
  or (_22357_, _22356_, _06563_);
  or (_22359_, _22357_, _22353_);
  or (_22360_, _22291_, _07241_);
  and (_22361_, _22360_, _06189_);
  and (_22362_, _22361_, _22359_);
  and (_22363_, _15477_, _07940_);
  or (_22364_, _22363_, _22286_);
  and (_22365_, _22364_, _06188_);
  or (_22366_, _22365_, _01456_);
  or (_22367_, _22366_, _22362_);
  or (_22368_, _01452_, \oc8051_golden_model_1.TL1 [5]);
  and (_22370_, _22368_, _43223_);
  and (_43817_, _22370_, _22367_);
  and (_22371_, _11673_, \oc8051_golden_model_1.TL1 [6]);
  and (_22372_, _15512_, _07940_);
  or (_22373_, _22372_, _22371_);
  or (_22374_, _22373_, _06252_);
  and (_22375_, _07940_, \oc8051_golden_model_1.ACC [6]);
  or (_22376_, _22375_, _22371_);
  and (_22377_, _22376_, _07123_);
  and (_22378_, _07124_, \oc8051_golden_model_1.TL1 [6]);
  or (_22380_, _22378_, _06251_);
  or (_22381_, _22380_, _22377_);
  and (_22382_, _22381_, _07142_);
  and (_22383_, _22382_, _22374_);
  nor (_22384_, _08106_, _11673_);
  or (_22385_, _22384_, _22371_);
  and (_22386_, _22385_, _06468_);
  or (_22387_, _22386_, _22383_);
  and (_22388_, _22387_, _06801_);
  and (_22389_, _22376_, _06466_);
  or (_22391_, _22389_, _07187_);
  or (_22392_, _22391_, _22388_);
  or (_22393_, _22385_, _07188_);
  and (_22394_, _22393_, _22392_);
  or (_22395_, _22394_, _07182_);
  and (_22396_, _09067_, _07940_);
  or (_22397_, _22371_, _07183_);
  or (_22398_, _22397_, _22396_);
  and (_22399_, _22398_, _06336_);
  and (_22400_, _22399_, _22395_);
  and (_22402_, _15601_, _07940_);
  or (_22403_, _22402_, _22371_);
  and (_22404_, _22403_, _05968_);
  or (_22405_, _22404_, _06371_);
  or (_22406_, _22405_, _22400_);
  and (_22407_, _15608_, _07940_);
  or (_22408_, _22407_, _22371_);
  or (_22409_, _22408_, _07198_);
  and (_22410_, _22409_, _22406_);
  or (_22411_, _22410_, _06367_);
  and (_22413_, _15618_, _07940_);
  or (_22414_, _22413_, _22371_);
  or (_22415_, _22414_, _07218_);
  and (_22416_, _22415_, _07216_);
  and (_22417_, _22416_, _22411_);
  and (_22418_, _11202_, _07940_);
  or (_22419_, _22418_, _22371_);
  and (_22420_, _22419_, _06533_);
  or (_22421_, _22420_, _22417_);
  and (_22422_, _22421_, _07213_);
  or (_22424_, _22371_, _08109_);
  and (_22425_, _22408_, _06366_);
  and (_22426_, _22425_, _22424_);
  or (_22427_, _22426_, _22422_);
  and (_22428_, _22427_, _07210_);
  and (_22429_, _22376_, _06541_);
  and (_22430_, _22429_, _22424_);
  or (_22431_, _22430_, _06383_);
  or (_22432_, _22431_, _22428_);
  and (_22433_, _15615_, _07940_);
  or (_22435_, _22371_, _07231_);
  or (_22436_, _22435_, _22433_);
  and (_22437_, _22436_, _07229_);
  and (_22438_, _22437_, _22432_);
  nor (_22439_, _11201_, _11673_);
  or (_22440_, _22439_, _22371_);
  and (_22441_, _22440_, _06528_);
  or (_22442_, _22441_, _06563_);
  or (_22443_, _22442_, _22438_);
  or (_22444_, _22373_, _07241_);
  and (_22446_, _22444_, _06189_);
  and (_22447_, _22446_, _22443_);
  and (_22448_, _15676_, _07940_);
  or (_22449_, _22448_, _22371_);
  and (_22450_, _22449_, _06188_);
  or (_22451_, _22450_, _01456_);
  or (_22452_, _22451_, _22447_);
  or (_22453_, _01452_, \oc8051_golden_model_1.TL1 [6]);
  and (_22454_, _22453_, _43223_);
  and (_43818_, _22454_, _22452_);
  and (_22456_, _01456_, \oc8051_golden_model_1.TL0 [0]);
  and (_22457_, _11751_, \oc8051_golden_model_1.TL0 [0]);
  and (_22458_, _07893_, \oc8051_golden_model_1.ACC [0]);
  and (_22459_, _22458_, _08351_);
  or (_22460_, _22459_, _22457_);
  or (_22461_, _22460_, _07210_);
  nor (_22462_, _08351_, _11767_);
  or (_22463_, _22462_, _22457_);
  or (_22464_, _22463_, _06252_);
  or (_22465_, _22458_, _22457_);
  and (_22467_, _22465_, _07123_);
  and (_22468_, _07124_, \oc8051_golden_model_1.TL0 [0]);
  or (_22469_, _22468_, _06251_);
  or (_22470_, _22469_, _22467_);
  and (_22471_, _22470_, _07142_);
  and (_22472_, _22471_, _22464_);
  and (_22473_, _08139_, _07325_);
  or (_22474_, _22473_, _22457_);
  and (_22475_, _22474_, _06468_);
  or (_22476_, _22475_, _22472_);
  and (_22478_, _22476_, _06801_);
  and (_22479_, _22465_, _06466_);
  or (_22480_, _22479_, _07187_);
  or (_22481_, _22480_, _22478_);
  or (_22482_, _22474_, _07188_);
  and (_22483_, _22482_, _22481_);
  or (_22484_, _22483_, _07182_);
  or (_22485_, _22457_, _07183_);
  and (_22486_, _09342_, _07893_);
  or (_22487_, _22486_, _22485_);
  and (_22488_, _22487_, _22484_);
  or (_22489_, _22488_, _05968_);
  and (_22490_, _14427_, _08139_);
  or (_22491_, _22457_, _06336_);
  or (_22492_, _22491_, _22490_);
  and (_22493_, _22492_, _07198_);
  and (_22494_, _22493_, _22489_);
  and (_22495_, _07893_, _08908_);
  or (_22496_, _22495_, _22457_);
  and (_22497_, _22496_, _06371_);
  or (_22500_, _22497_, _06367_);
  or (_22501_, _22500_, _22494_);
  and (_22502_, _14442_, _07893_);
  or (_22503_, _22502_, _22457_);
  or (_22504_, _22503_, _07218_);
  and (_22505_, _22504_, _07216_);
  and (_22506_, _22505_, _22501_);
  nor (_22507_, _12526_, _11767_);
  or (_22508_, _22507_, _22457_);
  nor (_22509_, _22459_, _07216_);
  and (_22511_, _22509_, _22508_);
  or (_22512_, _22511_, _22506_);
  and (_22513_, _22512_, _07213_);
  nand (_22514_, _22496_, _06366_);
  nor (_22515_, _22514_, _22462_);
  or (_22516_, _22515_, _06541_);
  or (_22517_, _22516_, _22513_);
  and (_22518_, _22517_, _22461_);
  or (_22519_, _22518_, _06383_);
  and (_22520_, _14325_, _08139_);
  or (_22522_, _22457_, _07231_);
  or (_22523_, _22522_, _22520_);
  and (_22524_, _22523_, _07229_);
  and (_22525_, _22524_, _22519_);
  and (_22526_, _22508_, _06528_);
  or (_22527_, _22526_, _19442_);
  or (_22528_, _22527_, _22525_);
  or (_22529_, _22463_, _06756_);
  and (_22530_, _22529_, _01452_);
  and (_22531_, _22530_, _22528_);
  or (_22533_, _22531_, _22456_);
  and (_43820_, _22533_, _43223_);
  and (_22534_, _01456_, \oc8051_golden_model_1.TL0 [1]);
  and (_22535_, _11751_, \oc8051_golden_model_1.TL0 [1]);
  or (_22536_, _22535_, _07183_);
  and (_22537_, _09297_, _07893_);
  or (_22538_, _22537_, _22536_);
  nor (_22539_, _11767_, _07120_);
  or (_22540_, _22535_, _19463_);
  or (_22541_, _22540_, _22539_);
  and (_22543_, _07893_, \oc8051_golden_model_1.ACC [1]);
  or (_22544_, _22543_, _22535_);
  and (_22545_, _22544_, _06466_);
  or (_22546_, _22545_, _07187_);
  or (_22547_, _07893_, \oc8051_golden_model_1.TL0 [1]);
  and (_22548_, _14503_, _08139_);
  not (_22549_, _22548_);
  and (_22550_, _22549_, _22547_);
  and (_22551_, _22550_, _06251_);
  and (_22552_, _07124_, \oc8051_golden_model_1.TL0 [1]);
  and (_22554_, _22544_, _07123_);
  or (_22555_, _22554_, _22552_);
  and (_22556_, _22555_, _06252_);
  or (_22557_, _22556_, _06468_);
  or (_22558_, _22557_, _22551_);
  and (_22559_, _22558_, _06801_);
  or (_22560_, _22559_, _22546_);
  and (_22561_, _22560_, _22541_);
  or (_22562_, _22561_, _07182_);
  and (_22563_, _22562_, _06336_);
  and (_22565_, _22563_, _22538_);
  and (_22566_, _14609_, _07893_);
  or (_22567_, _22566_, _22535_);
  and (_22568_, _22567_, _05968_);
  or (_22569_, _22568_, _22565_);
  and (_22570_, _22569_, _07198_);
  and (_22571_, _22547_, _06371_);
  nand (_22572_, _08139_, _07018_);
  and (_22573_, _22572_, _22571_);
  or (_22574_, _22573_, _22570_);
  and (_22576_, _22574_, _07218_);
  or (_22577_, _14625_, _11767_);
  and (_22578_, _22547_, _06367_);
  and (_22579_, _22578_, _22577_);
  or (_22580_, _22579_, _06533_);
  or (_22581_, _22580_, _22576_);
  nor (_22582_, _11216_, _11767_);
  or (_22583_, _22582_, _22535_);
  nand (_22584_, _11215_, _08139_);
  and (_22585_, _22584_, _22583_);
  or (_22587_, _22585_, _07216_);
  and (_22588_, _22587_, _07213_);
  and (_22589_, _22588_, _22581_);
  or (_22590_, _14623_, _11767_);
  and (_22591_, _22547_, _06366_);
  and (_22592_, _22591_, _22590_);
  or (_22593_, _22592_, _06541_);
  or (_22594_, _22593_, _22589_);
  nor (_22595_, _22535_, _07210_);
  nand (_22596_, _22595_, _22584_);
  and (_22597_, _22596_, _07231_);
  and (_22598_, _22597_, _22594_);
  or (_22599_, _22572_, _08302_);
  and (_22600_, _22547_, _06383_);
  and (_22601_, _22600_, _22599_);
  or (_22602_, _22601_, _06528_);
  or (_22603_, _22602_, _22598_);
  or (_22604_, _22583_, _07229_);
  and (_22605_, _22604_, _07241_);
  and (_22606_, _22605_, _22603_);
  and (_22609_, _22550_, _06563_);
  or (_22610_, _22609_, _06188_);
  or (_22611_, _22610_, _22606_);
  or (_22612_, _22535_, _06189_);
  or (_22613_, _22612_, _22548_);
  and (_22614_, _22613_, _01452_);
  and (_22615_, _22614_, _22611_);
  or (_22616_, _22615_, _22534_);
  and (_43821_, _22616_, _43223_);
  and (_22617_, _01456_, \oc8051_golden_model_1.TL0 [2]);
  and (_22619_, _11751_, \oc8051_golden_model_1.TL0 [2]);
  nor (_22620_, _11767_, _07578_);
  or (_22621_, _22620_, _22619_);
  or (_22622_, _22621_, _07188_);
  and (_22623_, _14712_, _08139_);
  or (_22624_, _22623_, _22619_);
  and (_22625_, _22624_, _06251_);
  and (_22626_, _07124_, \oc8051_golden_model_1.TL0 [2]);
  and (_22627_, _07893_, \oc8051_golden_model_1.ACC [2]);
  or (_22628_, _22627_, _22619_);
  and (_22630_, _22628_, _07123_);
  or (_22631_, _22630_, _22626_);
  and (_22632_, _22631_, _06252_);
  or (_22633_, _22632_, _06468_);
  or (_22634_, _22633_, _22625_);
  or (_22635_, _22621_, _07142_);
  and (_22636_, _22635_, _06801_);
  and (_22637_, _22636_, _22634_);
  and (_22638_, _22628_, _06466_);
  or (_22639_, _22638_, _07187_);
  or (_22641_, _22639_, _22637_);
  and (_22642_, _22641_, _22622_);
  or (_22643_, _22642_, _07182_);
  or (_22644_, _22619_, _07183_);
  and (_22645_, _09251_, _07893_);
  or (_22646_, _22645_, _22644_);
  and (_22647_, _22646_, _22643_);
  or (_22648_, _22647_, _05968_);
  and (_22649_, _14808_, _08139_);
  or (_22650_, _22619_, _06336_);
  or (_22652_, _22650_, _22649_);
  and (_22653_, _22652_, _07198_);
  and (_22654_, _22653_, _22648_);
  and (_22655_, _07893_, _08945_);
  or (_22656_, _22655_, _22619_);
  and (_22657_, _22656_, _06371_);
  or (_22658_, _22657_, _06367_);
  or (_22659_, _22658_, _22654_);
  and (_22660_, _14824_, _07893_);
  or (_22661_, _22660_, _22619_);
  or (_22663_, _22661_, _07218_);
  and (_22664_, _22663_, _07216_);
  and (_22665_, _22664_, _22659_);
  and (_22666_, _11214_, _07893_);
  or (_22667_, _22666_, _22619_);
  and (_22668_, _22667_, _06533_);
  or (_22669_, _22668_, _22665_);
  and (_22670_, _22669_, _07213_);
  or (_22671_, _22619_, _08397_);
  and (_22672_, _22656_, _06366_);
  and (_22674_, _22672_, _22671_);
  or (_22675_, _22674_, _22670_);
  and (_22676_, _22675_, _07210_);
  and (_22677_, _22628_, _06541_);
  and (_22678_, _22677_, _22671_);
  or (_22679_, _22678_, _06383_);
  or (_22680_, _22679_, _22676_);
  and (_22681_, _14821_, _08139_);
  or (_22682_, _22619_, _07231_);
  or (_22683_, _22682_, _22681_);
  and (_22685_, _22683_, _07229_);
  and (_22686_, _22685_, _22680_);
  nor (_22687_, _11213_, _11767_);
  or (_22688_, _22687_, _22619_);
  and (_22689_, _22688_, _06528_);
  or (_22690_, _22689_, _22686_);
  and (_22691_, _22690_, _07241_);
  and (_22692_, _22624_, _06563_);
  or (_22693_, _22692_, _06188_);
  or (_22694_, _22693_, _22691_);
  and (_22696_, _14884_, _08139_);
  or (_22697_, _22619_, _06189_);
  or (_22698_, _22697_, _22696_);
  and (_22699_, _22698_, _01452_);
  and (_22700_, _22699_, _22694_);
  or (_22701_, _22700_, _22617_);
  and (_43822_, _22701_, _43223_);
  and (_22702_, _11751_, \oc8051_golden_model_1.TL0 [3]);
  and (_22703_, _14898_, _08139_);
  or (_22704_, _22703_, _22702_);
  or (_22706_, _22704_, _06252_);
  and (_22707_, _07893_, \oc8051_golden_model_1.ACC [3]);
  or (_22708_, _22707_, _22702_);
  and (_22709_, _22708_, _07123_);
  and (_22710_, _07124_, \oc8051_golden_model_1.TL0 [3]);
  or (_22711_, _22710_, _06251_);
  or (_22712_, _22711_, _22709_);
  and (_22713_, _22712_, _07142_);
  and (_22714_, _22713_, _22706_);
  nor (_22715_, _11767_, _07713_);
  or (_22717_, _22715_, _22702_);
  and (_22718_, _22717_, _06468_);
  or (_22719_, _22718_, _22714_);
  and (_22720_, _22719_, _06801_);
  and (_22721_, _22708_, _06466_);
  or (_22722_, _22721_, _07187_);
  or (_22723_, _22722_, _22720_);
  or (_22724_, _22717_, _07188_);
  and (_22725_, _22724_, _22723_);
  or (_22726_, _22725_, _07182_);
  and (_22728_, _09205_, _07893_);
  or (_22729_, _22702_, _07183_);
  or (_22730_, _22729_, _22728_);
  and (_22731_, _22730_, _06336_);
  and (_22732_, _22731_, _22726_);
  and (_22733_, _15003_, _07893_);
  or (_22734_, _22733_, _22702_);
  and (_22735_, _22734_, _05968_);
  or (_22736_, _22735_, _06371_);
  or (_22737_, _22736_, _22732_);
  and (_22739_, _07893_, _08872_);
  or (_22740_, _22739_, _22702_);
  or (_22741_, _22740_, _07198_);
  and (_22742_, _22741_, _22737_);
  or (_22743_, _22742_, _06367_);
  and (_22744_, _15018_, _07893_);
  or (_22745_, _22744_, _22702_);
  or (_22746_, _22745_, _07218_);
  and (_22747_, _22746_, _07216_);
  and (_22748_, _22747_, _22743_);
  and (_22750_, _12523_, _07893_);
  or (_22751_, _22750_, _22702_);
  and (_22752_, _22751_, _06533_);
  or (_22753_, _22752_, _22748_);
  and (_22754_, _22753_, _07213_);
  or (_22755_, _22702_, _08257_);
  and (_22756_, _22740_, _06366_);
  and (_22757_, _22756_, _22755_);
  or (_22758_, _22757_, _22754_);
  and (_22759_, _22758_, _07210_);
  and (_22761_, _22708_, _06541_);
  and (_22762_, _22761_, _22755_);
  or (_22763_, _22762_, _06383_);
  or (_22764_, _22763_, _22759_);
  and (_22765_, _15015_, _08139_);
  or (_22766_, _22702_, _07231_);
  or (_22767_, _22766_, _22765_);
  and (_22768_, _22767_, _07229_);
  and (_22769_, _22768_, _22764_);
  nor (_22770_, _11211_, _11767_);
  or (_22772_, _22770_, _22702_);
  and (_22773_, _22772_, _06528_);
  or (_22774_, _22773_, _06563_);
  or (_22775_, _22774_, _22769_);
  or (_22776_, _22704_, _07241_);
  and (_22777_, _22776_, _06189_);
  and (_22778_, _22777_, _22775_);
  and (_22779_, _15075_, _08139_);
  or (_22780_, _22779_, _22702_);
  and (_22781_, _22780_, _06188_);
  or (_22783_, _22781_, _01456_);
  or (_22784_, _22783_, _22778_);
  or (_22785_, _01452_, \oc8051_golden_model_1.TL0 [3]);
  and (_22786_, _22785_, _43223_);
  and (_43823_, _22786_, _22784_);
  and (_22787_, _11751_, \oc8051_golden_model_1.TL0 [4]);
  nor (_22788_, _08494_, _11767_);
  or (_22789_, _22788_, _22787_);
  or (_22790_, _22789_, _07188_);
  and (_22791_, _15108_, _08139_);
  or (_22793_, _22791_, _22787_);
  or (_22794_, _22793_, _06252_);
  and (_22795_, _07893_, \oc8051_golden_model_1.ACC [4]);
  or (_22796_, _22795_, _22787_);
  and (_22797_, _22796_, _07123_);
  and (_22798_, _07124_, \oc8051_golden_model_1.TL0 [4]);
  or (_22799_, _22798_, _06251_);
  or (_22800_, _22799_, _22797_);
  and (_22801_, _22800_, _07142_);
  and (_22802_, _22801_, _22794_);
  and (_22804_, _22789_, _06468_);
  or (_22805_, _22804_, _22802_);
  and (_22806_, _22805_, _06801_);
  and (_22807_, _22796_, _06466_);
  or (_22808_, _22807_, _07187_);
  or (_22809_, _22808_, _22806_);
  and (_22810_, _22809_, _22790_);
  or (_22811_, _22810_, _07182_);
  or (_22812_, _22787_, _07183_);
  and (_22813_, _09159_, _07893_);
  or (_22814_, _22813_, _22812_);
  and (_22815_, _22814_, _22811_);
  or (_22816_, _22815_, _05968_);
  and (_22817_, _15198_, _08139_);
  or (_22818_, _22787_, _06336_);
  or (_22819_, _22818_, _22817_);
  and (_22820_, _22819_, _07198_);
  and (_22821_, _22820_, _22816_);
  and (_22822_, _08892_, _07893_);
  or (_22823_, _22822_, _22787_);
  and (_22826_, _22823_, _06371_);
  or (_22827_, _22826_, _06367_);
  or (_22828_, _22827_, _22821_);
  and (_22829_, _15214_, _07893_);
  or (_22830_, _22829_, _22787_);
  or (_22831_, _22830_, _07218_);
  and (_22832_, _22831_, _07216_);
  and (_22833_, _22832_, _22828_);
  and (_22834_, _11209_, _07893_);
  or (_22835_, _22834_, _22787_);
  and (_22837_, _22835_, _06533_);
  or (_22838_, _22837_, _22833_);
  and (_22839_, _22838_, _07213_);
  or (_22840_, _22787_, _08497_);
  and (_22841_, _22823_, _06366_);
  and (_22842_, _22841_, _22840_);
  or (_22843_, _22842_, _22839_);
  and (_22844_, _22843_, _07210_);
  and (_22845_, _22796_, _06541_);
  and (_22846_, _22845_, _22840_);
  or (_22848_, _22846_, _06383_);
  or (_22849_, _22848_, _22844_);
  and (_22850_, _15211_, _08139_);
  or (_22851_, _22787_, _07231_);
  or (_22852_, _22851_, _22850_);
  and (_22853_, _22852_, _07229_);
  and (_22854_, _22853_, _22849_);
  nor (_22855_, _11208_, _11767_);
  or (_22856_, _22855_, _22787_);
  and (_22857_, _22856_, _06528_);
  or (_22859_, _22857_, _06563_);
  or (_22860_, _22859_, _22854_);
  or (_22861_, _22793_, _07241_);
  and (_22862_, _22861_, _06189_);
  and (_22863_, _22862_, _22860_);
  and (_22864_, _15280_, _08139_);
  or (_22865_, _22864_, _22787_);
  and (_22866_, _22865_, _06188_);
  or (_22867_, _22866_, _01456_);
  or (_22868_, _22867_, _22863_);
  or (_22870_, _01452_, \oc8051_golden_model_1.TL0 [4]);
  and (_22871_, _22870_, _43223_);
  and (_43824_, _22871_, _22868_);
  and (_22872_, _11751_, \oc8051_golden_model_1.TL0 [5]);
  nor (_22873_, _08209_, _11767_);
  or (_22874_, _22873_, _22872_);
  or (_22875_, _22874_, _07188_);
  and (_22876_, _15311_, _08139_);
  or (_22877_, _22876_, _22872_);
  or (_22878_, _22877_, _06252_);
  and (_22880_, _07893_, \oc8051_golden_model_1.ACC [5]);
  or (_22881_, _22880_, _22872_);
  and (_22882_, _22881_, _07123_);
  and (_22883_, _07124_, \oc8051_golden_model_1.TL0 [5]);
  or (_22884_, _22883_, _06251_);
  or (_22885_, _22884_, _22882_);
  and (_22886_, _22885_, _07142_);
  and (_22887_, _22886_, _22878_);
  and (_22888_, _22874_, _06468_);
  or (_22889_, _22888_, _22887_);
  and (_22891_, _22889_, _06801_);
  and (_22892_, _22881_, _06466_);
  or (_22893_, _22892_, _07187_);
  or (_22894_, _22893_, _22891_);
  and (_22895_, _22894_, _22875_);
  or (_22896_, _22895_, _07182_);
  or (_22897_, _22872_, _07183_);
  and (_22898_, _09113_, _07893_);
  or (_22899_, _22898_, _22897_);
  and (_22900_, _22899_, _06336_);
  and (_22902_, _22900_, _22896_);
  and (_22903_, _15400_, _07893_);
  or (_22904_, _22903_, _22872_);
  and (_22905_, _22904_, _05968_);
  or (_22906_, _22905_, _06371_);
  or (_22907_, _22906_, _22902_);
  and (_22908_, _08888_, _07893_);
  or (_22909_, _22908_, _22872_);
  or (_22910_, _22909_, _07198_);
  and (_22911_, _22910_, _22907_);
  or (_22913_, _22911_, _06367_);
  and (_22914_, _15416_, _07893_);
  or (_22915_, _22914_, _22872_);
  or (_22916_, _22915_, _07218_);
  and (_22917_, _22916_, _07216_);
  and (_22918_, _22917_, _22913_);
  and (_22919_, _11205_, _07893_);
  or (_22920_, _22919_, _22872_);
  and (_22921_, _22920_, _06533_);
  or (_22922_, _22921_, _22918_);
  and (_22924_, _22922_, _07213_);
  or (_22925_, _22872_, _08212_);
  and (_22926_, _22909_, _06366_);
  and (_22927_, _22926_, _22925_);
  or (_22928_, _22927_, _22924_);
  and (_22929_, _22928_, _07210_);
  and (_22930_, _22881_, _06541_);
  and (_22931_, _22930_, _22925_);
  or (_22932_, _22931_, _06383_);
  or (_22933_, _22932_, _22929_);
  and (_22935_, _15413_, _08139_);
  or (_22936_, _22872_, _07231_);
  or (_22937_, _22936_, _22935_);
  and (_22938_, _22937_, _07229_);
  and (_22939_, _22938_, _22933_);
  nor (_22940_, _11204_, _11767_);
  or (_22941_, _22940_, _22872_);
  and (_22942_, _22941_, _06528_);
  or (_22943_, _22942_, _06563_);
  or (_22944_, _22943_, _22939_);
  or (_22946_, _22877_, _07241_);
  and (_22947_, _22946_, _06189_);
  and (_22948_, _22947_, _22944_);
  and (_22949_, _15477_, _08139_);
  or (_22950_, _22949_, _22872_);
  and (_22951_, _22950_, _06188_);
  or (_22952_, _22951_, _01456_);
  or (_22953_, _22952_, _22948_);
  or (_22954_, _01452_, \oc8051_golden_model_1.TL0 [5]);
  and (_22955_, _22954_, _43223_);
  and (_43825_, _22955_, _22953_);
  and (_22957_, _11751_, \oc8051_golden_model_1.TL0 [6]);
  nor (_22958_, _08106_, _11767_);
  or (_22959_, _22958_, _22957_);
  or (_22960_, _22959_, _07188_);
  and (_22961_, _15512_, _08139_);
  or (_22962_, _22961_, _22957_);
  or (_22963_, _22962_, _06252_);
  and (_22964_, _07893_, \oc8051_golden_model_1.ACC [6]);
  or (_22965_, _22964_, _22957_);
  and (_22967_, _22965_, _07123_);
  and (_22968_, _07124_, \oc8051_golden_model_1.TL0 [6]);
  or (_22969_, _22968_, _06251_);
  or (_22970_, _22969_, _22967_);
  and (_22971_, _22970_, _07142_);
  and (_22972_, _22971_, _22963_);
  and (_22973_, _22959_, _06468_);
  or (_22974_, _22973_, _22972_);
  and (_22975_, _22974_, _06801_);
  and (_22976_, _22965_, _06466_);
  or (_22978_, _22976_, _07187_);
  or (_22979_, _22978_, _22975_);
  and (_22980_, _22979_, _22960_);
  or (_22981_, _22980_, _07182_);
  or (_22982_, _22957_, _07183_);
  and (_22983_, _09067_, _07893_);
  or (_22984_, _22983_, _22982_);
  and (_22985_, _22984_, _06336_);
  and (_22986_, _22985_, _22981_);
  and (_22987_, _15601_, _07893_);
  or (_22989_, _22987_, _22957_);
  and (_22990_, _22989_, _05968_);
  or (_22991_, _22990_, _06371_);
  or (_22992_, _22991_, _22986_);
  and (_22993_, _15608_, _07893_);
  or (_22994_, _22993_, _22957_);
  or (_22995_, _22994_, _07198_);
  and (_22996_, _22995_, _22992_);
  or (_22997_, _22996_, _06367_);
  and (_22998_, _15618_, _07893_);
  or (_23000_, _22998_, _22957_);
  or (_23001_, _23000_, _07218_);
  and (_23002_, _23001_, _07216_);
  and (_23003_, _23002_, _22997_);
  and (_23004_, _11202_, _07893_);
  or (_23005_, _23004_, _22957_);
  and (_23006_, _23005_, _06533_);
  or (_23007_, _23006_, _23003_);
  and (_23008_, _23007_, _07213_);
  or (_23009_, _22957_, _08109_);
  and (_23011_, _22994_, _06366_);
  and (_23012_, _23011_, _23009_);
  or (_23013_, _23012_, _23008_);
  and (_23014_, _23013_, _07210_);
  and (_23015_, _22965_, _06541_);
  and (_23016_, _23015_, _23009_);
  or (_23017_, _23016_, _06383_);
  or (_23018_, _23017_, _23014_);
  and (_23019_, _15615_, _08139_);
  or (_23020_, _22957_, _07231_);
  or (_23022_, _23020_, _23019_);
  and (_23023_, _23022_, _07229_);
  and (_23024_, _23023_, _23018_);
  nor (_23025_, _11201_, _11767_);
  or (_23026_, _23025_, _22957_);
  and (_23027_, _23026_, _06528_);
  or (_23028_, _23027_, _06563_);
  or (_23029_, _23028_, _23024_);
  or (_23030_, _22962_, _07241_);
  and (_23031_, _23030_, _06189_);
  and (_23033_, _23031_, _23029_);
  and (_23034_, _15676_, _08139_);
  or (_23035_, _23034_, _22957_);
  and (_23036_, _23035_, _06188_);
  or (_23037_, _23036_, _01456_);
  or (_23038_, _23037_, _23033_);
  or (_23039_, _01452_, \oc8051_golden_model_1.TL0 [6]);
  and (_23040_, _23039_, _43223_);
  and (_43826_, _23040_, _23038_);
  not (_23041_, \oc8051_golden_model_1.TCON [0]);
  nor (_23043_, _01452_, _23041_);
  nand (_23044_, _11218_, _07897_);
  nor (_23045_, _07897_, _23041_);
  nor (_23046_, _23045_, _07210_);
  nand (_23047_, _23046_, _23044_);
  and (_23048_, _07897_, _07325_);
  or (_23049_, _23048_, _23045_);
  or (_23050_, _23049_, _07188_);
  nor (_23051_, _08351_, _11831_);
  or (_23052_, _23051_, _23045_);
  and (_23054_, _23052_, _06251_);
  nor (_23055_, _07123_, _23041_);
  and (_23056_, _07897_, \oc8051_golden_model_1.ACC [0]);
  or (_23057_, _23056_, _23045_);
  and (_23058_, _23057_, _07123_);
  or (_23059_, _23058_, _23055_);
  and (_23060_, _23059_, _06252_);
  or (_23061_, _23060_, _06475_);
  or (_23062_, _23061_, _23054_);
  and (_23063_, _14341_, _08528_);
  nor (_23065_, _08528_, _23041_);
  or (_23066_, _23065_, _06476_);
  or (_23067_, _23066_, _23063_);
  and (_23068_, _23067_, _07142_);
  and (_23069_, _23068_, _23062_);
  and (_23070_, _23049_, _06468_);
  or (_23071_, _23070_, _06466_);
  or (_23072_, _23071_, _23069_);
  or (_23073_, _23057_, _06801_);
  and (_23074_, _23073_, _06484_);
  and (_23075_, _23074_, _23072_);
  and (_23076_, _23045_, _06483_);
  or (_23077_, _23076_, _06461_);
  or (_23078_, _23077_, _23075_);
  or (_23079_, _23052_, _07164_);
  and (_23080_, _23079_, _06242_);
  and (_23081_, _23080_, _23078_);
  and (_23082_, _14372_, _08528_);
  or (_23083_, _23082_, _23065_);
  and (_23084_, _23083_, _06241_);
  or (_23087_, _23084_, _07187_);
  or (_23088_, _23087_, _23081_);
  and (_23089_, _23088_, _23050_);
  or (_23090_, _23089_, _07182_);
  and (_23091_, _09342_, _07897_);
  or (_23092_, _23045_, _07183_);
  or (_23093_, _23092_, _23091_);
  and (_23094_, _23093_, _23090_);
  or (_23095_, _23094_, _05968_);
  and (_23096_, _14427_, _07897_);
  or (_23098_, _23045_, _06336_);
  or (_23099_, _23098_, _23096_);
  and (_23100_, _23099_, _07198_);
  and (_23101_, _23100_, _23095_);
  and (_23102_, _07897_, _08908_);
  or (_23103_, _23102_, _23045_);
  and (_23104_, _23103_, _06371_);
  or (_23105_, _23104_, _06367_);
  or (_23106_, _23105_, _23101_);
  and (_23107_, _14442_, _07897_);
  or (_23109_, _23107_, _23045_);
  or (_23110_, _23109_, _07218_);
  and (_23111_, _23110_, _07216_);
  and (_23112_, _23111_, _23106_);
  nor (_23113_, _12526_, _11831_);
  or (_23114_, _23113_, _23045_);
  and (_23115_, _23044_, _06533_);
  and (_23116_, _23115_, _23114_);
  or (_23117_, _23116_, _23112_);
  and (_23118_, _23117_, _07213_);
  nand (_23120_, _23103_, _06366_);
  nor (_23121_, _23120_, _23051_);
  or (_23122_, _23121_, _06541_);
  or (_23123_, _23122_, _23118_);
  and (_23124_, _23123_, _23047_);
  or (_23125_, _23124_, _06383_);
  and (_23126_, _14325_, _07897_);
  or (_23127_, _23045_, _07231_);
  or (_23128_, _23127_, _23126_);
  and (_23129_, _23128_, _07229_);
  and (_23131_, _23129_, _23125_);
  and (_23132_, _23114_, _06528_);
  or (_23133_, _23132_, _06563_);
  or (_23134_, _23133_, _23131_);
  or (_23135_, _23052_, _07241_);
  and (_23136_, _23135_, _23134_);
  or (_23137_, _23136_, _06199_);
  or (_23138_, _23045_, _06571_);
  and (_23139_, _23138_, _23137_);
  or (_23140_, _23139_, _06188_);
  or (_23142_, _23052_, _06189_);
  and (_23143_, _23142_, _01452_);
  and (_23144_, _23143_, _23140_);
  or (_23145_, _23144_, _23043_);
  and (_43828_, _23145_, _43223_);
  not (_23146_, \oc8051_golden_model_1.TCON [1]);
  nor (_23147_, _01452_, _23146_);
  nor (_23148_, _07897_, _23146_);
  nor (_23149_, _11216_, _11831_);
  or (_23150_, _23149_, _23148_);
  or (_23152_, _23150_, _07229_);
  nor (_23153_, _11831_, _07120_);
  or (_23154_, _23153_, _23148_);
  or (_23155_, _23154_, _07142_);
  or (_23156_, _07897_, \oc8051_golden_model_1.TCON [1]);
  and (_23157_, _14503_, _07897_);
  not (_23158_, _23157_);
  and (_23159_, _23158_, _23156_);
  or (_23160_, _23159_, _06252_);
  and (_23161_, _07897_, \oc8051_golden_model_1.ACC [1]);
  or (_23163_, _23161_, _23148_);
  and (_23164_, _23163_, _07123_);
  nor (_23165_, _07123_, _23146_);
  or (_23166_, _23165_, _06251_);
  or (_23167_, _23166_, _23164_);
  and (_23168_, _23167_, _06476_);
  and (_23169_, _23168_, _23160_);
  nor (_23170_, _08528_, _23146_);
  and (_23171_, _14510_, _08528_);
  or (_23172_, _23171_, _23170_);
  and (_23174_, _23172_, _06475_);
  or (_23175_, _23174_, _06468_);
  or (_23176_, _23175_, _23169_);
  and (_23177_, _23176_, _23155_);
  or (_23178_, _23177_, _06466_);
  or (_23179_, _23163_, _06801_);
  and (_23180_, _23179_, _06484_);
  and (_23181_, _23180_, _23178_);
  and (_23182_, _14513_, _08528_);
  or (_23183_, _23182_, _23170_);
  and (_23185_, _23183_, _06483_);
  or (_23186_, _23185_, _06461_);
  or (_23187_, _23186_, _23181_);
  or (_23188_, _23170_, _14509_);
  and (_23189_, _23188_, _23172_);
  or (_23190_, _23189_, _07164_);
  and (_23191_, _23190_, _06242_);
  and (_23192_, _23191_, _23187_);
  or (_23193_, _23170_, _14553_);
  and (_23194_, _23193_, _06241_);
  and (_23196_, _23194_, _23172_);
  or (_23197_, _23196_, _07187_);
  or (_23198_, _23197_, _23192_);
  or (_23199_, _23154_, _07188_);
  and (_23200_, _23199_, _23198_);
  or (_23201_, _23200_, _07182_);
  and (_23202_, _09297_, _07897_);
  or (_23203_, _23148_, _07183_);
  or (_23204_, _23203_, _23202_);
  and (_23205_, _23204_, _06336_);
  and (_23207_, _23205_, _23201_);
  and (_23208_, _14609_, _07897_);
  or (_23209_, _23208_, _23148_);
  and (_23210_, _23209_, _05968_);
  or (_23211_, _23210_, _23207_);
  and (_23212_, _23211_, _07198_);
  nand (_23213_, _07897_, _07018_);
  and (_23214_, _23156_, _06371_);
  and (_23215_, _23214_, _23213_);
  or (_23216_, _23215_, _23212_);
  and (_23218_, _23216_, _07218_);
  or (_23219_, _14625_, _11831_);
  and (_23220_, _23156_, _06367_);
  and (_23221_, _23220_, _23219_);
  or (_23222_, _23221_, _06533_);
  or (_23223_, _23222_, _23218_);
  nand (_23224_, _11215_, _07897_);
  and (_23225_, _23224_, _23150_);
  or (_23226_, _23225_, _07216_);
  and (_23227_, _23226_, _07213_);
  and (_23229_, _23227_, _23223_);
  or (_23230_, _14623_, _11831_);
  and (_23231_, _23156_, _06366_);
  and (_23232_, _23231_, _23230_);
  or (_23233_, _23232_, _06541_);
  or (_23234_, _23233_, _23229_);
  nor (_23235_, _23148_, _07210_);
  nand (_23236_, _23235_, _23224_);
  and (_23237_, _23236_, _07231_);
  and (_23238_, _23237_, _23234_);
  or (_23240_, _23213_, _08302_);
  and (_23241_, _23156_, _06383_);
  and (_23242_, _23241_, _23240_);
  or (_23243_, _23242_, _06528_);
  or (_23244_, _23243_, _23238_);
  and (_23245_, _23244_, _23152_);
  or (_23246_, _23245_, _06563_);
  or (_23247_, _23159_, _07241_);
  and (_23248_, _23247_, _06571_);
  and (_23249_, _23248_, _23246_);
  and (_23251_, _23183_, _06199_);
  or (_23252_, _23251_, _06188_);
  or (_23253_, _23252_, _23249_);
  or (_23254_, _23148_, _06189_);
  or (_23255_, _23254_, _23157_);
  and (_23256_, _23255_, _01452_);
  and (_23257_, _23256_, _23253_);
  or (_23258_, _23257_, _23147_);
  and (_43829_, _23258_, _43223_);
  and (_23259_, _01456_, \oc8051_golden_model_1.TCON [2]);
  and (_23261_, _11831_, \oc8051_golden_model_1.TCON [2]);
  nor (_23262_, _11831_, _07578_);
  or (_23263_, _23262_, _23261_);
  or (_23264_, _23263_, _07188_);
  and (_23265_, _14712_, _07897_);
  or (_23266_, _23265_, _23261_);
  or (_23267_, _23266_, _06252_);
  and (_23268_, _07897_, \oc8051_golden_model_1.ACC [2]);
  or (_23269_, _23268_, _23261_);
  and (_23270_, _23269_, _07123_);
  and (_23272_, _07124_, \oc8051_golden_model_1.TCON [2]);
  or (_23273_, _23272_, _06251_);
  or (_23274_, _23273_, _23270_);
  and (_23275_, _23274_, _06476_);
  and (_23276_, _23275_, _23267_);
  and (_23277_, _11851_, \oc8051_golden_model_1.TCON [2]);
  and (_23278_, _14702_, _08528_);
  or (_23279_, _23278_, _23277_);
  and (_23280_, _23279_, _06475_);
  or (_23281_, _23280_, _06468_);
  or (_23283_, _23281_, _23276_);
  or (_23284_, _23263_, _07142_);
  and (_23285_, _23284_, _23283_);
  or (_23286_, _23285_, _06466_);
  or (_23287_, _23269_, _06801_);
  and (_23288_, _23287_, _06484_);
  and (_23289_, _23288_, _23286_);
  and (_23290_, _14706_, _08528_);
  or (_23291_, _23290_, _23277_);
  and (_23292_, _23291_, _06483_);
  or (_23294_, _23292_, _06461_);
  or (_23295_, _23294_, _23289_);
  or (_23296_, _23277_, _14739_);
  and (_23297_, _23296_, _23279_);
  or (_23298_, _23297_, _07164_);
  and (_23299_, _23298_, _06242_);
  and (_23300_, _23299_, _23295_);
  or (_23301_, _23277_, _14703_);
  and (_23302_, _23301_, _06241_);
  and (_23303_, _23302_, _23279_);
  or (_23305_, _23303_, _07187_);
  or (_23306_, _23305_, _23300_);
  and (_23307_, _23306_, _23264_);
  or (_23308_, _23307_, _07182_);
  and (_23309_, _09251_, _07897_);
  or (_23310_, _23261_, _07183_);
  or (_23311_, _23310_, _23309_);
  and (_23312_, _23311_, _06336_);
  and (_23313_, _23312_, _23308_);
  and (_23314_, _14808_, _07897_);
  or (_23316_, _23314_, _23261_);
  and (_23317_, _23316_, _05968_);
  or (_23318_, _23317_, _06371_);
  or (_23319_, _23318_, _23313_);
  and (_23320_, _07897_, _08945_);
  or (_23321_, _23320_, _23261_);
  or (_23322_, _23321_, _07198_);
  and (_23323_, _23322_, _23319_);
  or (_23324_, _23323_, _06367_);
  and (_23325_, _14824_, _07897_);
  or (_23327_, _23325_, _23261_);
  or (_23328_, _23327_, _07218_);
  and (_23329_, _23328_, _07216_);
  and (_23330_, _23329_, _23324_);
  and (_23331_, _11214_, _07897_);
  or (_23332_, _23331_, _23261_);
  and (_23333_, _23332_, _06533_);
  or (_23334_, _23333_, _23330_);
  and (_23335_, _23334_, _07213_);
  or (_23336_, _23261_, _08397_);
  and (_23338_, _23321_, _06366_);
  and (_23339_, _23338_, _23336_);
  or (_23340_, _23339_, _23335_);
  and (_23341_, _23340_, _07210_);
  and (_23342_, _23269_, _06541_);
  and (_23343_, _23342_, _23336_);
  or (_23344_, _23343_, _06383_);
  or (_23345_, _23344_, _23341_);
  and (_23346_, _14821_, _07897_);
  or (_23347_, _23261_, _07231_);
  or (_23349_, _23347_, _23346_);
  and (_23350_, _23349_, _07229_);
  and (_23351_, _23350_, _23345_);
  nor (_23352_, _11213_, _11831_);
  or (_23353_, _23352_, _23261_);
  and (_23354_, _23353_, _06528_);
  or (_23355_, _23354_, _06563_);
  or (_23356_, _23355_, _23351_);
  or (_23357_, _23266_, _07241_);
  and (_23358_, _23357_, _06571_);
  and (_23359_, _23358_, _23356_);
  and (_23360_, _23291_, _06199_);
  or (_23361_, _23360_, _06188_);
  or (_23362_, _23361_, _23359_);
  and (_23363_, _14884_, _07897_);
  or (_23364_, _23261_, _06189_);
  or (_23365_, _23364_, _23363_);
  and (_23366_, _23365_, _01452_);
  and (_23367_, _23366_, _23362_);
  or (_23368_, _23367_, _23259_);
  and (_43830_, _23368_, _43223_);
  and (_23371_, _01456_, \oc8051_golden_model_1.TCON [3]);
  and (_23372_, _11831_, \oc8051_golden_model_1.TCON [3]);
  nor (_23373_, _11831_, _07713_);
  or (_23374_, _23373_, _23372_);
  or (_23375_, _23374_, _07188_);
  or (_23376_, _23374_, _07142_);
  and (_23377_, _14898_, _07897_);
  or (_23378_, _23377_, _23372_);
  or (_23379_, _23378_, _06252_);
  and (_23381_, _07897_, \oc8051_golden_model_1.ACC [3]);
  or (_23382_, _23381_, _23372_);
  and (_23383_, _23382_, _07123_);
  and (_23384_, _07124_, \oc8051_golden_model_1.TCON [3]);
  or (_23385_, _23384_, _06251_);
  or (_23386_, _23385_, _23383_);
  and (_23387_, _23386_, _06476_);
  and (_23388_, _23387_, _23379_);
  and (_23389_, _11851_, \oc8051_golden_model_1.TCON [3]);
  and (_23390_, _14906_, _08528_);
  or (_23392_, _23390_, _23389_);
  and (_23393_, _23392_, _06475_);
  or (_23394_, _23393_, _06468_);
  or (_23395_, _23394_, _23388_);
  and (_23396_, _23395_, _23376_);
  or (_23397_, _23396_, _06466_);
  or (_23398_, _23382_, _06801_);
  and (_23399_, _23398_, _06484_);
  and (_23400_, _23399_, _23397_);
  and (_23401_, _14904_, _08528_);
  or (_23403_, _23401_, _23389_);
  and (_23404_, _23403_, _06483_);
  or (_23405_, _23404_, _06461_);
  or (_23406_, _23405_, _23400_);
  or (_23407_, _23389_, _14931_);
  and (_23408_, _23407_, _23392_);
  or (_23409_, _23408_, _07164_);
  and (_23410_, _23409_, _06242_);
  and (_23411_, _23410_, _23406_);
  or (_23412_, _23389_, _14947_);
  and (_23414_, _23412_, _06241_);
  and (_23415_, _23414_, _23392_);
  or (_23416_, _23415_, _07187_);
  or (_23417_, _23416_, _23411_);
  and (_23418_, _23417_, _23375_);
  or (_23419_, _23418_, _07182_);
  and (_23420_, _09205_, _07897_);
  or (_23421_, _23372_, _07183_);
  or (_23422_, _23421_, _23420_);
  and (_23423_, _23422_, _06336_);
  and (_23425_, _23423_, _23419_);
  and (_23426_, _15003_, _07897_);
  or (_23427_, _23426_, _23372_);
  and (_23428_, _23427_, _05968_);
  or (_23429_, _23428_, _06371_);
  or (_23430_, _23429_, _23425_);
  and (_23431_, _07897_, _08872_);
  or (_23432_, _23431_, _23372_);
  or (_23433_, _23432_, _07198_);
  and (_23434_, _23433_, _23430_);
  or (_23436_, _23434_, _06367_);
  and (_23437_, _15018_, _07897_);
  or (_23438_, _23437_, _23372_);
  or (_23439_, _23438_, _07218_);
  and (_23440_, _23439_, _07216_);
  and (_23441_, _23440_, _23436_);
  and (_23442_, _12523_, _07897_);
  or (_23443_, _23442_, _23372_);
  and (_23444_, _23443_, _06533_);
  or (_23445_, _23444_, _23441_);
  and (_23447_, _23445_, _07213_);
  or (_23448_, _23372_, _08257_);
  and (_23449_, _23432_, _06366_);
  and (_23450_, _23449_, _23448_);
  or (_23451_, _23450_, _23447_);
  and (_23452_, _23451_, _07210_);
  and (_23453_, _23382_, _06541_);
  and (_23454_, _23453_, _23448_);
  or (_23455_, _23454_, _06383_);
  or (_23456_, _23455_, _23452_);
  and (_23458_, _15015_, _07897_);
  or (_23459_, _23372_, _07231_);
  or (_23460_, _23459_, _23458_);
  and (_23461_, _23460_, _07229_);
  and (_23462_, _23461_, _23456_);
  nor (_23463_, _11211_, _11831_);
  or (_23464_, _23463_, _23372_);
  and (_23465_, _23464_, _06528_);
  or (_23466_, _23465_, _06563_);
  or (_23467_, _23466_, _23462_);
  or (_23469_, _23378_, _07241_);
  and (_23470_, _23469_, _06571_);
  and (_23471_, _23470_, _23467_);
  and (_23472_, _23403_, _06199_);
  or (_23473_, _23472_, _06188_);
  or (_23474_, _23473_, _23471_);
  and (_23475_, _15075_, _07897_);
  or (_23476_, _23372_, _06189_);
  or (_23477_, _23476_, _23475_);
  and (_23478_, _23477_, _01452_);
  and (_23480_, _23478_, _23474_);
  or (_23481_, _23480_, _23371_);
  and (_43832_, _23481_, _43223_);
  and (_23482_, _01456_, \oc8051_golden_model_1.TCON [4]);
  and (_23483_, _11831_, \oc8051_golden_model_1.TCON [4]);
  nor (_23484_, _08494_, _11831_);
  or (_23485_, _23484_, _23483_);
  or (_23486_, _23485_, _07188_);
  and (_23487_, _11851_, \oc8051_golden_model_1.TCON [4]);
  and (_23488_, _15089_, _08528_);
  or (_23490_, _23488_, _23487_);
  and (_23491_, _23490_, _06483_);
  or (_23492_, _23485_, _07142_);
  and (_23493_, _15108_, _07897_);
  or (_23494_, _23493_, _23483_);
  or (_23495_, _23494_, _06252_);
  and (_23496_, _07897_, \oc8051_golden_model_1.ACC [4]);
  or (_23497_, _23496_, _23483_);
  and (_23498_, _23497_, _07123_);
  and (_23499_, _07124_, \oc8051_golden_model_1.TCON [4]);
  or (_23501_, _23499_, _06251_);
  or (_23502_, _23501_, _23498_);
  and (_23503_, _23502_, _06476_);
  and (_23504_, _23503_, _23495_);
  and (_23505_, _15091_, _08528_);
  or (_23506_, _23505_, _23487_);
  and (_23507_, _23506_, _06475_);
  or (_23508_, _23507_, _06468_);
  or (_23509_, _23508_, _23504_);
  and (_23510_, _23509_, _23492_);
  or (_23512_, _23510_, _06466_);
  or (_23513_, _23497_, _06801_);
  and (_23514_, _23513_, _06484_);
  and (_23515_, _23514_, _23512_);
  or (_23516_, _23515_, _23491_);
  and (_23517_, _23516_, _07164_);
  or (_23518_, _23487_, _15125_);
  and (_23519_, _23518_, _06461_);
  and (_23520_, _23519_, _23506_);
  or (_23521_, _23520_, _23517_);
  and (_23523_, _23521_, _06242_);
  or (_23524_, _23487_, _15141_);
  and (_23525_, _23524_, _06241_);
  and (_23526_, _23525_, _23506_);
  or (_23527_, _23526_, _07187_);
  or (_23528_, _23527_, _23523_);
  and (_23529_, _23528_, _23486_);
  or (_23530_, _23529_, _07182_);
  and (_23531_, _09159_, _07897_);
  or (_23532_, _23483_, _07183_);
  or (_23534_, _23532_, _23531_);
  and (_23535_, _23534_, _06336_);
  and (_23536_, _23535_, _23530_);
  and (_23537_, _15198_, _07897_);
  or (_23538_, _23537_, _23483_);
  and (_23539_, _23538_, _05968_);
  or (_23540_, _23539_, _06371_);
  or (_23541_, _23540_, _23536_);
  and (_23542_, _08892_, _07897_);
  or (_23543_, _23542_, _23483_);
  or (_23545_, _23543_, _07198_);
  and (_23546_, _23545_, _23541_);
  or (_23547_, _23546_, _06367_);
  and (_23548_, _15214_, _07897_);
  or (_23549_, _23548_, _23483_);
  or (_23550_, _23549_, _07218_);
  and (_23551_, _23550_, _07216_);
  and (_23552_, _23551_, _23547_);
  and (_23553_, _11209_, _07897_);
  or (_23554_, _23553_, _23483_);
  and (_23556_, _23554_, _06533_);
  or (_23557_, _23556_, _23552_);
  and (_23558_, _23557_, _07213_);
  or (_23559_, _23483_, _08497_);
  and (_23560_, _23543_, _06366_);
  and (_23561_, _23560_, _23559_);
  or (_23562_, _23561_, _23558_);
  and (_23563_, _23562_, _07210_);
  and (_23564_, _23497_, _06541_);
  and (_23565_, _23564_, _23559_);
  or (_23567_, _23565_, _06383_);
  or (_23568_, _23567_, _23563_);
  and (_23569_, _15211_, _07897_);
  or (_23570_, _23483_, _07231_);
  or (_23571_, _23570_, _23569_);
  and (_23572_, _23571_, _07229_);
  and (_23573_, _23572_, _23568_);
  nor (_23574_, _11208_, _11831_);
  or (_23575_, _23574_, _23483_);
  and (_23576_, _23575_, _06528_);
  or (_23578_, _23576_, _06563_);
  or (_23579_, _23578_, _23573_);
  or (_23580_, _23494_, _07241_);
  and (_23581_, _23580_, _06571_);
  and (_23582_, _23581_, _23579_);
  and (_23583_, _23490_, _06199_);
  or (_23584_, _23583_, _06188_);
  or (_23585_, _23584_, _23582_);
  and (_23586_, _15280_, _07897_);
  or (_23587_, _23483_, _06189_);
  or (_23589_, _23587_, _23586_);
  and (_23590_, _23589_, _01452_);
  and (_23591_, _23590_, _23585_);
  or (_23592_, _23591_, _23482_);
  and (_43833_, _23592_, _43223_);
  and (_23593_, _01456_, \oc8051_golden_model_1.TCON [5]);
  and (_23594_, _11831_, \oc8051_golden_model_1.TCON [5]);
  nor (_23595_, _08209_, _11831_);
  or (_23596_, _23595_, _23594_);
  or (_23597_, _23596_, _07142_);
  and (_23599_, _15311_, _07897_);
  or (_23600_, _23599_, _23594_);
  or (_23601_, _23600_, _06252_);
  and (_23602_, _07897_, \oc8051_golden_model_1.ACC [5]);
  or (_23603_, _23602_, _23594_);
  and (_23604_, _23603_, _07123_);
  and (_23605_, _07124_, \oc8051_golden_model_1.TCON [5]);
  or (_23606_, _23605_, _06251_);
  or (_23607_, _23606_, _23604_);
  and (_23608_, _23607_, _06476_);
  and (_23610_, _23608_, _23601_);
  and (_23611_, _11851_, \oc8051_golden_model_1.TCON [5]);
  and (_23612_, _15296_, _08528_);
  or (_23613_, _23612_, _23611_);
  and (_23614_, _23613_, _06475_);
  or (_23615_, _23614_, _06468_);
  or (_23616_, _23615_, _23610_);
  and (_23617_, _23616_, _23597_);
  or (_23618_, _23617_, _06466_);
  or (_23619_, _23603_, _06801_);
  and (_23621_, _23619_, _06484_);
  and (_23622_, _23621_, _23618_);
  and (_23623_, _15294_, _08528_);
  or (_23624_, _23623_, _23611_);
  and (_23625_, _23624_, _06483_);
  or (_23626_, _23625_, _06461_);
  or (_23627_, _23626_, _23622_);
  or (_23628_, _23611_, _15328_);
  and (_23629_, _23628_, _23613_);
  or (_23630_, _23629_, _07164_);
  and (_23631_, _23630_, _06242_);
  and (_23632_, _23631_, _23627_);
  or (_23633_, _23611_, _15344_);
  and (_23634_, _23633_, _06241_);
  and (_23635_, _23634_, _23613_);
  or (_23636_, _23635_, _07187_);
  or (_23637_, _23636_, _23632_);
  or (_23638_, _23596_, _07188_);
  and (_23639_, _23638_, _23637_);
  or (_23640_, _23639_, _07182_);
  and (_23642_, _09113_, _07897_);
  or (_23643_, _23594_, _07183_);
  or (_23644_, _23643_, _23642_);
  and (_23645_, _23644_, _06336_);
  and (_23646_, _23645_, _23640_);
  and (_23647_, _15400_, _07897_);
  or (_23648_, _23647_, _23594_);
  and (_23649_, _23648_, _05968_);
  or (_23650_, _23649_, _06371_);
  or (_23651_, _23650_, _23646_);
  and (_23653_, _08888_, _07897_);
  or (_23654_, _23653_, _23594_);
  or (_23655_, _23654_, _07198_);
  and (_23656_, _23655_, _23651_);
  or (_23657_, _23656_, _06367_);
  and (_23658_, _15416_, _07897_);
  or (_23659_, _23658_, _23594_);
  or (_23660_, _23659_, _07218_);
  and (_23661_, _23660_, _07216_);
  and (_23662_, _23661_, _23657_);
  and (_23664_, _11205_, _07897_);
  or (_23665_, _23664_, _23594_);
  and (_23666_, _23665_, _06533_);
  or (_23667_, _23666_, _23662_);
  and (_23668_, _23667_, _07213_);
  or (_23669_, _23594_, _08212_);
  and (_23670_, _23654_, _06366_);
  and (_23671_, _23670_, _23669_);
  or (_23672_, _23671_, _23668_);
  and (_23673_, _23672_, _07210_);
  and (_23674_, _23603_, _06541_);
  and (_23675_, _23674_, _23669_);
  or (_23676_, _23675_, _06383_);
  or (_23677_, _23676_, _23673_);
  and (_23678_, _15413_, _07897_);
  or (_23679_, _23594_, _07231_);
  or (_23680_, _23679_, _23678_);
  and (_23681_, _23680_, _07229_);
  and (_23682_, _23681_, _23677_);
  nor (_23683_, _11204_, _11831_);
  or (_23685_, _23683_, _23594_);
  and (_23686_, _23685_, _06528_);
  or (_23687_, _23686_, _06563_);
  or (_23688_, _23687_, _23682_);
  or (_23689_, _23600_, _07241_);
  and (_23690_, _23689_, _06571_);
  and (_23691_, _23690_, _23688_);
  and (_23692_, _23624_, _06199_);
  or (_23693_, _23692_, _06188_);
  or (_23694_, _23693_, _23691_);
  and (_23695_, _15477_, _07897_);
  or (_23696_, _23594_, _06189_);
  or (_23697_, _23696_, _23695_);
  and (_23698_, _23697_, _01452_);
  and (_23699_, _23698_, _23694_);
  or (_23700_, _23699_, _23593_);
  and (_43834_, _23700_, _43223_);
  and (_23701_, _01456_, \oc8051_golden_model_1.TCON [6]);
  and (_23702_, _11831_, \oc8051_golden_model_1.TCON [6]);
  nor (_23703_, _08106_, _11831_);
  or (_23705_, _23703_, _23702_);
  or (_23706_, _23705_, _07142_);
  and (_23707_, _15512_, _07897_);
  or (_23708_, _23707_, _23702_);
  or (_23709_, _23708_, _06252_);
  and (_23710_, _07897_, \oc8051_golden_model_1.ACC [6]);
  or (_23711_, _23710_, _23702_);
  and (_23712_, _23711_, _07123_);
  and (_23713_, _07124_, \oc8051_golden_model_1.TCON [6]);
  or (_23714_, _23713_, _06251_);
  or (_23716_, _23714_, _23712_);
  and (_23717_, _23716_, _06476_);
  and (_23718_, _23717_, _23709_);
  and (_23719_, _11851_, \oc8051_golden_model_1.TCON [6]);
  and (_23720_, _15499_, _08528_);
  or (_23721_, _23720_, _23719_);
  and (_23722_, _23721_, _06475_);
  or (_23723_, _23722_, _06468_);
  or (_23724_, _23723_, _23718_);
  and (_23725_, _23724_, _23706_);
  or (_23726_, _23725_, _06466_);
  or (_23727_, _23711_, _06801_);
  and (_23728_, _23727_, _06484_);
  and (_23729_, _23728_, _23726_);
  and (_23730_, _15497_, _08528_);
  or (_23731_, _23730_, _23719_);
  and (_23732_, _23731_, _06483_);
  or (_23733_, _23732_, _06461_);
  or (_23734_, _23733_, _23729_);
  or (_23735_, _23719_, _15529_);
  and (_23737_, _23735_, _23721_);
  or (_23738_, _23737_, _07164_);
  and (_23739_, _23738_, _06242_);
  and (_23740_, _23739_, _23734_);
  or (_23741_, _23719_, _15545_);
  and (_23742_, _23741_, _06241_);
  and (_23743_, _23742_, _23721_);
  or (_23744_, _23743_, _07187_);
  or (_23745_, _23744_, _23740_);
  or (_23746_, _23705_, _07188_);
  and (_23748_, _23746_, _23745_);
  or (_23749_, _23748_, _07182_);
  and (_23750_, _09067_, _07897_);
  or (_23751_, _23702_, _07183_);
  or (_23752_, _23751_, _23750_);
  and (_23753_, _23752_, _06336_);
  and (_23754_, _23753_, _23749_);
  and (_23755_, _15601_, _07897_);
  or (_23756_, _23755_, _23702_);
  and (_23757_, _23756_, _05968_);
  or (_23758_, _23757_, _06371_);
  or (_23759_, _23758_, _23754_);
  and (_23760_, _15608_, _07897_);
  or (_23761_, _23760_, _23702_);
  or (_23762_, _23761_, _07198_);
  and (_23763_, _23762_, _23759_);
  or (_23764_, _23763_, _06367_);
  and (_23765_, _15618_, _07897_);
  or (_23766_, _23765_, _23702_);
  or (_23767_, _23766_, _07218_);
  and (_23769_, _23767_, _07216_);
  and (_23770_, _23769_, _23764_);
  and (_23771_, _11202_, _07897_);
  or (_23772_, _23771_, _23702_);
  and (_23773_, _23772_, _06533_);
  or (_23774_, _23773_, _23770_);
  and (_23775_, _23774_, _07213_);
  or (_23776_, _23702_, _08109_);
  and (_23777_, _23761_, _06366_);
  and (_23778_, _23777_, _23776_);
  or (_23780_, _23778_, _23775_);
  and (_23781_, _23780_, _07210_);
  and (_23782_, _23711_, _06541_);
  and (_23783_, _23782_, _23776_);
  or (_23784_, _23783_, _06383_);
  or (_23785_, _23784_, _23781_);
  and (_23786_, _15615_, _07897_);
  or (_23787_, _23702_, _07231_);
  or (_23788_, _23787_, _23786_);
  and (_23789_, _23788_, _07229_);
  and (_23790_, _23789_, _23785_);
  nor (_23791_, _11201_, _11831_);
  or (_23792_, _23791_, _23702_);
  and (_23793_, _23792_, _06528_);
  or (_23794_, _23793_, _06563_);
  or (_23795_, _23794_, _23790_);
  or (_23796_, _23708_, _07241_);
  and (_23797_, _23796_, _06571_);
  and (_23798_, _23797_, _23795_);
  and (_23799_, _23731_, _06199_);
  or (_23801_, _23799_, _06188_);
  or (_23802_, _23801_, _23798_);
  and (_23803_, _15676_, _07897_);
  or (_23804_, _23702_, _06189_);
  or (_23805_, _23804_, _23803_);
  and (_23806_, _23805_, _01452_);
  and (_23807_, _23806_, _23802_);
  or (_23808_, _23807_, _23701_);
  and (_43835_, _23808_, _43223_);
  and (_23809_, _01456_, \oc8051_golden_model_1.TH1 [0]);
  and (_23811_, _07879_, \oc8051_golden_model_1.ACC [0]);
  and (_23812_, _23811_, _08351_);
  and (_23813_, _11933_, \oc8051_golden_model_1.TH1 [0]);
  or (_23814_, _23813_, _07210_);
  or (_23815_, _23814_, _23812_);
  and (_23816_, _07879_, _07325_);
  or (_23817_, _23816_, _23813_);
  or (_23818_, _23817_, _07188_);
  nor (_23819_, _08351_, _11933_);
  or (_23820_, _23819_, _23813_);
  or (_23821_, _23820_, _06252_);
  or (_23822_, _23813_, _23811_);
  and (_23823_, _23822_, _07123_);
  and (_23824_, _07124_, \oc8051_golden_model_1.TH1 [0]);
  or (_23825_, _23824_, _06251_);
  or (_23826_, _23825_, _23823_);
  and (_23827_, _23826_, _07142_);
  and (_23828_, _23827_, _23821_);
  and (_23829_, _23817_, _06468_);
  or (_23830_, _23829_, _23828_);
  and (_23832_, _23830_, _06801_);
  and (_23833_, _23822_, _06466_);
  or (_23834_, _23833_, _07187_);
  or (_23835_, _23834_, _23832_);
  and (_23836_, _23835_, _23818_);
  or (_23837_, _23836_, _07182_);
  and (_23838_, _09342_, _07879_);
  or (_23839_, _23813_, _07183_);
  or (_23840_, _23839_, _23838_);
  and (_23841_, _23840_, _23837_);
  or (_23843_, _23841_, _05968_);
  and (_23844_, _14427_, _07879_);
  or (_23845_, _23813_, _06336_);
  or (_23846_, _23845_, _23844_);
  and (_23847_, _23846_, _07198_);
  and (_23848_, _23847_, _23843_);
  and (_23849_, _07879_, _08908_);
  or (_23850_, _23849_, _23813_);
  and (_23851_, _23850_, _06371_);
  or (_23852_, _23851_, _06367_);
  or (_23853_, _23852_, _23848_);
  and (_23854_, _14442_, _07879_);
  or (_23855_, _23854_, _23813_);
  or (_23856_, _23855_, _07218_);
  and (_23857_, _23856_, _07216_);
  and (_23858_, _23857_, _23853_);
  nor (_23859_, _12526_, _11933_);
  or (_23860_, _23859_, _23813_);
  nor (_23861_, _23812_, _07216_);
  and (_23862_, _23861_, _23860_);
  or (_23864_, _23862_, _23858_);
  and (_23865_, _23864_, _07213_);
  nand (_23866_, _23850_, _06366_);
  nor (_23867_, _23866_, _23819_);
  or (_23868_, _23867_, _06541_);
  or (_23869_, _23868_, _23865_);
  and (_23870_, _23869_, _23815_);
  or (_23871_, _23870_, _06383_);
  and (_23872_, _14325_, _07879_);
  or (_23873_, _23813_, _07231_);
  or (_23875_, _23873_, _23872_);
  and (_23876_, _23875_, _07229_);
  and (_23877_, _23876_, _23871_);
  and (_23878_, _23860_, _06528_);
  or (_23879_, _23878_, _19442_);
  or (_23880_, _23879_, _23877_);
  or (_23881_, _23820_, _06756_);
  and (_23882_, _23881_, _01452_);
  and (_23883_, _23882_, _23880_);
  or (_23884_, _23883_, _23809_);
  and (_43837_, _23884_, _43223_);
  and (_23885_, _01456_, \oc8051_golden_model_1.TH1 [1]);
  nand (_23886_, _07879_, _07018_);
  or (_23887_, _07879_, \oc8051_golden_model_1.TH1 [1]);
  and (_23888_, _23887_, _06371_);
  and (_23889_, _23888_, _23886_);
  and (_23890_, _09297_, _07879_);
  and (_23891_, _11933_, \oc8051_golden_model_1.TH1 [1]);
  or (_23892_, _23891_, _07183_);
  or (_23893_, _23892_, _23890_);
  nor (_23895_, _11933_, _07120_);
  or (_23896_, _23891_, _19463_);
  or (_23897_, _23896_, _23895_);
  and (_23898_, _07879_, \oc8051_golden_model_1.ACC [1]);
  or (_23899_, _23898_, _23891_);
  and (_23900_, _23899_, _06466_);
  or (_23901_, _23900_, _07187_);
  and (_23902_, _14503_, _07879_);
  not (_23903_, _23902_);
  and (_23904_, _23903_, _23887_);
  and (_23906_, _23904_, _06251_);
  and (_23907_, _07124_, \oc8051_golden_model_1.TH1 [1]);
  and (_23908_, _23899_, _07123_);
  or (_23909_, _23908_, _23907_);
  and (_23910_, _23909_, _06252_);
  or (_23911_, _23910_, _06468_);
  or (_23912_, _23911_, _23906_);
  and (_23913_, _23912_, _06801_);
  or (_23914_, _23913_, _23901_);
  and (_23915_, _23914_, _23897_);
  or (_23916_, _23915_, _07182_);
  and (_23917_, _23916_, _06336_);
  and (_23918_, _23917_, _23893_);
  or (_23919_, _14609_, _11933_);
  and (_23920_, _23887_, _05968_);
  and (_23921_, _23920_, _23919_);
  or (_23922_, _23921_, _23918_);
  and (_23923_, _23922_, _07198_);
  or (_23924_, _23923_, _23889_);
  and (_23925_, _23924_, _07218_);
  or (_23927_, _14625_, _11933_);
  and (_23928_, _23887_, _06367_);
  and (_23929_, _23928_, _23927_);
  or (_23930_, _23929_, _06533_);
  or (_23931_, _23930_, _23925_);
  and (_23932_, _11217_, _07879_);
  or (_23933_, _23932_, _23891_);
  or (_23934_, _23933_, _07216_);
  and (_23935_, _23934_, _07213_);
  and (_23936_, _23935_, _23931_);
  or (_23938_, _14623_, _11933_);
  and (_23939_, _23887_, _06366_);
  and (_23940_, _23939_, _23938_);
  or (_23941_, _23940_, _06541_);
  or (_23942_, _23941_, _23936_);
  and (_23943_, _23898_, _08302_);
  or (_23944_, _23891_, _07210_);
  or (_23945_, _23944_, _23943_);
  and (_23946_, _23945_, _07231_);
  and (_23947_, _23946_, _23942_);
  or (_23948_, _23886_, _08302_);
  and (_23949_, _23887_, _06383_);
  and (_23950_, _23949_, _23948_);
  or (_23951_, _23950_, _06528_);
  or (_23952_, _23951_, _23947_);
  nor (_23953_, _11216_, _11933_);
  or (_23954_, _23953_, _23891_);
  or (_23955_, _23954_, _07229_);
  and (_23956_, _23955_, _07241_);
  and (_23957_, _23956_, _23952_);
  and (_23959_, _23904_, _06563_);
  or (_23960_, _23959_, _06188_);
  or (_23961_, _23960_, _23957_);
  or (_23962_, _23891_, _06189_);
  or (_23963_, _23962_, _23902_);
  and (_23964_, _23963_, _01452_);
  and (_23965_, _23964_, _23961_);
  or (_23966_, _23965_, _23885_);
  and (_43838_, _23966_, _43223_);
  and (_23967_, _01456_, \oc8051_golden_model_1.TH1 [2]);
  and (_23968_, _11933_, \oc8051_golden_model_1.TH1 [2]);
  and (_23969_, _09251_, _07879_);
  or (_23970_, _23969_, _23968_);
  and (_23971_, _23970_, _07182_);
  and (_23972_, _14712_, _07879_);
  or (_23973_, _23972_, _23968_);
  or (_23974_, _23973_, _06252_);
  and (_23975_, _07879_, \oc8051_golden_model_1.ACC [2]);
  or (_23976_, _23975_, _23968_);
  and (_23977_, _23976_, _07123_);
  and (_23979_, _07124_, \oc8051_golden_model_1.TH1 [2]);
  or (_23980_, _23979_, _06251_);
  or (_23981_, _23980_, _23977_);
  and (_23982_, _23981_, _07142_);
  and (_23983_, _23982_, _23974_);
  nor (_23984_, _11933_, _07578_);
  or (_23985_, _23984_, _23968_);
  and (_23986_, _23985_, _06468_);
  or (_23987_, _23986_, _23983_);
  and (_23988_, _23987_, _06801_);
  and (_23990_, _23976_, _06466_);
  or (_23991_, _23990_, _07187_);
  or (_23992_, _23991_, _23988_);
  or (_23993_, _23985_, _07188_);
  and (_23994_, _23993_, _07183_);
  and (_23995_, _23994_, _23992_);
  or (_23996_, _23995_, _05968_);
  or (_23997_, _23996_, _23971_);
  and (_23998_, _14808_, _07879_);
  or (_23999_, _23968_, _06336_);
  or (_24001_, _23999_, _23998_);
  and (_24002_, _24001_, _07198_);
  and (_24003_, _24002_, _23997_);
  and (_24004_, _07879_, _08945_);
  or (_24005_, _24004_, _23968_);
  and (_24006_, _24005_, _06371_);
  or (_24007_, _24006_, _06367_);
  or (_24008_, _24007_, _24003_);
  and (_24009_, _14824_, _07879_);
  or (_24010_, _24009_, _23968_);
  or (_24011_, _24010_, _07218_);
  and (_24012_, _24011_, _07216_);
  and (_24013_, _24012_, _24008_);
  and (_24014_, _11214_, _07879_);
  or (_24015_, _24014_, _23968_);
  and (_24016_, _24015_, _06533_);
  or (_24017_, _24016_, _24013_);
  and (_24018_, _24017_, _07213_);
  or (_24019_, _23968_, _08397_);
  and (_24020_, _24005_, _06366_);
  and (_24022_, _24020_, _24019_);
  or (_24023_, _24022_, _24018_);
  and (_24024_, _24023_, _07210_);
  and (_24025_, _23976_, _06541_);
  and (_24026_, _24025_, _24019_);
  or (_24027_, _24026_, _06383_);
  or (_24028_, _24027_, _24024_);
  and (_24029_, _14821_, _07879_);
  or (_24030_, _23968_, _07231_);
  or (_24031_, _24030_, _24029_);
  and (_24033_, _24031_, _07229_);
  and (_24034_, _24033_, _24028_);
  nor (_24035_, _11213_, _11933_);
  or (_24036_, _24035_, _23968_);
  and (_24037_, _24036_, _06528_);
  or (_24038_, _24037_, _24034_);
  and (_24039_, _24038_, _07241_);
  and (_24040_, _23973_, _06563_);
  or (_24041_, _24040_, _06188_);
  or (_24042_, _24041_, _24039_);
  and (_24044_, _14884_, _07879_);
  or (_24045_, _23968_, _06189_);
  or (_24046_, _24045_, _24044_);
  and (_24047_, _24046_, _01452_);
  and (_24048_, _24047_, _24042_);
  or (_24049_, _24048_, _23967_);
  and (_43839_, _24049_, _43223_);
  and (_24050_, _11933_, \oc8051_golden_model_1.TH1 [3]);
  and (_24051_, _14898_, _07879_);
  or (_24052_, _24051_, _24050_);
  or (_24053_, _24052_, _06252_);
  and (_24054_, _07879_, \oc8051_golden_model_1.ACC [3]);
  or (_24055_, _24054_, _24050_);
  and (_24056_, _24055_, _07123_);
  and (_24057_, _07124_, \oc8051_golden_model_1.TH1 [3]);
  or (_24058_, _24057_, _06251_);
  or (_24059_, _24058_, _24056_);
  and (_24060_, _24059_, _07142_);
  and (_24061_, _24060_, _24053_);
  nor (_24062_, _11933_, _07713_);
  or (_24064_, _24062_, _24050_);
  and (_24065_, _24064_, _06468_);
  or (_24066_, _24065_, _24061_);
  and (_24067_, _24066_, _06801_);
  and (_24068_, _24055_, _06466_);
  or (_24069_, _24068_, _07187_);
  or (_24070_, _24069_, _24067_);
  or (_24071_, _24064_, _07188_);
  and (_24072_, _24071_, _07183_);
  and (_24073_, _24072_, _24070_);
  and (_24075_, _09205_, _07879_);
  or (_24076_, _24075_, _24050_);
  and (_24077_, _24076_, _07182_);
  or (_24078_, _24077_, _05968_);
  or (_24079_, _24078_, _24073_);
  and (_24080_, _15003_, _07879_);
  or (_24081_, _24050_, _06336_);
  or (_24082_, _24081_, _24080_);
  and (_24083_, _24082_, _07198_);
  and (_24084_, _24083_, _24079_);
  and (_24085_, _07879_, _08872_);
  or (_24086_, _24085_, _24050_);
  and (_24087_, _24086_, _06371_);
  or (_24088_, _24087_, _06367_);
  or (_24089_, _24088_, _24084_);
  and (_24090_, _15018_, _07879_);
  or (_24091_, _24090_, _24050_);
  or (_24092_, _24091_, _07218_);
  and (_24093_, _24092_, _07216_);
  and (_24094_, _24093_, _24089_);
  and (_24096_, _12523_, _07879_);
  or (_24097_, _24096_, _24050_);
  and (_24098_, _24097_, _06533_);
  or (_24099_, _24098_, _24094_);
  and (_24100_, _24099_, _07213_);
  or (_24101_, _24050_, _08257_);
  and (_24102_, _24086_, _06366_);
  and (_24103_, _24102_, _24101_);
  or (_24104_, _24103_, _24100_);
  and (_24105_, _24104_, _07210_);
  and (_24107_, _24055_, _06541_);
  and (_24108_, _24107_, _24101_);
  or (_24109_, _24108_, _06383_);
  or (_24110_, _24109_, _24105_);
  and (_24111_, _15015_, _07879_);
  or (_24112_, _24050_, _07231_);
  or (_24113_, _24112_, _24111_);
  and (_24114_, _24113_, _07229_);
  and (_24115_, _24114_, _24110_);
  nor (_24116_, _11211_, _11933_);
  or (_24118_, _24116_, _24050_);
  and (_24119_, _24118_, _06528_);
  or (_24120_, _24119_, _06563_);
  or (_24121_, _24120_, _24115_);
  or (_24122_, _24052_, _07241_);
  and (_24123_, _24122_, _06189_);
  and (_24124_, _24123_, _24121_);
  and (_24125_, _15075_, _07879_);
  or (_24126_, _24125_, _24050_);
  and (_24127_, _24126_, _06188_);
  or (_24128_, _24127_, _01456_);
  or (_24129_, _24128_, _24124_);
  or (_24130_, _01452_, \oc8051_golden_model_1.TH1 [3]);
  and (_24131_, _24130_, _43223_);
  and (_43840_, _24131_, _24129_);
  and (_24132_, _11933_, \oc8051_golden_model_1.TH1 [4]);
  nor (_24133_, _08494_, _11933_);
  or (_24134_, _24133_, _24132_);
  or (_24135_, _24134_, _07188_);
  and (_24136_, _15108_, _07879_);
  or (_24138_, _24136_, _24132_);
  or (_24139_, _24138_, _06252_);
  and (_24140_, _07879_, \oc8051_golden_model_1.ACC [4]);
  or (_24141_, _24140_, _24132_);
  and (_24142_, _24141_, _07123_);
  and (_24143_, _07124_, \oc8051_golden_model_1.TH1 [4]);
  or (_24144_, _24143_, _06251_);
  or (_24145_, _24144_, _24142_);
  and (_24146_, _24145_, _07142_);
  and (_24147_, _24146_, _24139_);
  and (_24149_, _24134_, _06468_);
  or (_24150_, _24149_, _24147_);
  and (_24151_, _24150_, _06801_);
  and (_24152_, _24141_, _06466_);
  or (_24153_, _24152_, _07187_);
  or (_24154_, _24153_, _24151_);
  and (_24155_, _24154_, _24135_);
  or (_24156_, _24155_, _07182_);
  and (_24157_, _09159_, _07879_);
  or (_24158_, _24132_, _07183_);
  or (_24159_, _24158_, _24157_);
  and (_24160_, _24159_, _24156_);
  or (_24161_, _24160_, _05968_);
  and (_24162_, _15198_, _07879_);
  or (_24163_, _24132_, _06336_);
  or (_24164_, _24163_, _24162_);
  and (_24165_, _24164_, _07198_);
  and (_24166_, _24165_, _24161_);
  and (_24167_, _08892_, _07879_);
  or (_24168_, _24167_, _24132_);
  and (_24170_, _24168_, _06371_);
  or (_24171_, _24170_, _06367_);
  or (_24172_, _24171_, _24166_);
  and (_24173_, _15214_, _07879_);
  or (_24174_, _24173_, _24132_);
  or (_24175_, _24174_, _07218_);
  and (_24176_, _24175_, _07216_);
  and (_24177_, _24176_, _24172_);
  and (_24178_, _11209_, _07879_);
  or (_24179_, _24178_, _24132_);
  and (_24181_, _24179_, _06533_);
  or (_24182_, _24181_, _24177_);
  and (_24183_, _24182_, _07213_);
  or (_24184_, _24132_, _08497_);
  and (_24185_, _24168_, _06366_);
  and (_24186_, _24185_, _24184_);
  or (_24187_, _24186_, _24183_);
  and (_24188_, _24187_, _07210_);
  and (_24189_, _24141_, _06541_);
  and (_24190_, _24189_, _24184_);
  or (_24192_, _24190_, _06383_);
  or (_24193_, _24192_, _24188_);
  and (_24194_, _15211_, _07879_);
  or (_24195_, _24132_, _07231_);
  or (_24196_, _24195_, _24194_);
  and (_24197_, _24196_, _07229_);
  and (_24198_, _24197_, _24193_);
  nor (_24199_, _11208_, _11933_);
  or (_24200_, _24199_, _24132_);
  and (_24201_, _24200_, _06528_);
  or (_24203_, _24201_, _06563_);
  or (_24204_, _24203_, _24198_);
  or (_24205_, _24138_, _07241_);
  and (_24206_, _24205_, _06189_);
  and (_24207_, _24206_, _24204_);
  and (_24208_, _15280_, _07879_);
  or (_24209_, _24208_, _24132_);
  and (_24210_, _24209_, _06188_);
  or (_24211_, _24210_, _01456_);
  or (_24212_, _24211_, _24207_);
  or (_24214_, _01452_, \oc8051_golden_model_1.TH1 [4]);
  and (_24215_, _24214_, _43223_);
  and (_43841_, _24215_, _24212_);
  and (_24216_, _11933_, \oc8051_golden_model_1.TH1 [5]);
  and (_24217_, _15311_, _07879_);
  or (_24218_, _24217_, _24216_);
  or (_24219_, _24218_, _06252_);
  and (_24220_, _07879_, \oc8051_golden_model_1.ACC [5]);
  or (_24221_, _24220_, _24216_);
  and (_24222_, _24221_, _07123_);
  and (_24224_, _07124_, \oc8051_golden_model_1.TH1 [5]);
  or (_24225_, _24224_, _06251_);
  or (_24226_, _24225_, _24222_);
  and (_24227_, _24226_, _07142_);
  and (_24228_, _24227_, _24219_);
  nor (_24229_, _08209_, _11933_);
  or (_24230_, _24229_, _24216_);
  and (_24231_, _24230_, _06468_);
  or (_24232_, _24231_, _24228_);
  and (_24233_, _24232_, _06801_);
  and (_24235_, _24221_, _06466_);
  or (_24236_, _24235_, _07187_);
  or (_24237_, _24236_, _24233_);
  or (_24238_, _24230_, _07188_);
  and (_24239_, _24238_, _24237_);
  or (_24240_, _24239_, _07182_);
  and (_24241_, _09113_, _07879_);
  or (_24242_, _24216_, _07183_);
  or (_24243_, _24242_, _24241_);
  and (_24244_, _24243_, _06336_);
  and (_24246_, _24244_, _24240_);
  and (_24247_, _15400_, _07879_);
  or (_24248_, _24247_, _24216_);
  and (_24249_, _24248_, _05968_);
  or (_24250_, _24249_, _06371_);
  or (_24251_, _24250_, _24246_);
  and (_24252_, _08888_, _07879_);
  or (_24253_, _24252_, _24216_);
  or (_24254_, _24253_, _07198_);
  and (_24255_, _24254_, _24251_);
  or (_24257_, _24255_, _06367_);
  and (_24258_, _15416_, _07879_);
  or (_24259_, _24258_, _24216_);
  or (_24260_, _24259_, _07218_);
  and (_24261_, _24260_, _07216_);
  and (_24262_, _24261_, _24257_);
  and (_24263_, _11205_, _07879_);
  or (_24264_, _24263_, _24216_);
  and (_24265_, _24264_, _06533_);
  or (_24266_, _24265_, _24262_);
  and (_24268_, _24266_, _07213_);
  or (_24269_, _24216_, _08212_);
  and (_24270_, _24253_, _06366_);
  and (_24271_, _24270_, _24269_);
  or (_24272_, _24271_, _24268_);
  and (_24273_, _24272_, _07210_);
  and (_24274_, _24221_, _06541_);
  and (_24275_, _24274_, _24269_);
  or (_24276_, _24275_, _06383_);
  or (_24277_, _24276_, _24273_);
  and (_24278_, _15413_, _07879_);
  or (_24279_, _24216_, _07231_);
  or (_24280_, _24279_, _24278_);
  and (_24281_, _24280_, _07229_);
  and (_24282_, _24281_, _24277_);
  nor (_24283_, _11204_, _11933_);
  or (_24284_, _24283_, _24216_);
  and (_24285_, _24284_, _06528_);
  or (_24286_, _24285_, _06563_);
  or (_24287_, _24286_, _24282_);
  or (_24289_, _24218_, _07241_);
  and (_24290_, _24289_, _06189_);
  and (_24291_, _24290_, _24287_);
  and (_24292_, _15477_, _07879_);
  or (_24293_, _24292_, _24216_);
  and (_24294_, _24293_, _06188_);
  or (_24295_, _24294_, _01456_);
  or (_24296_, _24295_, _24291_);
  or (_24297_, _01452_, \oc8051_golden_model_1.TH1 [5]);
  and (_24298_, _24297_, _43223_);
  and (_43842_, _24298_, _24296_);
  and (_24300_, _11933_, \oc8051_golden_model_1.TH1 [6]);
  nor (_24301_, _08106_, _11933_);
  or (_24302_, _24301_, _24300_);
  or (_24303_, _24302_, _07188_);
  and (_24304_, _15512_, _07879_);
  or (_24305_, _24304_, _24300_);
  or (_24306_, _24305_, _06252_);
  and (_24307_, _07879_, \oc8051_golden_model_1.ACC [6]);
  or (_24308_, _24307_, _24300_);
  and (_24310_, _24308_, _07123_);
  and (_24311_, _07124_, \oc8051_golden_model_1.TH1 [6]);
  or (_24312_, _24311_, _06251_);
  or (_24313_, _24312_, _24310_);
  and (_24314_, _24313_, _07142_);
  and (_24315_, _24314_, _24306_);
  and (_24316_, _24302_, _06468_);
  or (_24317_, _24316_, _24315_);
  and (_24318_, _24317_, _06801_);
  and (_24319_, _24308_, _06466_);
  or (_24321_, _24319_, _07187_);
  or (_24322_, _24321_, _24318_);
  and (_24323_, _24322_, _24303_);
  or (_24324_, _24323_, _07182_);
  and (_24325_, _09067_, _07879_);
  or (_24326_, _24300_, _07183_);
  or (_24327_, _24326_, _24325_);
  and (_24328_, _24327_, _06336_);
  and (_24329_, _24328_, _24324_);
  and (_24330_, _15601_, _07879_);
  or (_24332_, _24330_, _24300_);
  and (_24333_, _24332_, _05968_);
  or (_24334_, _24333_, _06371_);
  or (_24335_, _24334_, _24329_);
  and (_24336_, _15608_, _07879_);
  or (_24337_, _24336_, _24300_);
  or (_24338_, _24337_, _07198_);
  and (_24339_, _24338_, _24335_);
  or (_24340_, _24339_, _06367_);
  and (_24341_, _15618_, _07879_);
  or (_24343_, _24341_, _24300_);
  or (_24344_, _24343_, _07218_);
  and (_24345_, _24344_, _07216_);
  and (_24346_, _24345_, _24340_);
  and (_24347_, _11202_, _07879_);
  or (_24348_, _24347_, _24300_);
  and (_24349_, _24348_, _06533_);
  or (_24350_, _24349_, _24346_);
  and (_24351_, _24350_, _07213_);
  or (_24352_, _24300_, _08109_);
  and (_24354_, _24337_, _06366_);
  and (_24355_, _24354_, _24352_);
  or (_24356_, _24355_, _24351_);
  and (_24357_, _24356_, _07210_);
  and (_24358_, _24308_, _06541_);
  and (_24359_, _24358_, _24352_);
  or (_24360_, _24359_, _06383_);
  or (_24361_, _24360_, _24357_);
  and (_24362_, _15615_, _07879_);
  or (_24363_, _24300_, _07231_);
  or (_24365_, _24363_, _24362_);
  and (_24366_, _24365_, _07229_);
  and (_24367_, _24366_, _24361_);
  nor (_24368_, _11201_, _11933_);
  or (_24369_, _24368_, _24300_);
  and (_24370_, _24369_, _06528_);
  or (_24371_, _24370_, _06563_);
  or (_24372_, _24371_, _24367_);
  or (_24373_, _24305_, _07241_);
  and (_24374_, _24373_, _06189_);
  and (_24376_, _24374_, _24372_);
  and (_24377_, _15676_, _07879_);
  or (_24378_, _24377_, _24300_);
  and (_24379_, _24378_, _06188_);
  or (_24380_, _24379_, _01456_);
  or (_24381_, _24380_, _24376_);
  or (_24382_, _01452_, \oc8051_golden_model_1.TH1 [6]);
  and (_24383_, _24382_, _43223_);
  and (_43843_, _24383_, _24381_);
  and (_24384_, _01456_, \oc8051_golden_model_1.TH0 [0]);
  and (_24386_, _07889_, \oc8051_golden_model_1.ACC [0]);
  and (_24387_, _24386_, _08351_);
  and (_24388_, _12011_, \oc8051_golden_model_1.TH0 [0]);
  or (_24389_, _24388_, _07210_);
  or (_24390_, _24389_, _24387_);
  or (_24391_, _24388_, _24386_);
  and (_24392_, _24391_, _06466_);
  or (_24393_, _24392_, _07187_);
  nor (_24394_, _08351_, _12011_);
  or (_24395_, _24394_, _24388_);
  and (_24397_, _24395_, _06251_);
  and (_24398_, _07124_, \oc8051_golden_model_1.TH0 [0]);
  and (_24399_, _24391_, _07123_);
  or (_24400_, _24399_, _24398_);
  and (_24401_, _24400_, _06252_);
  or (_24402_, _24401_, _06468_);
  or (_24403_, _24402_, _24397_);
  and (_24404_, _24403_, _06801_);
  or (_24405_, _24404_, _24393_);
  and (_24406_, _07889_, _07325_);
  or (_24408_, _24388_, _19463_);
  or (_24409_, _24408_, _24406_);
  and (_24410_, _24409_, _24405_);
  or (_24411_, _24410_, _07182_);
  and (_24412_, _09342_, _07889_);
  or (_24413_, _24388_, _07183_);
  or (_24414_, _24413_, _24412_);
  and (_24415_, _24414_, _24411_);
  or (_24416_, _24415_, _05968_);
  and (_24417_, _14427_, _07889_);
  or (_24419_, _24388_, _06336_);
  or (_24420_, _24419_, _24417_);
  and (_24421_, _24420_, _07198_);
  and (_24422_, _24421_, _24416_);
  and (_24423_, _07889_, _08908_);
  or (_24424_, _24423_, _24388_);
  and (_24425_, _24424_, _06371_);
  or (_24426_, _24425_, _06367_);
  or (_24427_, _24426_, _24422_);
  and (_24428_, _14442_, _07889_);
  or (_24430_, _24428_, _24388_);
  or (_24431_, _24430_, _07218_);
  and (_24432_, _24431_, _07216_);
  and (_24433_, _24432_, _24427_);
  nor (_24434_, _12526_, _12011_);
  or (_24435_, _24434_, _24388_);
  nor (_24436_, _24387_, _07216_);
  and (_24437_, _24436_, _24435_);
  or (_24438_, _24437_, _24433_);
  and (_24439_, _24438_, _07213_);
  nand (_24441_, _24424_, _06366_);
  nor (_24442_, _24441_, _24394_);
  or (_24443_, _24442_, _06541_);
  or (_24444_, _24443_, _24439_);
  and (_24445_, _24444_, _24390_);
  or (_24446_, _24445_, _06383_);
  and (_24447_, _14325_, _07889_);
  or (_24448_, _24388_, _07231_);
  or (_24449_, _24448_, _24447_);
  and (_24450_, _24449_, _07229_);
  and (_24452_, _24450_, _24446_);
  and (_24453_, _24435_, _06528_);
  or (_24454_, _24453_, _19442_);
  or (_24455_, _24454_, _24452_);
  or (_24456_, _24395_, _06756_);
  and (_24457_, _24456_, _01452_);
  and (_24458_, _24457_, _24455_);
  or (_24459_, _24458_, _24384_);
  and (_43845_, _24459_, _43223_);
  not (_24460_, \oc8051_golden_model_1.TH0 [1]);
  nor (_24462_, _01452_, _24460_);
  or (_24463_, _07889_, \oc8051_golden_model_1.TH0 [1]);
  and (_24464_, _14503_, _07889_);
  not (_24465_, _24464_);
  and (_24466_, _24465_, _24463_);
  or (_24467_, _24466_, _06252_);
  nor (_24468_, _07889_, _24460_);
  and (_24469_, _07889_, \oc8051_golden_model_1.ACC [1]);
  or (_24470_, _24469_, _24468_);
  and (_24471_, _24470_, _07123_);
  nor (_24473_, _07123_, _24460_);
  or (_24474_, _24473_, _06251_);
  or (_24475_, _24474_, _24471_);
  and (_24476_, _24475_, _07142_);
  and (_24477_, _24476_, _24467_);
  nor (_24478_, _12011_, _07120_);
  or (_24479_, _24478_, _24468_);
  and (_24480_, _24479_, _06468_);
  or (_24481_, _24480_, _24477_);
  and (_24482_, _24481_, _06801_);
  and (_24484_, _24470_, _06466_);
  or (_24485_, _24484_, _07187_);
  or (_24486_, _24485_, _24482_);
  or (_24487_, _24479_, _07188_);
  and (_24488_, _24487_, _07183_);
  and (_24489_, _24488_, _24486_);
  or (_24490_, _09297_, _12011_);
  and (_24491_, _24463_, _07182_);
  and (_24492_, _24491_, _24490_);
  or (_24493_, _24492_, _24489_);
  and (_24494_, _24493_, _06336_);
  or (_24495_, _14609_, _12011_);
  and (_24496_, _24463_, _05968_);
  and (_24497_, _24496_, _24495_);
  or (_24498_, _24497_, _24494_);
  and (_24499_, _24498_, _07198_);
  nand (_24500_, _07889_, _07018_);
  and (_24501_, _24463_, _06371_);
  and (_24502_, _24501_, _24500_);
  or (_24503_, _24502_, _24499_);
  and (_24506_, _24503_, _07218_);
  or (_24507_, _14625_, _12011_);
  and (_24508_, _24463_, _06367_);
  and (_24509_, _24508_, _24507_);
  or (_24510_, _24509_, _06533_);
  or (_24511_, _24510_, _24506_);
  nor (_24512_, _11216_, _12011_);
  or (_24513_, _24512_, _24468_);
  nand (_24514_, _11215_, _07889_);
  and (_24515_, _24514_, _24513_);
  or (_24517_, _24515_, _07216_);
  and (_24518_, _24517_, _07213_);
  and (_24519_, _24518_, _24511_);
  or (_24520_, _14623_, _12011_);
  and (_24521_, _24463_, _06366_);
  and (_24522_, _24521_, _24520_);
  or (_24523_, _24522_, _06541_);
  or (_24524_, _24523_, _24519_);
  nor (_24525_, _24468_, _07210_);
  nand (_24526_, _24525_, _24514_);
  and (_24528_, _24526_, _07231_);
  and (_24529_, _24528_, _24524_);
  or (_24530_, _24500_, _08302_);
  and (_24531_, _24463_, _06383_);
  and (_24532_, _24531_, _24530_);
  or (_24533_, _24532_, _06528_);
  or (_24534_, _24533_, _24529_);
  or (_24535_, _24513_, _07229_);
  and (_24536_, _24535_, _07241_);
  and (_24537_, _24536_, _24534_);
  and (_24539_, _24466_, _06563_);
  or (_24540_, _24539_, _06188_);
  or (_24541_, _24540_, _24537_);
  or (_24542_, _24468_, _06189_);
  or (_24543_, _24542_, _24464_);
  and (_24544_, _24543_, _01452_);
  and (_24545_, _24544_, _24541_);
  or (_24546_, _24545_, _24462_);
  and (_43846_, _24546_, _43223_);
  and (_24547_, _01456_, \oc8051_golden_model_1.TH0 [2]);
  and (_24549_, _12011_, \oc8051_golden_model_1.TH0 [2]);
  and (_24550_, _09251_, _07889_);
  or (_24551_, _24550_, _24549_);
  and (_24552_, _24551_, _07182_);
  and (_24553_, _14712_, _07889_);
  or (_24554_, _24553_, _24549_);
  or (_24555_, _24554_, _06252_);
  and (_24556_, _07889_, \oc8051_golden_model_1.ACC [2]);
  or (_24557_, _24556_, _24549_);
  and (_24558_, _24557_, _07123_);
  and (_24560_, _07124_, \oc8051_golden_model_1.TH0 [2]);
  or (_24561_, _24560_, _06251_);
  or (_24562_, _24561_, _24558_);
  and (_24563_, _24562_, _07142_);
  and (_24564_, _24563_, _24555_);
  nor (_24565_, _12011_, _07578_);
  or (_24566_, _24565_, _24549_);
  and (_24567_, _24566_, _06468_);
  or (_24568_, _24567_, _24564_);
  and (_24569_, _24568_, _06801_);
  and (_24571_, _24557_, _06466_);
  or (_24572_, _24571_, _07187_);
  or (_24573_, _24572_, _24569_);
  or (_24574_, _24566_, _07188_);
  and (_24575_, _24574_, _07183_);
  and (_24576_, _24575_, _24573_);
  or (_24577_, _24576_, _05968_);
  or (_24578_, _24577_, _24552_);
  and (_24579_, _14808_, _07889_);
  or (_24580_, _24549_, _06336_);
  or (_24582_, _24580_, _24579_);
  and (_24583_, _24582_, _07198_);
  and (_24584_, _24583_, _24578_);
  and (_24585_, _07889_, _08945_);
  or (_24586_, _24585_, _24549_);
  and (_24587_, _24586_, _06371_);
  or (_24588_, _24587_, _06367_);
  or (_24589_, _24588_, _24584_);
  and (_24590_, _14824_, _07889_);
  or (_24591_, _24590_, _24549_);
  or (_24593_, _24591_, _07218_);
  and (_24594_, _24593_, _07216_);
  and (_24595_, _24594_, _24589_);
  and (_24596_, _11214_, _07889_);
  or (_24597_, _24596_, _24549_);
  and (_24598_, _24597_, _06533_);
  or (_24599_, _24598_, _24595_);
  and (_24600_, _24599_, _07213_);
  or (_24601_, _24549_, _08397_);
  and (_24602_, _24586_, _06366_);
  and (_24604_, _24602_, _24601_);
  or (_24605_, _24604_, _24600_);
  and (_24606_, _24605_, _07210_);
  and (_24607_, _24557_, _06541_);
  and (_24608_, _24607_, _24601_);
  or (_24609_, _24608_, _06383_);
  or (_24610_, _24609_, _24606_);
  and (_24611_, _14821_, _07889_);
  or (_24612_, _24549_, _07231_);
  or (_24613_, _24612_, _24611_);
  and (_24615_, _24613_, _07229_);
  and (_24616_, _24615_, _24610_);
  nor (_24617_, _11213_, _12011_);
  or (_24618_, _24617_, _24549_);
  and (_24619_, _24618_, _06528_);
  or (_24620_, _24619_, _24616_);
  and (_24621_, _24620_, _07241_);
  and (_24622_, _24554_, _06563_);
  or (_24623_, _24622_, _06188_);
  or (_24624_, _24623_, _24621_);
  and (_24626_, _14884_, _07889_);
  or (_24627_, _24549_, _06189_);
  or (_24628_, _24627_, _24626_);
  and (_24629_, _24628_, _01452_);
  and (_24630_, _24629_, _24624_);
  or (_24631_, _24630_, _24547_);
  and (_43847_, _24631_, _43223_);
  and (_24632_, _12011_, \oc8051_golden_model_1.TH0 [3]);
  and (_24633_, _14898_, _07889_);
  or (_24634_, _24633_, _24632_);
  or (_24636_, _24634_, _06252_);
  and (_24637_, _07889_, \oc8051_golden_model_1.ACC [3]);
  or (_24638_, _24637_, _24632_);
  and (_24639_, _24638_, _07123_);
  and (_24640_, _07124_, \oc8051_golden_model_1.TH0 [3]);
  or (_24641_, _24640_, _06251_);
  or (_24642_, _24641_, _24639_);
  and (_24643_, _24642_, _07142_);
  and (_24644_, _24643_, _24636_);
  nor (_24645_, _12011_, _07713_);
  or (_24647_, _24645_, _24632_);
  and (_24648_, _24647_, _06468_);
  or (_24649_, _24648_, _24644_);
  and (_24650_, _24649_, _06801_);
  and (_24651_, _24638_, _06466_);
  or (_24652_, _24651_, _07187_);
  or (_24653_, _24652_, _24650_);
  or (_24654_, _24647_, _07188_);
  and (_24655_, _24654_, _24653_);
  or (_24656_, _24655_, _07182_);
  and (_24658_, _09205_, _07889_);
  or (_24659_, _24632_, _07183_);
  or (_24660_, _24659_, _24658_);
  and (_24661_, _24660_, _06336_);
  and (_24662_, _24661_, _24656_);
  and (_24663_, _15003_, _07889_);
  or (_24664_, _24663_, _24632_);
  and (_24665_, _24664_, _05968_);
  or (_24666_, _24665_, _06371_);
  or (_24667_, _24666_, _24662_);
  and (_24669_, _07889_, _08872_);
  or (_24670_, _24669_, _24632_);
  or (_24671_, _24670_, _07198_);
  and (_24672_, _24671_, _24667_);
  or (_24673_, _24672_, _06367_);
  and (_24674_, _15018_, _07889_);
  or (_24675_, _24674_, _24632_);
  or (_24676_, _24675_, _07218_);
  and (_24677_, _24676_, _07216_);
  and (_24678_, _24677_, _24673_);
  and (_24680_, _12523_, _07889_);
  or (_24681_, _24680_, _24632_);
  and (_24682_, _24681_, _06533_);
  or (_24683_, _24682_, _24678_);
  and (_24684_, _24683_, _07213_);
  or (_24685_, _24632_, _08257_);
  and (_24686_, _24670_, _06366_);
  and (_24687_, _24686_, _24685_);
  or (_24688_, _24687_, _24684_);
  and (_24689_, _24688_, _07210_);
  and (_24691_, _24638_, _06541_);
  and (_24692_, _24691_, _24685_);
  or (_24693_, _24692_, _06383_);
  or (_24694_, _24693_, _24689_);
  and (_24695_, _15015_, _07889_);
  or (_24696_, _24632_, _07231_);
  or (_24697_, _24696_, _24695_);
  and (_24698_, _24697_, _07229_);
  and (_24699_, _24698_, _24694_);
  nor (_24700_, _11211_, _12011_);
  or (_24702_, _24700_, _24632_);
  and (_24703_, _24702_, _06528_);
  or (_24704_, _24703_, _06563_);
  or (_24705_, _24704_, _24699_);
  or (_24706_, _24634_, _07241_);
  and (_24707_, _24706_, _06189_);
  and (_24708_, _24707_, _24705_);
  and (_24709_, _15075_, _07889_);
  or (_24710_, _24709_, _24632_);
  and (_24711_, _24710_, _06188_);
  or (_24713_, _24711_, _01456_);
  or (_24714_, _24713_, _24708_);
  or (_24715_, _01452_, \oc8051_golden_model_1.TH0 [3]);
  and (_24716_, _24715_, _43223_);
  and (_43848_, _24716_, _24714_);
  and (_24717_, _12011_, \oc8051_golden_model_1.TH0 [4]);
  and (_24718_, _15108_, _07889_);
  or (_24719_, _24718_, _24717_);
  or (_24720_, _24719_, _06252_);
  and (_24721_, _07889_, \oc8051_golden_model_1.ACC [4]);
  or (_24723_, _24721_, _24717_);
  and (_24724_, _24723_, _07123_);
  and (_24725_, _07124_, \oc8051_golden_model_1.TH0 [4]);
  or (_24726_, _24725_, _06251_);
  or (_24727_, _24726_, _24724_);
  and (_24728_, _24727_, _07142_);
  and (_24729_, _24728_, _24720_);
  nor (_24730_, _08494_, _12011_);
  or (_24731_, _24730_, _24717_);
  and (_24732_, _24731_, _06468_);
  or (_24734_, _24732_, _24729_);
  and (_24735_, _24734_, _06801_);
  and (_24736_, _24723_, _06466_);
  or (_24737_, _24736_, _07187_);
  or (_24738_, _24737_, _24735_);
  or (_24739_, _24731_, _07188_);
  and (_24740_, _24739_, _24738_);
  or (_24741_, _24740_, _07182_);
  and (_24742_, _09159_, _07889_);
  or (_24743_, _24717_, _07183_);
  or (_24745_, _24743_, _24742_);
  and (_24746_, _24745_, _24741_);
  or (_24747_, _24746_, _05968_);
  and (_24748_, _15198_, _07889_);
  or (_24749_, _24717_, _06336_);
  or (_24750_, _24749_, _24748_);
  and (_24751_, _24750_, _07198_);
  and (_24752_, _24751_, _24747_);
  and (_24753_, _08892_, _07889_);
  or (_24754_, _24753_, _24717_);
  and (_24756_, _24754_, _06371_);
  or (_24757_, _24756_, _06367_);
  or (_24758_, _24757_, _24752_);
  and (_24759_, _15214_, _07889_);
  or (_24760_, _24759_, _24717_);
  or (_24761_, _24760_, _07218_);
  and (_24762_, _24761_, _07216_);
  and (_24763_, _24762_, _24758_);
  and (_24764_, _11209_, _07889_);
  or (_24765_, _24764_, _24717_);
  and (_24767_, _24765_, _06533_);
  or (_24768_, _24767_, _24763_);
  and (_24769_, _24768_, _07213_);
  or (_24770_, _24717_, _08497_);
  and (_24771_, _24754_, _06366_);
  and (_24772_, _24771_, _24770_);
  or (_24773_, _24772_, _24769_);
  and (_24774_, _24773_, _07210_);
  and (_24775_, _24723_, _06541_);
  and (_24776_, _24775_, _24770_);
  or (_24778_, _24776_, _06383_);
  or (_24779_, _24778_, _24774_);
  and (_24780_, _15211_, _07889_);
  or (_24781_, _24717_, _07231_);
  or (_24782_, _24781_, _24780_);
  and (_24783_, _24782_, _07229_);
  and (_24784_, _24783_, _24779_);
  nor (_24785_, _11208_, _12011_);
  or (_24786_, _24785_, _24717_);
  and (_24787_, _24786_, _06528_);
  or (_24789_, _24787_, _06563_);
  or (_24790_, _24789_, _24784_);
  or (_24791_, _24719_, _07241_);
  and (_24792_, _24791_, _06189_);
  and (_24793_, _24792_, _24790_);
  and (_24794_, _15280_, _07889_);
  or (_24795_, _24794_, _24717_);
  and (_24796_, _24795_, _06188_);
  or (_24797_, _24796_, _01456_);
  or (_24798_, _24797_, _24793_);
  or (_24800_, _01452_, \oc8051_golden_model_1.TH0 [4]);
  and (_24801_, _24800_, _43223_);
  and (_43849_, _24801_, _24798_);
  and (_24802_, _12011_, \oc8051_golden_model_1.TH0 [5]);
  nor (_24803_, _08209_, _12011_);
  or (_24804_, _24803_, _24802_);
  or (_24805_, _24804_, _07188_);
  and (_24806_, _15311_, _07889_);
  or (_24807_, _24806_, _24802_);
  or (_24808_, _24807_, _06252_);
  and (_24810_, _07889_, \oc8051_golden_model_1.ACC [5]);
  or (_24811_, _24810_, _24802_);
  and (_24812_, _24811_, _07123_);
  and (_24813_, _07124_, \oc8051_golden_model_1.TH0 [5]);
  or (_24814_, _24813_, _06251_);
  or (_24815_, _24814_, _24812_);
  and (_24816_, _24815_, _07142_);
  and (_24817_, _24816_, _24808_);
  and (_24818_, _24804_, _06468_);
  or (_24819_, _24818_, _24817_);
  and (_24821_, _24819_, _06801_);
  and (_24822_, _24811_, _06466_);
  or (_24823_, _24822_, _07187_);
  or (_24824_, _24823_, _24821_);
  and (_24825_, _24824_, _24805_);
  or (_24826_, _24825_, _07182_);
  and (_24827_, _09113_, _07889_);
  or (_24828_, _24802_, _07183_);
  or (_24829_, _24828_, _24827_);
  and (_24830_, _24829_, _06336_);
  and (_24832_, _24830_, _24826_);
  and (_24833_, _15400_, _07889_);
  or (_24834_, _24833_, _24802_);
  and (_24835_, _24834_, _05968_);
  or (_24836_, _24835_, _06371_);
  or (_24837_, _24836_, _24832_);
  and (_24838_, _08888_, _07889_);
  or (_24839_, _24838_, _24802_);
  or (_24840_, _24839_, _07198_);
  and (_24841_, _24840_, _24837_);
  or (_24843_, _24841_, _06367_);
  and (_24844_, _15416_, _07889_);
  or (_24845_, _24844_, _24802_);
  or (_24846_, _24845_, _07218_);
  and (_24847_, _24846_, _07216_);
  and (_24848_, _24847_, _24843_);
  and (_24849_, _11205_, _07889_);
  or (_24850_, _24849_, _24802_);
  and (_24851_, _24850_, _06533_);
  or (_24852_, _24851_, _24848_);
  and (_24854_, _24852_, _07213_);
  or (_24855_, _24802_, _08212_);
  and (_24856_, _24839_, _06366_);
  and (_24857_, _24856_, _24855_);
  or (_24858_, _24857_, _24854_);
  and (_24859_, _24858_, _07210_);
  and (_24860_, _24811_, _06541_);
  and (_24861_, _24860_, _24855_);
  or (_24862_, _24861_, _06383_);
  or (_24863_, _24862_, _24859_);
  and (_24865_, _15413_, _07889_);
  or (_24866_, _24802_, _07231_);
  or (_24867_, _24866_, _24865_);
  and (_24868_, _24867_, _07229_);
  and (_24869_, _24868_, _24863_);
  nor (_24870_, _11204_, _12011_);
  or (_24871_, _24870_, _24802_);
  and (_24872_, _24871_, _06528_);
  or (_24873_, _24872_, _06563_);
  or (_24874_, _24873_, _24869_);
  or (_24876_, _24807_, _07241_);
  and (_24877_, _24876_, _06189_);
  and (_24878_, _24877_, _24874_);
  and (_24879_, _15477_, _07889_);
  or (_24880_, _24879_, _24802_);
  and (_24881_, _24880_, _06188_);
  or (_24882_, _24881_, _01456_);
  or (_24883_, _24882_, _24878_);
  or (_24884_, _01452_, \oc8051_golden_model_1.TH0 [5]);
  and (_24885_, _24884_, _43223_);
  and (_43851_, _24885_, _24883_);
  and (_24887_, _12011_, \oc8051_golden_model_1.TH0 [6]);
  nor (_24888_, _08106_, _12011_);
  or (_24889_, _24888_, _24887_);
  or (_24890_, _24889_, _07188_);
  and (_24891_, _15512_, _07889_);
  or (_24892_, _24891_, _24887_);
  or (_24893_, _24892_, _06252_);
  and (_24894_, _07889_, \oc8051_golden_model_1.ACC [6]);
  or (_24895_, _24894_, _24887_);
  and (_24897_, _24895_, _07123_);
  and (_24898_, _07124_, \oc8051_golden_model_1.TH0 [6]);
  or (_24899_, _24898_, _06251_);
  or (_24900_, _24899_, _24897_);
  and (_24901_, _24900_, _07142_);
  and (_24902_, _24901_, _24893_);
  and (_24903_, _24889_, _06468_);
  or (_24904_, _24903_, _24902_);
  and (_24905_, _24904_, _06801_);
  and (_24906_, _24895_, _06466_);
  or (_24908_, _24906_, _07187_);
  or (_24909_, _24908_, _24905_);
  and (_24910_, _24909_, _24890_);
  or (_24911_, _24910_, _07182_);
  and (_24912_, _09067_, _07889_);
  or (_24913_, _24887_, _07183_);
  or (_24914_, _24913_, _24912_);
  and (_24915_, _24914_, _06336_);
  and (_24916_, _24915_, _24911_);
  and (_24917_, _15601_, _07889_);
  or (_24919_, _24917_, _24887_);
  and (_24920_, _24919_, _05968_);
  or (_24921_, _24920_, _06371_);
  or (_24922_, _24921_, _24916_);
  and (_24923_, _15608_, _07889_);
  or (_24924_, _24923_, _24887_);
  or (_24925_, _24924_, _07198_);
  and (_24926_, _24925_, _24922_);
  or (_24927_, _24926_, _06367_);
  and (_24928_, _15618_, _07889_);
  or (_24930_, _24928_, _24887_);
  or (_24931_, _24930_, _07218_);
  and (_24932_, _24931_, _07216_);
  and (_24933_, _24932_, _24927_);
  and (_24934_, _11202_, _07889_);
  or (_24935_, _24934_, _24887_);
  and (_24936_, _24935_, _06533_);
  or (_24937_, _24936_, _24933_);
  and (_24938_, _24937_, _07213_);
  or (_24939_, _24887_, _08109_);
  and (_24941_, _24924_, _06366_);
  and (_24942_, _24941_, _24939_);
  or (_24943_, _24942_, _24938_);
  and (_24944_, _24943_, _07210_);
  and (_24945_, _24895_, _06541_);
  and (_24946_, _24945_, _24939_);
  or (_24947_, _24946_, _06383_);
  or (_24948_, _24947_, _24944_);
  and (_24949_, _15615_, _07889_);
  or (_24950_, _24887_, _07231_);
  or (_24952_, _24950_, _24949_);
  and (_24953_, _24952_, _07229_);
  and (_24954_, _24953_, _24948_);
  nor (_24955_, _11201_, _12011_);
  or (_24956_, _24955_, _24887_);
  and (_24957_, _24956_, _06528_);
  or (_24958_, _24957_, _06563_);
  or (_24959_, _24958_, _24954_);
  or (_24960_, _24892_, _07241_);
  and (_24961_, _24960_, _06189_);
  and (_24963_, _24961_, _24959_);
  and (_24964_, _15676_, _07889_);
  or (_24965_, _24964_, _24887_);
  and (_24966_, _24965_, _06188_);
  or (_24967_, _24966_, _01456_);
  or (_24968_, _24967_, _24963_);
  or (_24969_, _01452_, \oc8051_golden_model_1.TH0 [6]);
  and (_24970_, _24969_, _43223_);
  and (_43852_, _24970_, _24968_);
  and (_24971_, _13025_, _05557_);
  and (_24973_, _12954_, \oc8051_golden_model_1.PC [0]);
  and (_24974_, _06912_, \oc8051_golden_model_1.PC [0]);
  nor (_24975_, _24974_, _12312_);
  nor (_24976_, _24975_, _12954_);
  nor (_24977_, _24976_, _24973_);
  and (_24978_, _24977_, _06199_);
  and (_24979_, _12984_, _12991_);
  nor (_24980_, _24979_, _05557_);
  and (_24981_, _12105_, _12966_);
  nor (_24982_, _24981_, _05557_);
  and (_24984_, _12756_, _11081_);
  nor (_24985_, _24984_, _05557_);
  nor (_24986_, _06912_, _05922_);
  and (_24987_, _12736_, _07231_);
  nor (_24988_, _24987_, _05557_);
  nor (_24989_, _10855_, _05557_);
  and (_24990_, _10855_, _05557_);
  nor (_24991_, _24990_, _24989_);
  nor (_24992_, _24991_, _12724_);
  and (_24993_, _12226_, _07213_);
  nor (_24995_, _24993_, _05557_);
  and (_24996_, _12232_, _07218_);
  nor (_24997_, _24996_, _05557_);
  and (_24998_, _06371_, _05557_);
  nor (_24999_, _06912_, _08723_);
  and (_25000_, _12533_, _05557_);
  not (_25001_, _24975_);
  nor (_25002_, _25001_, _12533_);
  nor (_25003_, _25002_, _25000_);
  nor (_25004_, _25003_, _12536_);
  and (_25006_, _12392_, _05557_);
  not (_25007_, _25006_);
  nor (_25008_, _25001_, _12392_);
  nor (_25009_, _25008_, _06345_);
  and (_25010_, _25009_, _25007_);
  nor (_25011_, _06912_, _05953_);
  and (_25012_, _06912_, _06705_);
  nor (_25013_, _12427_, _05557_);
  nor (_25014_, _12420_, _05557_);
  and (_25015_, _12420_, _05557_);
  nor (_25017_, _25015_, _25014_);
  and (_25018_, _12427_, _07272_);
  not (_25019_, _25018_);
  nor (_25020_, _25019_, _25017_);
  nor (_25021_, _25020_, _25013_);
  not (_25022_, _25021_);
  nor (_25023_, _25022_, _25012_);
  nor (_25024_, _25023_, _08572_);
  and (_25025_, _12412_, \oc8051_golden_model_1.PC [0]);
  and (_25026_, _06802_, _05557_);
  nor (_25028_, _25026_, _12160_);
  and (_25029_, _25028_, _12414_);
  or (_25030_, _25029_, _25025_);
  nor (_25031_, _25030_, _08573_);
  nor (_25032_, _25031_, _25024_);
  nor (_25033_, _25032_, _07134_);
  and (_25034_, _07134_, \oc8051_golden_model_1.PC [0]);
  nor (_25035_, _25034_, _25033_);
  and (_25036_, _25035_, _06252_);
  and (_25037_, _12402_, _05557_);
  and (_25038_, _24975_, _12404_);
  or (_25039_, _25038_, _25037_);
  and (_25040_, _25039_, _06251_);
  nor (_25041_, _25040_, _12444_);
  not (_25042_, _25041_);
  nor (_25043_, _25042_, _25036_);
  nor (_25044_, _12443_, _05557_);
  nor (_25045_, _25044_, _07474_);
  not (_25046_, _25045_);
  nor (_25047_, _25046_, _25043_);
  nor (_25050_, _06912_, _05950_);
  and (_25051_, _12462_, _12451_);
  not (_25052_, _25051_);
  nor (_25053_, _25052_, _25050_);
  not (_25054_, _25053_);
  nor (_25055_, _25054_, _25047_);
  nor (_25056_, _25051_, _05557_);
  nor (_25057_, _25056_, _12466_);
  not (_25058_, _25057_);
  nor (_25059_, _25058_, _25055_);
  or (_25061_, _25059_, _12479_);
  nor (_25062_, _25061_, _25011_);
  and (_25063_, _12513_, _05557_);
  not (_25064_, _25063_);
  nor (_25065_, _25001_, _12513_);
  nor (_25066_, _25065_, _12478_);
  and (_25067_, _25066_, _25064_);
  nor (_25068_, _25067_, _25062_);
  nor (_25069_, _25068_, _06344_);
  nor (_25070_, _25069_, _06338_);
  not (_25072_, _25070_);
  nor (_25073_, _25072_, _25010_);
  nor (_25074_, _25073_, _25004_);
  nor (_25075_, _25074_, _06373_);
  and (_25076_, _12555_, _05557_);
  nor (_25077_, _25001_, _12555_);
  or (_25078_, _25077_, _25076_);
  and (_25079_, _25078_, _06373_);
  or (_25080_, _25079_, _25075_);
  and (_25081_, _25080_, _12246_);
  and (_25083_, _12245_, _05557_);
  or (_25084_, _25083_, _25081_);
  and (_25085_, _25084_, _05947_);
  nor (_25086_, _06912_, _05947_);
  nor (_25087_, _25086_, _12243_);
  not (_25088_, _25087_);
  nor (_25089_, _25088_, _25085_);
  not (_25090_, _05958_);
  nor (_25091_, _12242_, _05557_);
  nor (_25092_, _25091_, _25090_);
  not (_25094_, _25092_);
  nor (_25095_, _25094_, _25089_);
  nor (_25096_, _06912_, _05958_);
  and (_25097_, _12237_, _05977_);
  not (_25098_, _25097_);
  nor (_25099_, _25098_, _25096_);
  not (_25100_, _25099_);
  nor (_25101_, _25100_, _25095_);
  nor (_25102_, _25097_, _05557_);
  nor (_25103_, _25102_, _05970_);
  not (_25105_, _25103_);
  nor (_25106_, _25105_, _25101_);
  nor (_25107_, _06369_, _05968_);
  and (_25108_, _25107_, _12611_);
  not (_25109_, _25108_);
  or (_25110_, _25109_, _25106_);
  nor (_25111_, _25110_, _24999_);
  nor (_25112_, _25108_, _05557_);
  nor (_25113_, _25112_, _05900_);
  not (_25114_, _25113_);
  nor (_25116_, _25114_, _25111_);
  not (_25117_, _05900_);
  nor (_25118_, _06912_, _25117_);
  or (_25119_, _25118_, _12619_);
  nor (_25120_, _25119_, _25116_);
  nor (_25121_, _25028_, _12620_);
  nor (_25122_, _25121_, _25120_);
  and (_25123_, _25122_, _07198_);
  or (_25124_, _25123_, _24998_);
  and (_25125_, _25124_, _12635_);
  and (_25127_, _12634_, _06006_);
  or (_25128_, _25127_, _25125_);
  and (_25129_, _25128_, _13846_);
  nor (_25130_, _06912_, _13846_);
  or (_25131_, _25130_, _25129_);
  and (_25132_, _25131_, _12678_);
  not (_25133_, _24996_);
  nor (_25134_, _25028_, _11291_);
  and (_25135_, _11291_, _05557_);
  nor (_25136_, _25135_, _12678_);
  not (_25138_, _25136_);
  nor (_25139_, _25138_, _25134_);
  nor (_25140_, _25139_, _25133_);
  not (_25141_, _25140_);
  nor (_25142_, _25141_, _25132_);
  nor (_25143_, _25142_, _24997_);
  and (_25144_, _25143_, _05890_);
  nor (_25145_, _06912_, _05890_);
  or (_25146_, _25145_, _25144_);
  and (_25147_, _25146_, _12702_);
  not (_25149_, _24993_);
  nor (_25150_, _11291_, _05557_);
  and (_25151_, _25028_, _11291_);
  or (_25152_, _25151_, _25150_);
  and (_25153_, _25152_, _12701_);
  nor (_25154_, _25153_, _25149_);
  not (_25155_, _25154_);
  nor (_25156_, _25155_, _25147_);
  nor (_25157_, _25156_, _24995_);
  and (_25158_, _25157_, _05919_);
  nor (_25160_, _06912_, _05919_);
  or (_25161_, _25160_, _25158_);
  and (_25162_, _25161_, _12724_);
  not (_25163_, _24987_);
  or (_25164_, _25163_, _25162_);
  nor (_25165_, _25164_, _24992_);
  or (_25166_, _25165_, _12746_);
  nor (_25167_, _25166_, _24988_);
  nor (_25168_, _25167_, _24986_);
  nor (_25169_, _25168_, _12215_);
  and (_25171_, _10849_, \oc8051_golden_model_1.PC [0]);
  nor (_25172_, _10849_, \oc8051_golden_model_1.PC [0]);
  nor (_25173_, _25172_, _25171_);
  and (_25174_, _25173_, _12215_);
  nor (_25175_, _25174_, _25169_);
  and (_25176_, _25175_, _24984_);
  or (_25177_, _25176_, _06547_);
  nor (_25178_, _25177_, _24985_);
  and (_25179_, _09342_, _06547_);
  or (_25180_, _25179_, _25178_);
  and (_25182_, _25180_, _05916_);
  nor (_25183_, _06912_, _05916_);
  or (_25184_, _25183_, _25182_);
  and (_25185_, _25184_, _06946_);
  and (_25186_, _25001_, _12954_);
  nor (_25187_, _12954_, _05557_);
  or (_25188_, _25187_, _06946_);
  or (_25189_, _25188_, _25186_);
  and (_25190_, _25189_, _24981_);
  not (_25191_, _25190_);
  nor (_25193_, _25191_, _25185_);
  nor (_25194_, _25193_, _24982_);
  and (_25195_, _25194_, _06261_);
  and (_25196_, _09342_, _06260_);
  or (_25197_, _25196_, _25195_);
  and (_25198_, _25197_, _05924_);
  nor (_25199_, _06912_, _05924_);
  nor (_25200_, _25199_, _25198_);
  nor (_25201_, _25200_, _06377_);
  not (_25202_, _24979_);
  and (_25204_, _24977_, _06377_);
  nor (_25205_, _25204_, _25202_);
  not (_25206_, _25205_);
  nor (_25207_, _25206_, _25201_);
  nor (_25208_, _25207_, _24980_);
  nor (_25209_, _25208_, _07812_);
  and (_25210_, _07812_, _06912_);
  nor (_25211_, _25210_, _06199_);
  not (_25212_, _25211_);
  nor (_25213_, _25212_, _25209_);
  nor (_25215_, _25213_, _24978_);
  and (_25216_, _13006_, _13013_);
  not (_25217_, _25216_);
  nor (_25218_, _25217_, _25215_);
  nor (_25219_, _06342_, _05907_);
  not (_25220_, _25219_);
  nor (_25221_, _25216_, \oc8051_golden_model_1.PC [0]);
  nor (_25222_, _25221_, _25220_);
  not (_25223_, _25222_);
  nor (_25224_, _25223_, _25218_);
  and (_25226_, _25220_, _06912_);
  nor (_25227_, _25226_, _13025_);
  not (_25228_, _25227_);
  nor (_25229_, _25228_, _25224_);
  nor (_25230_, _25229_, _24971_);
  nand (_25231_, _25230_, _01452_);
  or (_25232_, _01452_, \oc8051_golden_model_1.PC [0]);
  and (_25233_, _25232_, _43223_);
  and (_43854_, _25233_, _25231_);
  nor (_25234_, _13013_, _05978_);
  nor (_25236_, _12991_, _05978_);
  nor (_25237_, _09012_, _05978_);
  nor (_25238_, _12105_, _05978_);
  and (_25239_, _10525_, _05938_);
  nor (_25240_, _12736_, _05978_);
  nor (_25241_, _12226_, _05978_);
  nor (_25242_, _12228_, _05550_);
  nor (_25243_, _17747_, _18386_);
  and (_25244_, _25243_, _17189_);
  and (_25245_, _25244_, _10917_);
  nor (_25247_, _25245_, _05978_);
  nor (_25248_, _08972_, _05550_);
  and (_25249_, _14150_, _05938_);
  and (_25250_, _12245_, _05938_);
  and (_25251_, _12513_, _05938_);
  nor (_25252_, _12314_, _12312_);
  nor (_25253_, _25252_, _12315_);
  not (_25254_, _25253_);
  nor (_25255_, _25254_, _12513_);
  or (_25256_, _25255_, _25251_);
  nor (_25258_, _25256_, _12478_);
  nor (_25259_, _12462_, _05978_);
  and (_25260_, _07134_, _05978_);
  not (_25261_, _25260_);
  not (_25262_, _12426_);
  nor (_25263_, _10704_, _05978_);
  nor (_25264_, _07018_, _07272_);
  nor (_25265_, _12419_, _05557_);
  nor (_25266_, _25265_, _07123_);
  and (_25267_, _25266_, _05550_);
  nor (_25269_, _25266_, _05550_);
  nor (_25270_, _25269_, _25267_);
  nor (_25271_, _25270_, _06808_);
  and (_25272_, _06808_, _05938_);
  nor (_25273_, _25272_, _25271_);
  and (_25274_, _25273_, _07272_);
  nor (_25275_, _25274_, _17204_);
  not (_25276_, _25275_);
  nor (_25277_, _25276_, _25264_);
  nor (_25278_, _25277_, _25263_);
  nor (_25280_, _25278_, _25262_);
  nor (_25281_, _12426_, _05978_);
  nor (_25282_, _25281_, _08572_);
  not (_25283_, _25282_);
  nor (_25284_, _25283_, _25280_);
  or (_25285_, _12414_, _05550_);
  nor (_25286_, _12162_, _12160_);
  nor (_25287_, _25286_, _12163_);
  or (_25288_, _25287_, _12412_);
  and (_25289_, _25288_, _08572_);
  and (_25291_, _25289_, _25285_);
  or (_25292_, _25291_, _25284_);
  nand (_25293_, _25292_, _07338_);
  and (_25294_, _25293_, _25261_);
  or (_25295_, _25294_, _06251_);
  or (_25296_, _25254_, _12402_);
  or (_25297_, _12404_, _05978_);
  and (_25298_, _25297_, _25296_);
  or (_25299_, _25298_, _06252_);
  and (_25300_, _25299_, _12443_);
  nand (_25301_, _25300_, _25295_);
  nor (_25302_, _12443_, _05978_);
  nor (_25303_, _25302_, _06475_);
  nand (_25304_, _25303_, _25301_);
  and (_25305_, _06475_, _05550_);
  nor (_25306_, _25305_, _07474_);
  nand (_25307_, _25306_, _25304_);
  and (_25308_, _07018_, _07474_);
  nor (_25309_, _25308_, _06468_);
  nand (_25310_, _25309_, _25307_);
  and (_25313_, _06468_, _05550_);
  nor (_25314_, _25313_, _12452_);
  nand (_25315_, _25314_, _25310_);
  nor (_25316_, _12451_, _05978_);
  nor (_25317_, _25316_, _06466_);
  nand (_25318_, _25317_, _25315_);
  and (_25319_, _06466_, _05550_);
  nor (_25320_, _25319_, _12464_);
  and (_25321_, _25320_, _25318_);
  or (_25322_, _25321_, _25259_);
  nand (_25324_, _25322_, _06484_);
  and (_25325_, _06483_, \oc8051_golden_model_1.PC [1]);
  nor (_25326_, _25325_, _12466_);
  and (_25327_, _25326_, _25324_);
  nor (_25328_, _07018_, _05953_);
  or (_25329_, _25328_, _25327_);
  nand (_25330_, _25329_, _07523_);
  and (_25331_, _06247_, _05550_);
  nor (_25332_, _25331_, _12479_);
  and (_25333_, _25332_, _25330_);
  or (_25335_, _25333_, _25258_);
  nand (_25336_, _25335_, _06345_);
  nand (_25337_, _12392_, _05938_);
  or (_25338_, _25254_, _12392_);
  and (_25339_, _25338_, _06344_);
  nand (_25340_, _25339_, _25337_);
  and (_25341_, _25340_, _12536_);
  nand (_25342_, _25341_, _25336_);
  and (_25343_, _12533_, _05978_);
  nor (_25344_, _25253_, _12533_);
  or (_25346_, _25344_, _12536_);
  or (_25347_, _25346_, _25343_);
  nand (_25348_, _25347_, _25342_);
  nand (_25349_, _25348_, _12522_);
  and (_25350_, _12555_, _05938_);
  nor (_25351_, _25254_, _12555_);
  or (_25352_, _25351_, _25350_);
  and (_25353_, _25352_, _06373_);
  nor (_25354_, _25353_, _12245_);
  and (_25355_, _25354_, _25349_);
  or (_25357_, _25355_, _25250_);
  nand (_25358_, _25357_, _07164_);
  and (_25359_, _06461_, \oc8051_golden_model_1.PC [1]);
  nor (_25360_, _25359_, _07471_);
  nand (_25361_, _25360_, _25358_);
  nor (_25362_, _07018_, _05947_);
  nor (_25363_, _06194_, _06358_);
  or (_25364_, _25363_, _05957_);
  and (_25365_, _25364_, _12568_);
  not (_25366_, _25365_);
  nor (_25368_, _25366_, _25362_);
  nand (_25369_, _25368_, _25361_);
  nor (_25370_, _25365_, _05550_);
  nor (_25371_, _25370_, _12239_);
  and (_25372_, _25371_, _25369_);
  and (_25373_, _12241_, _05938_);
  nor (_25374_, _25373_, _12242_);
  or (_25375_, _25374_, _25372_);
  nor (_25376_, _12241_, _05978_);
  nor (_25377_, _25376_, _06505_);
  nand (_25379_, _25377_, _25375_);
  and (_25380_, _06505_, _05550_);
  nor (_25381_, _25380_, _25090_);
  nand (_25382_, _25381_, _25379_);
  and (_25383_, _07018_, _25090_);
  nor (_25384_, _25383_, _06504_);
  nand (_25385_, _25384_, _25382_);
  and (_25386_, _06504_, _05550_);
  nor (_25387_, _25386_, _14150_);
  and (_25388_, _25387_, _25385_);
  or (_25390_, _25388_, _25249_);
  and (_25391_, _07129_, _05969_);
  nor (_25392_, _17815_, _25391_);
  nand (_25393_, _25392_, _25390_);
  nor (_25394_, _25392_, _05978_);
  nor (_25395_, _25394_, _17755_);
  nand (_25396_, _25395_, _25393_);
  and (_25397_, _17755_, _05978_);
  nor (_25398_, _25397_, _12589_);
  nand (_25399_, _25398_, _25396_);
  nor (_25401_, _12588_, _05550_);
  nor (_25402_, _25401_, _05976_);
  nand (_25403_, _25402_, _25399_);
  and (_25404_, _05976_, _05978_);
  nor (_25405_, _25404_, _06241_);
  and (_25406_, _25405_, _25403_);
  and (_25407_, _06241_, \oc8051_golden_model_1.PC [1]);
  or (_25408_, _25407_, _25406_);
  nand (_25409_, _25408_, _08723_);
  and (_25410_, _07018_, _05970_);
  nor (_25412_, _25410_, _06369_);
  nand (_25413_, _25412_, _25409_);
  and (_25414_, _06369_, _05938_);
  nor (_25415_, _25414_, _12604_);
  nand (_25416_, _25415_, _25413_);
  nor (_25417_, _12603_, _05550_);
  nor (_25418_, _25417_, _05968_);
  nand (_25419_, _25418_, _25416_);
  and (_25420_, _05968_, _05938_);
  nor (_25421_, _25420_, _12615_);
  nand (_25423_, _25421_, _25419_);
  nor (_25424_, _12611_, _05978_);
  nor (_25425_, _25424_, _06332_);
  nand (_25426_, _25425_, _25423_);
  and (_25427_, _06332_, _05550_);
  nor (_25428_, _25427_, _05900_);
  nand (_25429_, _25428_, _25426_);
  and (_25430_, _07018_, _05900_);
  nor (_25431_, _25430_, _12619_);
  nand (_25432_, _25431_, _25429_);
  and (_25434_, _25287_, _12619_);
  nor (_25435_, _25434_, _08973_);
  and (_25436_, _25435_, _25432_);
  or (_25437_, _25436_, _25248_);
  nand (_25438_, _25437_, _07198_);
  and (_25439_, _06371_, _05978_);
  nor (_25440_, _25439_, _10904_);
  nand (_25441_, _25440_, _25438_);
  and (_25442_, _10904_, _05550_);
  nor (_25443_, _25442_, _12634_);
  nand (_25445_, _25443_, _25441_);
  nor (_25446_, _12635_, _05987_);
  nor (_25447_, _25446_, _06331_);
  nand (_25448_, _25447_, _25445_);
  and (_25449_, _06331_, _05550_);
  nor (_25450_, _25449_, _05895_);
  nand (_25451_, _25450_, _25448_);
  and (_25452_, _07018_, _05895_);
  nor (_25453_, _25452_, _12677_);
  nand (_25454_, _25453_, _25451_);
  not (_25456_, _25245_);
  and (_25457_, _11291_, _05550_);
  and (_25458_, _25287_, _12684_);
  or (_25459_, _25458_, _25457_);
  and (_25460_, _25459_, _12677_);
  nor (_25461_, _25460_, _25456_);
  and (_25462_, _25461_, _25454_);
  or (_25463_, _25462_, _25247_);
  nor (_25464_, _18236_, _17915_);
  nand (_25465_, _25464_, _25463_);
  nor (_25467_, _25464_, _05978_);
  nor (_25468_, _25467_, _18067_);
  nand (_25469_, _25468_, _25465_);
  and (_25470_, _18067_, _05978_);
  nor (_25471_, _25470_, _12229_);
  and (_25472_, _25471_, _25469_);
  or (_25473_, _25472_, _25242_);
  nand (_25474_, _25473_, _07218_);
  and (_25475_, _06367_, _05978_);
  nor (_25476_, _25475_, _06533_);
  nand (_25478_, _25476_, _25474_);
  and (_25479_, _06533_, _05550_);
  nor (_25480_, _25479_, _05889_);
  nand (_25481_, _25480_, _25478_);
  and (_25482_, _07018_, _05889_);
  nor (_25483_, _25482_, _12701_);
  nand (_25484_, _25483_, _25481_);
  nor (_25485_, _25287_, _12684_);
  nor (_25486_, _11291_, _05550_);
  nor (_25487_, _25486_, _12702_);
  not (_25489_, _25487_);
  nor (_25490_, _25489_, _25485_);
  nor (_25491_, _25490_, _12710_);
  and (_25492_, _25491_, _25484_);
  or (_25493_, _25492_, _25241_);
  nand (_25494_, _25493_, _10967_);
  nor (_25495_, _10967_, _05550_);
  nor (_25496_, _25495_, _06366_);
  nand (_25497_, _25496_, _25494_);
  and (_25498_, _06366_, _05938_);
  nor (_25500_, _25498_, _06541_);
  and (_25501_, _25500_, _25497_);
  and (_25502_, _06541_, \oc8051_golden_model_1.PC [1]);
  or (_25503_, _25502_, _25501_);
  nand (_25504_, _25503_, _05919_);
  and (_25505_, _07018_, _07209_);
  nor (_25506_, _25505_, _12723_);
  nand (_25507_, _25506_, _25504_);
  nor (_25508_, _25287_, \oc8051_golden_model_1.PSW [7]);
  and (_25509_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor (_25511_, _25509_, _12724_);
  not (_25512_, _25511_);
  nor (_25513_, _25512_, _25508_);
  nor (_25514_, _25513_, _12738_);
  and (_25515_, _25514_, _25507_);
  or (_25516_, _25515_, _25240_);
  nand (_25517_, _25516_, _11005_);
  nor (_25518_, _11005_, _05550_);
  nor (_25519_, _25518_, _06383_);
  nand (_25520_, _25519_, _25517_);
  and (_25522_, _06383_, _05938_);
  nor (_25523_, _25522_, _06528_);
  and (_25524_, _25523_, _25520_);
  and (_25525_, _06528_, \oc8051_golden_model_1.PC [1]);
  or (_25526_, _25525_, _25524_);
  nand (_25527_, _25526_, _05922_);
  and (_25528_, _07018_, _12746_);
  nor (_25529_, _25528_, _12215_);
  nand (_25530_, _25529_, _25527_);
  nor (_25531_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_25533_, _25287_, \oc8051_golden_model_1.PSW [7]);
  or (_25534_, _25533_, _25531_);
  and (_25535_, _25534_, _12215_);
  nor (_25536_, _25535_, _10525_);
  and (_25537_, _25536_, _25530_);
  or (_25538_, _25537_, _25239_);
  nand (_25539_, _25538_, _17668_);
  nor (_25540_, _17668_, _05978_);
  nor (_25541_, _25540_, _17673_);
  nand (_25542_, _25541_, _25539_);
  and (_25544_, _17673_, _05978_);
  nor (_25545_, _25544_, _11052_);
  nand (_25546_, _25545_, _25542_);
  nor (_25547_, _11051_, _05550_);
  nor (_25548_, _25547_, _11080_);
  nand (_25549_, _25548_, _25546_);
  and (_25550_, _11080_, _05978_);
  nor (_25551_, _25550_, _06547_);
  and (_25552_, _25551_, _25549_);
  nor (_25553_, _09297_, _13873_);
  or (_25555_, _25553_, _25552_);
  nand (_25556_, _25555_, _05916_);
  and (_25557_, _07018_, _07228_);
  nor (_25558_, _25557_, _06381_);
  nand (_25559_, _25558_, _25556_);
  and (_25560_, _25254_, _12954_);
  not (_25561_, _25560_);
  nor (_25562_, _12954_, _05938_);
  nor (_25563_, _25562_, _06946_);
  and (_25564_, _25563_, _25561_);
  nor (_25566_, _25564_, _12774_);
  and (_25567_, _25566_, _25559_);
  or (_25568_, _25567_, _25238_);
  nand (_25569_, _25568_, _12963_);
  nor (_25570_, _12963_, _05550_);
  nor (_25571_, _25570_, _10448_);
  nand (_25572_, _25571_, _25569_);
  and (_25573_, _10448_, _05978_);
  nor (_25574_, _25573_, _06260_);
  and (_25575_, _25574_, _25572_);
  nor (_25577_, _09297_, _06261_);
  or (_25578_, _25577_, _25575_);
  nand (_25579_, _25578_, _05924_);
  and (_25580_, _07018_, _12089_);
  nor (_25581_, _25580_, _06377_);
  nand (_25582_, _25581_, _25579_);
  and (_25583_, _12954_, _05978_);
  nor (_25584_, _25253_, _12954_);
  nor (_25585_, _25584_, _25583_);
  and (_25586_, _25585_, _06377_);
  nor (_25588_, _25586_, _15238_);
  and (_25589_, _25588_, _25582_);
  or (_25590_, _25589_, _25237_);
  nor (_25591_, _07238_, _07243_);
  nand (_25592_, _25591_, _25590_);
  nor (_25593_, _25591_, _05978_);
  nor (_25594_, _25593_, _06563_);
  nand (_25595_, _25594_, _25592_);
  and (_25596_, _06563_, _05550_);
  nor (_25597_, _25596_, _12992_);
  and (_25599_, _25597_, _25595_);
  or (_25600_, _25599_, _25236_);
  nand (_25601_, _25600_, _07250_);
  and (_25602_, _07812_, _07018_);
  nor (_25603_, _25602_, _06199_);
  nand (_25604_, _25603_, _25601_);
  not (_25605_, _14678_);
  and (_25606_, _25585_, _06199_);
  nor (_25607_, _25606_, _25605_);
  and (_25608_, _25607_, _25604_);
  nor (_25609_, _14678_, _05978_);
  or (_25610_, _25609_, _25608_);
  nor (_25611_, _07256_, _07259_);
  nand (_25612_, _25611_, _25610_);
  nor (_25613_, _25611_, _05978_);
  nor (_25614_, _25613_, _06188_);
  nand (_25615_, _25614_, _25612_);
  and (_25616_, _06188_, _05550_);
  nor (_25617_, _25616_, _13014_);
  and (_25618_, _25617_, _25615_);
  or (_25621_, _25618_, _25234_);
  nand (_25622_, _25621_, _25219_);
  and (_25623_, _25220_, _07018_);
  nor (_25624_, _25623_, _13025_);
  and (_25625_, _25624_, _25622_);
  and (_25626_, _13025_, _05978_);
  or (_25627_, _25626_, _25625_);
  or (_25628_, _25627_, _01456_);
  or (_25629_, _01452_, \oc8051_golden_model_1.PC [1]);
  and (_25630_, _25629_, _43223_);
  and (_43855_, _25630_, _25628_);
  and (_25632_, _06188_, _06018_);
  and (_25633_, _06563_, _06018_);
  nor (_25634_, _09251_, _06261_);
  nor (_25635_, _12105_, _06024_);
  nor (_25636_, _12756_, _06024_);
  nor (_25637_, _12736_, _06024_);
  nor (_25638_, _12226_, _06024_);
  nor (_25639_, _12232_, _06024_);
  nand (_25640_, _05899_, _06192_);
  not (_25642_, _25640_);
  and (_25643_, _07490_, _08581_);
  nor (_25644_, _25643_, _25642_);
  nor (_25645_, _25644_, _06018_);
  not (_25646_, _06024_);
  and (_25647_, _12245_, _25646_);
  and (_25648_, _06651_, _06705_);
  nor (_25649_, _12427_, _06024_);
  or (_25650_, _12419_, _25646_);
  nand (_25651_, _12420_, \oc8051_golden_model_1.PC [2]);
  and (_25653_, _25651_, _25650_);
  or (_25654_, _25653_, _07123_);
  and (_25655_, _06808_, _06024_);
  nor (_25656_, _06808_, _06019_);
  and (_25657_, _25656_, _07123_);
  nor (_25658_, _25657_, _25655_);
  and (_25659_, _25658_, _25018_);
  and (_25660_, _25659_, _25654_);
  or (_25661_, _25660_, _25649_);
  nor (_25662_, _25661_, _25648_);
  nor (_25664_, _25662_, _08572_);
  or (_25665_, _12414_, _06019_);
  and (_25666_, _12167_, _12164_);
  nor (_25667_, _25666_, _12168_);
  nand (_25668_, _25667_, _12414_);
  and (_25669_, _25668_, _08572_);
  and (_25670_, _25669_, _25665_);
  or (_25671_, _25670_, _25664_);
  nand (_25672_, _25671_, _07338_);
  and (_25673_, _07134_, _25646_);
  nor (_25675_, _25673_, _06251_);
  nand (_25676_, _25675_, _25672_);
  and (_25677_, _12319_, _12316_);
  nor (_25678_, _25677_, _12320_);
  or (_25679_, _25678_, _12402_);
  or (_25680_, _12404_, _12308_);
  and (_25681_, _25680_, _06251_);
  nand (_25682_, _25681_, _25679_);
  and (_25683_, _25682_, _12443_);
  nand (_25684_, _25683_, _25676_);
  nor (_25686_, _12443_, _06024_);
  nor (_25687_, _25686_, _06475_);
  nand (_25688_, _25687_, _25684_);
  and (_25689_, _06475_, _06018_);
  nor (_25690_, _25689_, _07474_);
  nand (_25691_, _25690_, _25688_);
  and (_25692_, _06651_, _07474_);
  nor (_25693_, _25692_, _06468_);
  nand (_25694_, _25693_, _25691_);
  and (_25695_, _06468_, _06018_);
  nor (_25697_, _25695_, _12452_);
  nand (_25698_, _25697_, _25694_);
  nor (_25699_, _12451_, _06024_);
  nor (_25700_, _25699_, _06466_);
  nand (_25701_, _25700_, _25698_);
  and (_25702_, _06466_, _06018_);
  nor (_25703_, _25702_, _12464_);
  nand (_25704_, _25703_, _25701_);
  nor (_25705_, _12462_, _06024_);
  nor (_25706_, _25705_, _06483_);
  nand (_25708_, _25706_, _25704_);
  and (_25709_, _06483_, _06018_);
  nor (_25710_, _25709_, _12466_);
  nand (_25711_, _25710_, _25708_);
  and (_25712_, _06651_, _12466_);
  nor (_25713_, _25712_, _06247_);
  nand (_25714_, _25713_, _25711_);
  and (_25715_, _06247_, _06018_);
  nor (_25716_, _25715_, _12479_);
  and (_25717_, _25716_, _25714_);
  nor (_25719_, _25678_, _12513_);
  and (_25720_, _12513_, _12309_);
  nor (_25721_, _25720_, _25719_);
  nor (_25722_, _25721_, _12478_);
  or (_25723_, _25722_, _25717_);
  nand (_25724_, _25723_, _06345_);
  not (_25725_, _25678_);
  or (_25726_, _25725_, _12392_);
  nand (_25727_, _12392_, _12308_);
  and (_25728_, _25727_, _06344_);
  nand (_25730_, _25728_, _25726_);
  nand (_25731_, _25730_, _25724_);
  nand (_25732_, _25731_, _12536_);
  and (_25733_, _12533_, _12308_);
  not (_25734_, _25733_);
  nor (_25735_, _25725_, _12533_);
  nor (_25736_, _25735_, _12536_);
  and (_25737_, _25736_, _25734_);
  nor (_25738_, _25737_, _06373_);
  nand (_25739_, _25738_, _25732_);
  and (_25741_, _12555_, _12309_);
  nor (_25742_, _25678_, _12555_);
  or (_25743_, _25742_, _12522_);
  or (_25744_, _25743_, _25741_);
  and (_25745_, _25744_, _12246_);
  and (_25746_, _25745_, _25739_);
  or (_25747_, _25746_, _25647_);
  nand (_25748_, _25747_, _07164_);
  and (_25749_, _06461_, _06019_);
  nor (_25750_, _25749_, _07471_);
  nand (_25752_, _25750_, _25748_);
  nor (_25753_, _06651_, _05947_);
  nor (_25754_, _25753_, _25366_);
  and (_25755_, _25754_, _25752_);
  nor (_25756_, _25365_, _06018_);
  or (_25757_, _25756_, _25755_);
  nand (_25758_, _25757_, _12242_);
  nor (_25759_, _12242_, _06024_);
  nor (_25760_, _25759_, _06505_);
  nand (_25761_, _25760_, _25758_);
  and (_25763_, _06505_, _06018_);
  nor (_25764_, _25763_, _25090_);
  nand (_25765_, _25764_, _25761_);
  and (_25766_, _06651_, _25090_);
  nor (_25767_, _25766_, _06504_);
  nand (_25768_, _25767_, _25765_);
  and (_25769_, _06504_, _06018_);
  nor (_25770_, _25769_, _12582_);
  and (_25771_, _25770_, _25768_);
  nor (_25772_, _12237_, _06024_);
  or (_25774_, _25772_, _25771_);
  nand (_25775_, _25774_, _12588_);
  nor (_25776_, _12588_, _06018_);
  nor (_25777_, _25776_, _05976_);
  nand (_25778_, _25777_, _25775_);
  and (_25779_, _06024_, _05976_);
  nor (_25780_, _25779_, _06241_);
  and (_25781_, _25780_, _25778_);
  and (_25782_, _06241_, _06019_);
  or (_25783_, _25782_, _25781_);
  nand (_25785_, _25783_, _08723_);
  and (_25786_, _06651_, _05970_);
  nor (_25787_, _25786_, _06369_);
  nand (_25788_, _25787_, _25785_);
  and (_25789_, _12308_, _06369_);
  not (_25790_, _25789_);
  and (_25791_, _25790_, _25644_);
  and (_25792_, _25791_, _25788_);
  or (_25793_, _25792_, _25645_);
  and (_25794_, _05899_, _06348_);
  nor (_25796_, _07182_, _25794_);
  nand (_25797_, _25796_, _25793_);
  nor (_25798_, _25796_, _06018_);
  nor (_25799_, _25798_, _05968_);
  nand (_25800_, _25799_, _25797_);
  and (_25801_, _12308_, _05968_);
  nor (_25802_, _25801_, _12615_);
  nand (_25803_, _25802_, _25800_);
  nor (_25804_, _12611_, _06024_);
  nor (_25805_, _25804_, _06332_);
  and (_25807_, _25805_, _25803_);
  and (_25808_, _06332_, _06018_);
  or (_25809_, _25808_, _05900_);
  nor (_25810_, _25809_, _25807_);
  and (_25811_, _06651_, _05900_);
  or (_25812_, _25811_, _25810_);
  nand (_25813_, _25812_, _12620_);
  nor (_25814_, _25667_, _12620_);
  nor (_25815_, _25814_, _08968_);
  nand (_25816_, _25815_, _25813_);
  and (_25818_, _08968_, _06018_);
  not (_25819_, _25818_);
  nand (_25820_, _07438_, _05932_);
  and (_25821_, _25820_, _07460_);
  and (_25822_, _25821_, _25819_);
  nand (_25823_, _25822_, _25816_);
  nor (_25824_, _25821_, _06018_);
  and (_25825_, _05894_, _06817_);
  not (_25826_, _25825_);
  not (_25827_, _05894_);
  nor (_25829_, _07129_, _07455_);
  nor (_25830_, _25829_, _25827_);
  nor (_25831_, _25830_, _06916_);
  nand (_25832_, _25831_, _25826_);
  nor (_25833_, _25832_, _25824_);
  and (_25834_, _25833_, _25823_);
  and (_25835_, _25832_, _06018_);
  or (_25836_, _25835_, _06371_);
  or (_25837_, _25836_, _25834_);
  and (_25838_, _12309_, _06371_);
  nor (_25840_, _25838_, _10904_);
  nand (_25841_, _25840_, _25837_);
  and (_25842_, _10904_, _06018_);
  nor (_25843_, _25842_, _12634_);
  nand (_25844_, _25843_, _25841_);
  and (_25845_, _12634_, _06035_);
  nor (_25846_, _25845_, _06331_);
  and (_25847_, _25846_, _25844_);
  and (_25848_, _06331_, _06018_);
  or (_25849_, _25848_, _05895_);
  or (_25851_, _25849_, _25847_);
  and (_25852_, _06651_, _05895_);
  nor (_25853_, _25852_, _12677_);
  nand (_25854_, _25853_, _25851_);
  nor (_25855_, _25667_, _11291_);
  and (_25856_, _11291_, _06019_);
  nor (_25857_, _25856_, _12678_);
  not (_25858_, _25857_);
  nor (_25859_, _25858_, _25855_);
  nor (_25860_, _25859_, _12682_);
  and (_25862_, _25860_, _25854_);
  or (_25863_, _25862_, _25639_);
  nand (_25864_, _25863_, _12228_);
  nor (_25865_, _12228_, _06018_);
  nor (_25866_, _25865_, _06367_);
  and (_25867_, _25866_, _25864_);
  and (_25868_, _12308_, _06367_);
  or (_25869_, _25868_, _06533_);
  nor (_25870_, _25869_, _25867_);
  and (_25871_, _06533_, _06019_);
  or (_25873_, _25871_, _25870_);
  nand (_25874_, _25873_, _05890_);
  and (_25875_, _06651_, _05889_);
  nor (_25876_, _25875_, _12701_);
  nand (_25877_, _25876_, _25874_);
  nor (_25878_, _11291_, _06019_);
  and (_25879_, _25667_, _11291_);
  or (_25880_, _25879_, _25878_);
  and (_25881_, _25880_, _12701_);
  nor (_25882_, _25881_, _12710_);
  and (_25884_, _25882_, _25877_);
  or (_25885_, _25884_, _25638_);
  nand (_25886_, _25885_, _10967_);
  nor (_25887_, _10967_, _06018_);
  nor (_25888_, _25887_, _06366_);
  nand (_25889_, _25888_, _25886_);
  and (_25890_, _12308_, _06366_);
  nor (_25891_, _25890_, _06541_);
  and (_25892_, _25891_, _25889_);
  and (_25893_, _06541_, _06019_);
  or (_25895_, _25893_, _25892_);
  nand (_25896_, _25895_, _05919_);
  and (_25897_, _06651_, _07209_);
  nor (_25898_, _25897_, _12723_);
  nand (_25899_, _25898_, _25896_);
  nor (_25900_, _25667_, \oc8051_golden_model_1.PSW [7]);
  nor (_25901_, _06018_, _10854_);
  nor (_25902_, _25901_, _12724_);
  not (_25903_, _25902_);
  nor (_25904_, _25903_, _25900_);
  nor (_25906_, _25904_, _12738_);
  and (_25907_, _25906_, _25899_);
  or (_25908_, _25907_, _25637_);
  nand (_25909_, _25908_, _11005_);
  nor (_25910_, _11005_, _06018_);
  nor (_25911_, _25910_, _06383_);
  and (_25912_, _25911_, _25909_);
  and (_25913_, _12308_, _06383_);
  or (_25914_, _25913_, _06528_);
  nor (_25915_, _25914_, _25912_);
  and (_25917_, _06528_, _06019_);
  or (_25918_, _25917_, _25915_);
  nand (_25919_, _25918_, _05922_);
  and (_25920_, _06651_, _12746_);
  nor (_25921_, _25920_, _12215_);
  nand (_25922_, _25921_, _25919_);
  nor (_25923_, _25667_, _10854_);
  nor (_25924_, _06018_, \oc8051_golden_model_1.PSW [7]);
  nor (_25925_, _25924_, _12751_);
  not (_25926_, _25925_);
  nor (_25928_, _25926_, _25923_);
  nor (_25929_, _25928_, _12758_);
  and (_25930_, _25929_, _25922_);
  or (_25931_, _25930_, _25636_);
  nand (_25932_, _25931_, _11051_);
  nor (_25933_, _11051_, _06018_);
  nor (_25934_, _25933_, _11080_);
  nand (_25935_, _25934_, _25932_);
  and (_25936_, _11080_, _06024_);
  nor (_25937_, _25936_, _06547_);
  and (_25938_, _25937_, _25935_);
  nor (_25939_, _09251_, _13873_);
  or (_25940_, _25939_, _25938_);
  nand (_25941_, _25940_, _05916_);
  and (_25942_, _06651_, _07228_);
  nor (_25943_, _25942_, _06381_);
  nand (_25944_, _25943_, _25941_);
  and (_25945_, _25725_, _12954_);
  nor (_25946_, _12308_, _12954_);
  or (_25947_, _25946_, _06946_);
  or (_25950_, _25947_, _25945_);
  and (_25951_, _25950_, _12105_);
  and (_25952_, _25951_, _25944_);
  or (_25953_, _25952_, _25635_);
  nand (_25954_, _25953_, _12963_);
  nor (_25955_, _12963_, _06018_);
  nor (_25956_, _25955_, _10448_);
  nand (_25957_, _25956_, _25954_);
  and (_25958_, _10448_, _06024_);
  nor (_25959_, _25958_, _06260_);
  and (_25961_, _25959_, _25957_);
  or (_25962_, _25961_, _25634_);
  nand (_25963_, _25962_, _05924_);
  and (_25964_, _06651_, _12089_);
  nor (_25965_, _25964_, _06377_);
  nand (_25966_, _25965_, _25963_);
  nor (_25967_, _25678_, _12954_);
  and (_25968_, _12309_, _12954_);
  nor (_25969_, _25968_, _25967_);
  and (_25970_, _25969_, _06377_);
  nor (_25972_, _25970_, _12985_);
  nand (_25973_, _25972_, _25966_);
  nor (_25974_, _12984_, _06024_);
  nor (_25975_, _25974_, _06563_);
  and (_25976_, _25975_, _25973_);
  or (_25977_, _25976_, _25633_);
  nand (_25978_, _25977_, _12991_);
  nor (_25979_, _12991_, _25646_);
  nor (_25980_, _25979_, _07812_);
  nand (_25981_, _25980_, _25978_);
  and (_25983_, _07812_, _06651_);
  nor (_25984_, _25983_, _06199_);
  nand (_25985_, _25984_, _25981_);
  and (_25986_, _25969_, _06199_);
  nor (_25987_, _25986_, _13007_);
  nand (_25988_, _25987_, _25985_);
  nor (_25989_, _13006_, _06024_);
  nor (_25990_, _25989_, _06188_);
  and (_25991_, _25990_, _25988_);
  or (_25992_, _25991_, _25632_);
  nand (_25994_, _25992_, _13013_);
  nor (_25995_, _13013_, _25646_);
  nor (_25996_, _25995_, _25220_);
  nand (_25997_, _25996_, _25994_);
  and (_25998_, _25220_, _06651_);
  nor (_25999_, _25998_, _13025_);
  and (_26000_, _25999_, _25997_);
  and (_26001_, _13025_, _06024_);
  or (_26002_, _26001_, _26000_);
  or (_26003_, _26002_, _01456_);
  or (_26005_, _01452_, \oc8051_golden_model_1.PC [2]);
  and (_26006_, _26005_, _43223_);
  and (_43856_, _26006_, _26003_);
  and (_26007_, _06188_, _06075_);
  and (_26008_, _06563_, _06075_);
  nor (_26009_, _12105_, _06071_);
  nor (_26010_, _12756_, _06071_);
  nor (_26011_, _12736_, _06071_);
  nor (_26012_, _12226_, _06071_);
  nor (_26013_, _12232_, _06071_);
  nor (_26015_, _08972_, _06075_);
  and (_26016_, _06241_, _06095_);
  and (_26017_, _12245_, _06062_);
  or (_26018_, _12306_, _12305_);
  and (_26019_, _26018_, _12321_);
  nor (_26020_, _26018_, _12321_);
  nor (_26021_, _26020_, _26019_);
  not (_26022_, _26021_);
  nor (_26023_, _26022_, _12533_);
  and (_26024_, _12533_, _12303_);
  nor (_26026_, _26024_, _26023_);
  or (_26027_, _26026_, _12536_);
  nor (_26028_, _06458_, _07272_);
  and (_26029_, _07123_, _06095_);
  nor (_26030_, _26029_, _06808_);
  and (_26031_, _12419_, \oc8051_golden_model_1.PC [3]);
  or (_26032_, _26031_, _07123_);
  and (_26033_, _26032_, _26030_);
  or (_26034_, _12420_, _06062_);
  nand (_26035_, _26034_, _12427_);
  or (_26037_, _26035_, _26033_);
  and (_26038_, _26037_, _07272_);
  nor (_26039_, _26038_, _26028_);
  nor (_26040_, _12427_, _06071_);
  nor (_26041_, _26040_, _26039_);
  nor (_26042_, _26041_, _08572_);
  and (_26043_, _12412_, _06075_);
  not (_26044_, _26043_);
  or (_26045_, _12157_, _12156_);
  and (_26046_, _26045_, _12169_);
  nor (_26048_, _26045_, _12169_);
  nor (_26049_, _26048_, _26046_);
  and (_26050_, _26049_, _12414_);
  nor (_26051_, _26050_, _08573_);
  and (_26052_, _26051_, _26044_);
  nor (_26053_, _26052_, _26042_);
  nor (_26054_, _26053_, _07134_);
  and (_26055_, _07134_, _06062_);
  or (_26056_, _26055_, _26054_);
  or (_26057_, _26056_, _06251_);
  and (_26059_, _12402_, _12303_);
  and (_26060_, _26021_, _12404_);
  or (_26061_, _26060_, _26059_);
  and (_26062_, _26061_, _06251_);
  nor (_26063_, _26062_, _12444_);
  nand (_26064_, _26063_, _26057_);
  nor (_26065_, _12443_, _06071_);
  nor (_26066_, _26065_, _06475_);
  nand (_26067_, _26066_, _26064_);
  and (_26068_, _06475_, _06075_);
  nor (_26070_, _26068_, _07474_);
  nand (_26071_, _26070_, _26067_);
  and (_26072_, _06458_, _07474_);
  nor (_26073_, _26072_, _06468_);
  nand (_26074_, _26073_, _26071_);
  and (_26075_, _06468_, _06075_);
  nor (_26076_, _26075_, _12452_);
  nand (_26077_, _26076_, _26074_);
  nor (_26078_, _12451_, _06071_);
  nor (_26079_, _26078_, _06466_);
  nand (_26081_, _26079_, _26077_);
  and (_26082_, _06466_, _06075_);
  nor (_26083_, _26082_, _12464_);
  nand (_26084_, _26083_, _26081_);
  nor (_26085_, _12462_, _06071_);
  nor (_26086_, _26085_, _06483_);
  nand (_26087_, _26086_, _26084_);
  and (_26088_, _06483_, _06075_);
  nor (_26089_, _26088_, _12466_);
  nand (_26090_, _26089_, _26087_);
  and (_26092_, _06458_, _12466_);
  nor (_26093_, _26092_, _06247_);
  nand (_26094_, _26093_, _26090_);
  and (_26095_, _06247_, _06075_);
  nor (_26096_, _26095_, _12479_);
  and (_26097_, _26096_, _26094_);
  and (_26098_, _12513_, _12303_);
  nor (_26099_, _26022_, _12513_);
  or (_26100_, _26099_, _26098_);
  nor (_26101_, _26100_, _12478_);
  or (_26103_, _26101_, _26097_);
  and (_26104_, _26103_, _06345_);
  and (_26105_, _12392_, _12303_);
  nor (_26106_, _26022_, _12392_);
  or (_26107_, _26106_, _06345_);
  nor (_26108_, _26107_, _26105_);
  or (_26109_, _26108_, _26104_);
  or (_26110_, _26109_, _06338_);
  and (_26111_, _26110_, _26027_);
  or (_26112_, _26111_, _06373_);
  nor (_26114_, _26021_, _12555_);
  and (_26115_, _12555_, _12304_);
  or (_26116_, _26115_, _12522_);
  nor (_26117_, _26116_, _26114_);
  nor (_26118_, _26117_, _12245_);
  and (_26119_, _26118_, _26112_);
  or (_26120_, _26119_, _26017_);
  nand (_26121_, _26120_, _07164_);
  and (_26122_, _06461_, _06095_);
  nor (_26123_, _26122_, _07471_);
  nand (_26125_, _26123_, _26121_);
  nor (_26126_, _06458_, _05947_);
  nor (_26127_, _26126_, _25366_);
  and (_26128_, _26127_, _26125_);
  nor (_26129_, _25365_, _06075_);
  or (_26130_, _26129_, _26128_);
  nand (_26131_, _26130_, _12242_);
  nor (_26132_, _12242_, _06071_);
  nor (_26133_, _26132_, _06505_);
  nand (_26134_, _26133_, _26131_);
  and (_26136_, _06505_, _06075_);
  nor (_26137_, _26136_, _25090_);
  nand (_26138_, _26137_, _26134_);
  and (_26139_, _06458_, _25090_);
  nor (_26140_, _26139_, _06504_);
  nand (_26141_, _26140_, _26138_);
  and (_26142_, _06504_, _06075_);
  nor (_26143_, _26142_, _12582_);
  and (_26144_, _26143_, _26141_);
  nor (_26145_, _12237_, _06071_);
  or (_26147_, _26145_, _26144_);
  nand (_26148_, _26147_, _12588_);
  nor (_26149_, _12588_, _06075_);
  nor (_26150_, _26149_, _05976_);
  nand (_26151_, _26150_, _26148_);
  and (_26152_, _05976_, _06071_);
  nor (_26153_, _26152_, _06241_);
  and (_26154_, _26153_, _26151_);
  or (_26155_, _26154_, _26016_);
  nand (_26156_, _26155_, _08723_);
  and (_26158_, _06458_, _05970_);
  nor (_26159_, _26158_, _06369_);
  nand (_26160_, _26159_, _26156_);
  and (_26161_, _12303_, _06369_);
  nor (_26162_, _26161_, _12604_);
  nand (_26163_, _26162_, _26160_);
  nor (_26164_, _12603_, _06075_);
  nor (_26165_, _26164_, _05968_);
  nand (_26166_, _26165_, _26163_);
  and (_26167_, _12303_, _05968_);
  nor (_26169_, _26167_, _12615_);
  nand (_26170_, _26169_, _26166_);
  nor (_26171_, _12611_, _06071_);
  nor (_26172_, _26171_, _06332_);
  and (_26173_, _26172_, _26170_);
  and (_26174_, _06332_, _06075_);
  or (_26175_, _26174_, _05900_);
  or (_26176_, _26175_, _26173_);
  and (_26177_, _06458_, _05900_);
  nor (_26178_, _26177_, _12619_);
  nand (_26180_, _26178_, _26176_);
  and (_26181_, _26049_, _12619_);
  nor (_26182_, _26181_, _08973_);
  and (_26183_, _26182_, _26180_);
  or (_26184_, _26183_, _26015_);
  nand (_26185_, _26184_, _07198_);
  and (_26186_, _12304_, _06371_);
  nor (_26187_, _26186_, _10904_);
  nand (_26188_, _26187_, _26185_);
  and (_26189_, _10904_, _06075_);
  nor (_26191_, _26189_, _12634_);
  nand (_26192_, _26191_, _26188_);
  nor (_26193_, _12635_, _06086_);
  nor (_26194_, _26193_, _06331_);
  nand (_26195_, _26194_, _26192_);
  and (_26196_, _06331_, _06075_);
  nor (_26197_, _26196_, _05895_);
  nand (_26198_, _26197_, _26195_);
  and (_26199_, _06458_, _05895_);
  nor (_26200_, _26199_, _12677_);
  nand (_26202_, _26200_, _26198_);
  and (_26203_, _11291_, _06075_);
  and (_26204_, _26049_, _12684_);
  or (_26205_, _26204_, _26203_);
  and (_26206_, _26205_, _12677_);
  nor (_26207_, _26206_, _12682_);
  and (_26208_, _26207_, _26202_);
  or (_26209_, _26208_, _26013_);
  nand (_26210_, _26209_, _12228_);
  nor (_26211_, _12228_, _06075_);
  nor (_26213_, _26211_, _06367_);
  nand (_26214_, _26213_, _26210_);
  and (_26215_, _12303_, _06367_);
  nor (_26216_, _26215_, _06533_);
  and (_26217_, _26216_, _26214_);
  and (_26218_, _06533_, _06095_);
  or (_26219_, _26218_, _26217_);
  nand (_26220_, _26219_, _05890_);
  and (_26221_, _06458_, _05889_);
  nor (_26222_, _26221_, _12701_);
  nand (_26224_, _26222_, _26220_);
  nor (_26225_, _11291_, _06095_);
  and (_26226_, _26049_, _11291_);
  or (_26227_, _26226_, _26225_);
  and (_26228_, _26227_, _12701_);
  nor (_26229_, _26228_, _12710_);
  and (_26230_, _26229_, _26224_);
  or (_26231_, _26230_, _26012_);
  nand (_26232_, _26231_, _10967_);
  nor (_26233_, _10967_, _06075_);
  nor (_26235_, _26233_, _06366_);
  nand (_26236_, _26235_, _26232_);
  and (_26237_, _12303_, _06366_);
  nor (_26238_, _26237_, _06541_);
  and (_26239_, _26238_, _26236_);
  and (_26240_, _06541_, _06095_);
  or (_26241_, _26240_, _26239_);
  nand (_26242_, _26241_, _05919_);
  and (_26243_, _06458_, _07209_);
  nor (_26244_, _26243_, _12723_);
  nand (_26246_, _26244_, _26242_);
  nor (_26247_, _26049_, \oc8051_golden_model_1.PSW [7]);
  nor (_26248_, _06075_, _10854_);
  nor (_26249_, _26248_, _12724_);
  not (_26250_, _26249_);
  nor (_26251_, _26250_, _26247_);
  nor (_26252_, _26251_, _12738_);
  and (_26253_, _26252_, _26246_);
  or (_26254_, _26253_, _26011_);
  nand (_26255_, _26254_, _11005_);
  nor (_26257_, _11005_, _06075_);
  nor (_26258_, _26257_, _06383_);
  nand (_26259_, _26258_, _26255_);
  and (_26260_, _12303_, _06383_);
  nor (_26261_, _26260_, _06528_);
  and (_26262_, _26261_, _26259_);
  and (_26263_, _06528_, _06095_);
  or (_26264_, _26263_, _26262_);
  nand (_26265_, _26264_, _05922_);
  and (_26266_, _06458_, _12746_);
  nor (_26268_, _26266_, _12215_);
  nand (_26269_, _26268_, _26265_);
  and (_26270_, _06075_, _10854_);
  and (_26271_, _26049_, \oc8051_golden_model_1.PSW [7]);
  or (_26272_, _26271_, _26270_);
  and (_26273_, _26272_, _12215_);
  nor (_26274_, _26273_, _12758_);
  and (_26275_, _26274_, _26269_);
  or (_26276_, _26275_, _26010_);
  nand (_26277_, _26276_, _11051_);
  nor (_26279_, _11051_, _06075_);
  nor (_26280_, _26279_, _11080_);
  nand (_26281_, _26280_, _26277_);
  and (_26282_, _11080_, _06071_);
  nor (_26283_, _26282_, _06547_);
  and (_26284_, _26283_, _26281_);
  nor (_26285_, _09205_, _13873_);
  or (_26286_, _26285_, _26284_);
  nand (_26287_, _26286_, _05916_);
  and (_26288_, _06458_, _07228_);
  nor (_26290_, _26288_, _06381_);
  nand (_26291_, _26290_, _26287_);
  and (_26292_, _26022_, _12954_);
  nor (_26293_, _12303_, _12954_);
  or (_26294_, _26293_, _06946_);
  or (_26295_, _26294_, _26292_);
  and (_26296_, _26295_, _12105_);
  and (_26297_, _26296_, _26291_);
  or (_26298_, _26297_, _26009_);
  nand (_26299_, _26298_, _12963_);
  nor (_26301_, _12963_, _06075_);
  nor (_26302_, _26301_, _10448_);
  nand (_26303_, _26302_, _26299_);
  and (_26304_, _10448_, _06071_);
  nor (_26305_, _26304_, _06260_);
  and (_26306_, _26305_, _26303_);
  nor (_26307_, _09205_, _06261_);
  or (_26308_, _26307_, _26306_);
  nand (_26309_, _26308_, _05924_);
  and (_26310_, _06458_, _12089_);
  nor (_26312_, _26310_, _06377_);
  nand (_26313_, _26312_, _26309_);
  nor (_26314_, _26021_, _12954_);
  and (_26315_, _12304_, _12954_);
  nor (_26316_, _26315_, _26314_);
  and (_26317_, _26316_, _06377_);
  nor (_26318_, _26317_, _12985_);
  nand (_26319_, _26318_, _26313_);
  nor (_26320_, _12984_, _06071_);
  nor (_26321_, _26320_, _06563_);
  and (_26323_, _26321_, _26319_);
  or (_26324_, _26323_, _26008_);
  nand (_26325_, _26324_, _12991_);
  nor (_26326_, _12991_, _06062_);
  nor (_26327_, _26326_, _07812_);
  nand (_26328_, _26327_, _26325_);
  and (_26329_, _07812_, _06458_);
  nor (_26330_, _26329_, _06199_);
  nand (_26331_, _26330_, _26328_);
  and (_26332_, _26316_, _06199_);
  nor (_26334_, _26332_, _13007_);
  nand (_26335_, _26334_, _26331_);
  nor (_26336_, _13006_, _06071_);
  nor (_26337_, _26336_, _06188_);
  and (_26338_, _26337_, _26335_);
  or (_26339_, _26338_, _26007_);
  nand (_26340_, _26339_, _13013_);
  nor (_26341_, _13013_, _06062_);
  nor (_26342_, _26341_, _25220_);
  nand (_26343_, _26342_, _26340_);
  and (_26345_, _25220_, _06458_);
  nor (_26346_, _26345_, _13025_);
  and (_26347_, _26346_, _26343_);
  and (_26348_, _13025_, _06071_);
  or (_26349_, _26348_, _26347_);
  or (_26350_, _26349_, _01456_);
  or (_26351_, _01452_, \oc8051_golden_model_1.PC [3]);
  and (_26352_, _26351_, _43223_);
  and (_43858_, _26352_, _26350_);
  and (_26353_, _05571_, \oc8051_golden_model_1.PC [4]);
  nor (_26355_, _05571_, \oc8051_golden_model_1.PC [4]);
  nor (_26356_, _26355_, _26353_);
  and (_26357_, _26356_, _13025_);
  and (_26358_, _08834_, _07812_);
  and (_26359_, _12153_, _10854_);
  and (_26360_, _12174_, _12171_);
  nor (_26361_, _26360_, _12175_);
  and (_26362_, _26361_, \oc8051_golden_model_1.PSW [7]);
  or (_26363_, _26362_, _26359_);
  and (_26364_, _26363_, _12215_);
  nor (_26366_, _12153_, _08972_);
  and (_26367_, _12154_, _06241_);
  not (_26368_, _26356_);
  and (_26369_, _26368_, _12245_);
  and (_26370_, _12326_, _12323_);
  nor (_26371_, _26370_, _12327_);
  not (_26372_, _26371_);
  nor (_26373_, _26372_, _12533_);
  and (_26374_, _12533_, _12299_);
  nor (_26375_, _26374_, _26373_);
  nor (_26377_, _26375_, _12536_);
  and (_26378_, _12392_, _12300_);
  nor (_26379_, _26371_, _12392_);
  nor (_26380_, _26379_, _26378_);
  and (_26381_, _26380_, _06344_);
  and (_26382_, _12154_, _06483_);
  nand (_26383_, _12443_, _07338_);
  nand (_26384_, _26383_, _26368_);
  or (_26385_, _26371_, _12402_);
  or (_26386_, _12404_, _12299_);
  and (_26388_, _26386_, _26385_);
  or (_26389_, _26388_, _06252_);
  and (_26390_, _08834_, _06705_);
  and (_26391_, _12154_, _07123_);
  or (_26392_, _26391_, _06808_);
  nand (_26393_, _12419_, \oc8051_golden_model_1.PC [4]);
  and (_26394_, _26393_, _07124_);
  or (_26395_, _26394_, _26392_);
  or (_26396_, _26368_, _12420_);
  and (_26397_, _26396_, _07272_);
  and (_26399_, _26397_, _26395_);
  or (_26400_, _26399_, _12432_);
  or (_26401_, _26400_, _26390_);
  or (_26402_, _26368_, _12427_);
  and (_26403_, _26402_, _08573_);
  and (_26404_, _26403_, _26401_);
  nand (_26405_, _26361_, _12414_);
  and (_26406_, _26405_, _08572_);
  or (_26407_, _12414_, _12154_);
  and (_26408_, _26407_, _26406_);
  nor (_26410_, _26408_, _26404_);
  or (_26411_, _07134_, _06251_);
  or (_26412_, _26411_, _26410_);
  and (_26413_, _26412_, _26389_);
  or (_26414_, _26413_, _12444_);
  nand (_26415_, _26414_, _26384_);
  nand (_26416_, _26415_, _06476_);
  and (_26417_, _12154_, _06475_);
  nor (_26418_, _26417_, _07474_);
  and (_26419_, _26418_, _26416_);
  nor (_26420_, _08834_, _05950_);
  or (_26421_, _26420_, _06468_);
  nor (_26422_, _26421_, _26419_);
  and (_26423_, _12154_, _06468_);
  or (_26424_, _26423_, _26422_);
  and (_26425_, _26424_, _12451_);
  nor (_26426_, _26356_, _12451_);
  or (_26427_, _26426_, _26425_);
  nand (_26428_, _26427_, _06801_);
  and (_26429_, _12154_, _06466_);
  nor (_26432_, _26429_, _12464_);
  nand (_26433_, _26432_, _26428_);
  nor (_26434_, _26368_, _12462_);
  nor (_26435_, _26434_, _06483_);
  and (_26436_, _26435_, _26433_);
  or (_26437_, _26436_, _26382_);
  nand (_26438_, _26437_, _05953_);
  and (_26439_, _08834_, _12466_);
  nor (_26440_, _26439_, _06247_);
  nand (_26441_, _26440_, _26438_);
  and (_26443_, _12153_, _06247_);
  nor (_26444_, _26443_, _12479_);
  nand (_26445_, _26444_, _26441_);
  and (_26446_, _12513_, _12299_);
  nor (_26447_, _26372_, _12513_);
  or (_26448_, _26447_, _12478_);
  nor (_26449_, _26448_, _26446_);
  nor (_26450_, _26449_, _06344_);
  and (_26451_, _26450_, _26445_);
  or (_26452_, _26451_, _26381_);
  and (_26454_, _26452_, _12536_);
  or (_26455_, _26454_, _26377_);
  nand (_26456_, _26455_, _12522_);
  nor (_26457_, _26371_, _12555_);
  and (_26458_, _12555_, _12300_);
  or (_26459_, _26458_, _12522_);
  nor (_26460_, _26459_, _26457_);
  nor (_26461_, _26460_, _12245_);
  and (_26462_, _26461_, _26456_);
  or (_26463_, _26462_, _26369_);
  nand (_26465_, _26463_, _07164_);
  and (_26466_, _12154_, _06461_);
  nor (_26467_, _26466_, _07471_);
  nand (_26468_, _26467_, _26465_);
  nor (_26469_, _08834_, _05947_);
  nor (_26470_, _26469_, _25366_);
  nand (_26471_, _26470_, _26468_);
  nor (_26472_, _25365_, _12153_);
  nor (_26473_, _26472_, _12243_);
  and (_26474_, _26473_, _26471_);
  nor (_26476_, _26368_, _12242_);
  or (_26477_, _26476_, _06505_);
  nor (_26478_, _26477_, _26474_);
  and (_26479_, _12154_, _06505_);
  or (_26480_, _26479_, _26478_);
  nand (_26481_, _26480_, _05958_);
  and (_26482_, _08834_, _25090_);
  nor (_26483_, _26482_, _06504_);
  and (_26484_, _26483_, _26481_);
  and (_26485_, _12153_, _06504_);
  or (_26486_, _26485_, _26484_);
  nand (_26487_, _26486_, _12237_);
  nor (_26488_, _26368_, _12237_);
  nor (_26489_, _26488_, _12589_);
  nand (_26490_, _26489_, _26487_);
  nor (_26491_, _12588_, _12153_);
  nor (_26492_, _26491_, _05976_);
  nand (_26493_, _26492_, _26490_);
  and (_26494_, _26356_, _05976_);
  nor (_26495_, _26494_, _06241_);
  and (_26497_, _26495_, _26493_);
  or (_26498_, _26497_, _26367_);
  nand (_26499_, _26498_, _08723_);
  and (_26500_, _08834_, _05970_);
  nor (_26501_, _26500_, _06369_);
  nand (_26502_, _26501_, _26499_);
  and (_26503_, _12299_, _06369_);
  nor (_26504_, _26503_, _12604_);
  nand (_26505_, _26504_, _26502_);
  nor (_26506_, _12603_, _12153_);
  nor (_26508_, _26506_, _05968_);
  nand (_26509_, _26508_, _26505_);
  and (_26510_, _12299_, _05968_);
  nor (_26511_, _26510_, _12615_);
  nand (_26512_, _26511_, _26509_);
  nor (_26513_, _26356_, _12611_);
  nor (_26514_, _26513_, _06332_);
  and (_26515_, _26514_, _26512_);
  nor (_26516_, _12153_, _05900_);
  nor (_26517_, _26516_, _12613_);
  or (_26518_, _26517_, _26515_);
  and (_26519_, _08834_, _05900_);
  nor (_26520_, _26519_, _12619_);
  nand (_26521_, _26520_, _26518_);
  and (_26522_, _26361_, _12619_);
  nor (_26523_, _26522_, _08973_);
  and (_26524_, _26523_, _26521_);
  or (_26525_, _26524_, _26366_);
  nand (_26526_, _26525_, _07198_);
  and (_26527_, _12300_, _06371_);
  nor (_26528_, _26527_, _10904_);
  and (_26529_, _26528_, _26526_);
  and (_26530_, _12153_, _10904_);
  or (_26531_, _26530_, _26529_);
  nand (_26532_, _26531_, _12635_);
  and (_26533_, _12651_, _12648_);
  nor (_26534_, _26533_, _12652_);
  and (_26535_, _26534_, _12634_);
  nor (_26536_, _26535_, _06331_);
  and (_26537_, _26536_, _26532_);
  and (_26538_, _12154_, _06331_);
  or (_26539_, _26538_, _26537_);
  nand (_26540_, _26539_, _13846_);
  and (_26541_, _08834_, _05895_);
  nor (_26542_, _26541_, _12677_);
  and (_26543_, _26542_, _26540_);
  and (_26544_, _12153_, _11291_);
  and (_26545_, _26361_, _12684_);
  or (_26546_, _26545_, _26544_);
  and (_26547_, _26546_, _12677_);
  or (_26548_, _26547_, _26543_);
  nand (_26549_, _26548_, _12232_);
  nor (_26550_, _26368_, _12232_);
  nor (_26551_, _26550_, _12229_);
  nand (_26552_, _26551_, _26549_);
  nor (_26553_, _12153_, _12228_);
  nor (_26554_, _26553_, _06367_);
  nand (_26555_, _26554_, _26552_);
  and (_26556_, _12299_, _06367_);
  nor (_26557_, _26556_, _06533_);
  and (_26558_, _26557_, _26555_);
  and (_26559_, _12154_, _06533_);
  or (_26560_, _26559_, _26558_);
  nand (_26561_, _26560_, _05890_);
  and (_26562_, _08834_, _05889_);
  nor (_26563_, _26562_, _12701_);
  and (_26564_, _26563_, _26561_);
  nor (_26565_, _12154_, _11291_);
  and (_26566_, _26361_, _11291_);
  or (_26567_, _26566_, _26565_);
  and (_26569_, _26567_, _12701_);
  or (_26570_, _26569_, _26564_);
  nand (_26571_, _26570_, _12226_);
  nor (_26572_, _26368_, _12226_);
  nor (_26573_, _26572_, _10968_);
  nand (_26574_, _26573_, _26571_);
  nor (_26575_, _12153_, _10967_);
  nor (_26576_, _26575_, _06366_);
  nand (_26577_, _26576_, _26574_);
  and (_26578_, _12299_, _06366_);
  nor (_26580_, _26578_, _06541_);
  and (_26581_, _26580_, _26577_);
  and (_26582_, _12154_, _06541_);
  or (_26583_, _26582_, _26581_);
  nand (_26584_, _26583_, _05919_);
  and (_26585_, _08834_, _07209_);
  nor (_26586_, _26585_, _12723_);
  and (_26587_, _26586_, _26584_);
  and (_26588_, _12153_, \oc8051_golden_model_1.PSW [7]);
  and (_26589_, _26361_, _10854_);
  or (_26590_, _26589_, _26588_);
  and (_26591_, _26590_, _12723_);
  or (_26592_, _26591_, _26587_);
  nand (_26593_, _26592_, _12736_);
  nor (_26594_, _26368_, _12736_);
  nor (_26595_, _26594_, _11006_);
  nand (_26596_, _26595_, _26593_);
  nor (_26597_, _12153_, _11005_);
  nor (_26598_, _26597_, _06383_);
  nand (_26599_, _26598_, _26596_);
  and (_26601_, _12299_, _06383_);
  nor (_26602_, _26601_, _06528_);
  and (_26603_, _26602_, _26599_);
  and (_26604_, _12154_, _06528_);
  or (_26605_, _26604_, _26603_);
  nand (_26606_, _26605_, _05922_);
  and (_26607_, _08834_, _12746_);
  nor (_26608_, _26607_, _12215_);
  and (_26609_, _26608_, _26606_);
  or (_26610_, _26609_, _26364_);
  nand (_26612_, _26610_, _12756_);
  nor (_26613_, _26368_, _12756_);
  nor (_26614_, _26613_, _11052_);
  nand (_26615_, _26614_, _26612_);
  nor (_26616_, _12153_, _11051_);
  nor (_26617_, _26616_, _11080_);
  nand (_26618_, _26617_, _26615_);
  and (_26619_, _26356_, _11080_);
  nor (_26620_, _26619_, _06547_);
  and (_26621_, _26620_, _26618_);
  nor (_26623_, _09159_, _13873_);
  or (_26624_, _26623_, _26621_);
  nand (_26625_, _26624_, _05916_);
  and (_26626_, _08834_, _07228_);
  nor (_26627_, _26626_, _06381_);
  and (_26628_, _26627_, _26625_);
  nor (_26629_, _12300_, _12954_);
  and (_26630_, _26371_, _12954_);
  nor (_26631_, _26630_, _26629_);
  nor (_26632_, _26631_, _06946_);
  or (_26634_, _26632_, _26628_);
  nand (_26635_, _26634_, _12105_);
  nor (_26636_, _26368_, _12105_);
  nor (_26637_, _26636_, _12964_);
  nand (_26638_, _26637_, _26635_);
  nor (_26639_, _12963_, _12153_);
  nor (_26640_, _26639_, _10448_);
  nand (_26641_, _26640_, _26638_);
  and (_26642_, _26356_, _10448_);
  nor (_26643_, _26642_, _06260_);
  nand (_26644_, _26643_, _26641_);
  nor (_26645_, _09159_, _06261_);
  nor (_26646_, _26645_, _12089_);
  nand (_26647_, _26646_, _26644_);
  nor (_26648_, _08834_, _05924_);
  nor (_26649_, _26648_, _06377_);
  nand (_26650_, _26649_, _26647_);
  and (_26651_, _12300_, _12954_);
  nor (_26652_, _26371_, _12954_);
  nor (_26653_, _26652_, _26651_);
  nor (_26655_, _26653_, _06564_);
  nor (_26656_, _26655_, _12985_);
  nand (_26657_, _26656_, _26650_);
  nor (_26658_, _26368_, _12984_);
  nor (_26659_, _26658_, _06563_);
  nand (_26660_, _26659_, _26657_);
  and (_26661_, _12154_, _06563_);
  nor (_26662_, _26661_, _12992_);
  nand (_26663_, _26662_, _26660_);
  nor (_26664_, _26368_, _12991_);
  nor (_26666_, _26664_, _07812_);
  and (_26667_, _26666_, _26663_);
  or (_26668_, _26667_, _26358_);
  nand (_26669_, _26668_, _06571_);
  nor (_26670_, _26653_, _06571_);
  nor (_26671_, _26670_, _13007_);
  nand (_26672_, _26671_, _26669_);
  nor (_26673_, _26368_, _13006_);
  nor (_26674_, _26673_, _06188_);
  nand (_26675_, _26674_, _26672_);
  and (_26677_, _12154_, _06188_);
  nor (_26678_, _26677_, _13014_);
  nand (_26679_, _26678_, _26675_);
  nor (_26680_, _26368_, _13013_);
  nor (_26681_, _26680_, _25220_);
  nand (_26682_, _26681_, _26679_);
  and (_26683_, _25220_, _08834_);
  nor (_26684_, _26683_, _13025_);
  and (_26685_, _26684_, _26682_);
  or (_26686_, _26685_, _26357_);
  or (_26688_, _26686_, _01456_);
  or (_26689_, _01452_, \oc8051_golden_model_1.PC [4]);
  and (_26690_, _26689_, _43223_);
  and (_43859_, _26690_, _26688_);
  nor (_26691_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_26692_, _12148_, _05557_);
  nor (_26693_, _26692_, _26691_);
  and (_26694_, _26693_, _13025_);
  and (_26695_, _12148_, _06188_);
  and (_26696_, _12148_, _06563_);
  nor (_26698_, _26693_, _12105_);
  nor (_26699_, _26693_, _12756_);
  nor (_26700_, _26693_, _12736_);
  nor (_26701_, _26693_, _12226_);
  nor (_26702_, _26693_, _12232_);
  nor (_26703_, _12148_, _08972_);
  and (_26704_, _12149_, _06241_);
  nor (_26705_, _26693_, _12237_);
  not (_26706_, _26693_);
  and (_26707_, _26706_, _12245_);
  or (_26708_, _12297_, _12296_);
  not (_26709_, _26708_);
  nor (_26710_, _26709_, _12328_);
  and (_26711_, _26709_, _12328_);
  nor (_26712_, _26711_, _26710_);
  nor (_26713_, _26712_, _12533_);
  and (_26714_, _12533_, _12294_);
  nor (_26715_, _26714_, _26713_);
  or (_26716_, _26715_, _12536_);
  nor (_26717_, _08867_, _07272_);
  and (_26719_, _12149_, _07123_);
  nor (_26720_, _26719_, _06808_);
  and (_26721_, _12419_, \oc8051_golden_model_1.PC [5]);
  or (_26722_, _26721_, _07123_);
  and (_26723_, _26722_, _26720_);
  or (_26724_, _26706_, _12420_);
  nand (_26725_, _26724_, _12427_);
  or (_26726_, _26725_, _26723_);
  and (_26727_, _26726_, _07272_);
  nor (_26728_, _26727_, _26717_);
  nor (_26730_, _26693_, _12427_);
  nor (_26731_, _26730_, _26728_);
  nor (_26732_, _26731_, _08572_);
  or (_26733_, _12414_, _12149_);
  or (_26734_, _12151_, _12150_);
  and (_26735_, _26734_, _12176_);
  nor (_26736_, _26734_, _12176_);
  or (_26737_, _26736_, _26735_);
  or (_26738_, _26737_, _12412_);
  and (_26739_, _26738_, _08572_);
  and (_26741_, _26739_, _26733_);
  or (_26742_, _26741_, _26732_);
  nand (_26743_, _26742_, _07338_);
  and (_26744_, _26706_, _07134_);
  nor (_26745_, _26744_, _06251_);
  nand (_26746_, _26745_, _26743_);
  not (_26747_, _26712_);
  or (_26748_, _26747_, _12402_);
  and (_26749_, _26748_, _06251_);
  or (_26750_, _12404_, _12294_);
  nand (_26752_, _26750_, _26749_);
  and (_26753_, _26752_, _12443_);
  nand (_26754_, _26753_, _26746_);
  nor (_26755_, _26693_, _12443_);
  nor (_26756_, _26755_, _06475_);
  nand (_26757_, _26756_, _26754_);
  and (_26758_, _12148_, _06475_);
  nor (_26759_, _26758_, _07474_);
  nand (_26760_, _26759_, _26757_);
  and (_26761_, _08867_, _07474_);
  nor (_26763_, _26761_, _06468_);
  nand (_26764_, _26763_, _26760_);
  and (_26765_, _12148_, _06468_);
  nor (_26766_, _26765_, _12452_);
  nand (_26767_, _26766_, _26764_);
  nor (_26768_, _26693_, _12451_);
  nor (_26769_, _26768_, _06466_);
  nand (_26770_, _26769_, _26767_);
  and (_26771_, _12148_, _06466_);
  nor (_26772_, _26771_, _12464_);
  nand (_26773_, _26772_, _26770_);
  nor (_26774_, _26693_, _12462_);
  nor (_26775_, _26774_, _06483_);
  nand (_26776_, _26775_, _26773_);
  and (_26777_, _12148_, _06483_);
  nor (_26778_, _26777_, _12466_);
  nand (_26779_, _26778_, _26776_);
  and (_26780_, _08867_, _12466_);
  nor (_26781_, _26780_, _06247_);
  nand (_26782_, _26781_, _26779_);
  and (_26784_, _12148_, _06247_);
  nor (_26785_, _26784_, _12479_);
  and (_26786_, _26785_, _26782_);
  and (_26787_, _12513_, _12294_);
  nor (_26788_, _26712_, _12513_);
  or (_26789_, _26788_, _26787_);
  nor (_26790_, _26789_, _12478_);
  or (_26791_, _26790_, _26786_);
  nand (_26792_, _26791_, _06345_);
  or (_26793_, _26712_, _12392_);
  nand (_26795_, _12392_, _12294_);
  and (_26796_, _26795_, _06344_);
  nand (_26797_, _26796_, _26793_);
  nand (_26798_, _26797_, _26792_);
  or (_26799_, _26798_, _06338_);
  and (_26800_, _26799_, _26716_);
  or (_26801_, _26800_, _06373_);
  and (_26802_, _12555_, _12294_);
  nor (_26803_, _26712_, _12555_);
  or (_26804_, _26803_, _26802_);
  and (_26806_, _26804_, _06373_);
  nor (_26807_, _26806_, _12245_);
  and (_26808_, _26807_, _26801_);
  or (_26809_, _26808_, _26707_);
  nand (_26810_, _26809_, _07164_);
  and (_26811_, _12149_, _06461_);
  nor (_26812_, _26811_, _07471_);
  nand (_26813_, _26812_, _26810_);
  nor (_26814_, _08867_, _05947_);
  nor (_26815_, _26814_, _25366_);
  and (_26817_, _26815_, _26813_);
  nor (_26818_, _25365_, _12148_);
  or (_26819_, _26818_, _26817_);
  nand (_26820_, _26819_, _12242_);
  nor (_26821_, _26693_, _12242_);
  nor (_26822_, _26821_, _06505_);
  nand (_26823_, _26822_, _26820_);
  and (_26824_, _12148_, _06505_);
  nor (_26825_, _26824_, _25090_);
  nand (_26826_, _26825_, _26823_);
  and (_26828_, _08867_, _25090_);
  nor (_26829_, _26828_, _06504_);
  nand (_26830_, _26829_, _26826_);
  and (_26831_, _12148_, _06504_);
  nor (_26832_, _26831_, _12582_);
  and (_26833_, _26832_, _26830_);
  or (_26834_, _26833_, _26705_);
  nand (_26835_, _26834_, _12588_);
  nor (_26836_, _12588_, _12148_);
  nor (_26837_, _26836_, _05976_);
  nand (_26838_, _26837_, _26835_);
  and (_26839_, _26693_, _05976_);
  nor (_26840_, _26839_, _06241_);
  and (_26841_, _26840_, _26838_);
  or (_26842_, _26841_, _26704_);
  nand (_26843_, _26842_, _08723_);
  and (_26844_, _08867_, _05970_);
  nor (_26845_, _26844_, _06369_);
  nand (_26846_, _26845_, _26843_);
  and (_26847_, _12294_, _06369_);
  nor (_26849_, _26847_, _12604_);
  nand (_26850_, _26849_, _26846_);
  nor (_26851_, _12603_, _12148_);
  nor (_26852_, _26851_, _05968_);
  nand (_26853_, _26852_, _26850_);
  and (_26854_, _12294_, _05968_);
  nor (_26855_, _26854_, _12615_);
  nand (_26856_, _26855_, _26853_);
  nor (_26857_, _26693_, _12611_);
  nor (_26858_, _26857_, _06332_);
  and (_26860_, _26858_, _26856_);
  and (_26861_, _12148_, _06332_);
  or (_26862_, _26861_, _05900_);
  or (_26863_, _26862_, _26860_);
  and (_26864_, _08867_, _05900_);
  nor (_26865_, _26864_, _12619_);
  nand (_26866_, _26865_, _26863_);
  nor (_26867_, _26737_, _12620_);
  nor (_26868_, _26867_, _08973_);
  and (_26869_, _26868_, _26866_);
  or (_26871_, _26869_, _26703_);
  nand (_26872_, _26871_, _07198_);
  and (_26873_, _12295_, _06371_);
  nor (_26874_, _26873_, _10904_);
  nand (_26875_, _26874_, _26872_);
  and (_26876_, _12148_, _10904_);
  nor (_26877_, _26876_, _12634_);
  nand (_26878_, _26877_, _26875_);
  and (_26879_, _12653_, _12646_);
  nor (_26880_, _26879_, _12654_);
  nor (_26882_, _26880_, _12635_);
  nor (_26883_, _26882_, _06331_);
  nand (_26884_, _26883_, _26878_);
  and (_26885_, _12148_, _06331_);
  nor (_26886_, _26885_, _05895_);
  nand (_26887_, _26886_, _26884_);
  and (_26888_, _08867_, _05895_);
  nor (_26889_, _26888_, _12677_);
  nand (_26890_, _26889_, _26887_);
  and (_26891_, _12148_, _11291_);
  nor (_26893_, _26737_, _11291_);
  or (_26894_, _26893_, _26891_);
  and (_26895_, _26894_, _12677_);
  nor (_26896_, _26895_, _12682_);
  and (_26897_, _26896_, _26890_);
  or (_26898_, _26897_, _26702_);
  nand (_26899_, _26898_, _12228_);
  nor (_26900_, _12148_, _12228_);
  nor (_26901_, _26900_, _06367_);
  nand (_26902_, _26901_, _26899_);
  and (_26903_, _12294_, _06367_);
  nor (_26904_, _26903_, _06533_);
  and (_26905_, _26904_, _26902_);
  and (_26906_, _12149_, _06533_);
  or (_26907_, _26906_, _26905_);
  nand (_26908_, _26907_, _05890_);
  and (_26909_, _08867_, _05889_);
  nor (_26910_, _26909_, _12701_);
  nand (_26911_, _26910_, _26908_);
  nor (_26912_, _12149_, _11291_);
  nor (_26914_, _26737_, _12684_);
  or (_26915_, _26914_, _26912_);
  and (_26916_, _26915_, _12701_);
  nor (_26917_, _26916_, _12710_);
  and (_26918_, _26917_, _26911_);
  or (_26919_, _26918_, _26701_);
  nand (_26920_, _26919_, _10967_);
  nor (_26921_, _12148_, _10967_);
  nor (_26922_, _26921_, _06366_);
  nand (_26923_, _26922_, _26920_);
  and (_26925_, _12294_, _06366_);
  nor (_26926_, _26925_, _06541_);
  and (_26927_, _26926_, _26923_);
  and (_26928_, _12149_, _06541_);
  or (_26929_, _26928_, _26927_);
  nand (_26930_, _26929_, _05919_);
  and (_26931_, _08867_, _07209_);
  nor (_26932_, _26931_, _12723_);
  nand (_26933_, _26932_, _26930_);
  and (_26934_, _26737_, _10854_);
  nor (_26936_, _12148_, _10854_);
  nor (_26937_, _26936_, _12724_);
  not (_26938_, _26937_);
  nor (_26939_, _26938_, _26934_);
  nor (_26940_, _26939_, _12738_);
  and (_26941_, _26940_, _26933_);
  or (_26942_, _26941_, _26700_);
  nand (_26943_, _26942_, _11005_);
  nor (_26944_, _12148_, _11005_);
  nor (_26945_, _26944_, _06383_);
  nand (_26947_, _26945_, _26943_);
  and (_26948_, _12294_, _06383_);
  nor (_26949_, _26948_, _06528_);
  and (_26950_, _26949_, _26947_);
  and (_26951_, _12149_, _06528_);
  or (_26952_, _26951_, _26950_);
  nand (_26953_, _26952_, _05922_);
  and (_26954_, _08867_, _12746_);
  nor (_26955_, _26954_, _12215_);
  nand (_26956_, _26955_, _26953_);
  and (_26958_, _12148_, _10854_);
  nor (_26959_, _26737_, _10854_);
  or (_26960_, _26959_, _26958_);
  and (_26961_, _26960_, _12215_);
  nor (_26962_, _26961_, _12758_);
  and (_26963_, _26962_, _26956_);
  or (_26964_, _26963_, _26699_);
  nand (_26965_, _26964_, _11051_);
  nor (_26966_, _12148_, _11051_);
  nor (_26967_, _26966_, _11080_);
  nand (_26969_, _26967_, _26965_);
  and (_26970_, _26693_, _11080_);
  nor (_26971_, _26970_, _06547_);
  and (_26972_, _26971_, _26969_);
  nor (_26973_, _09113_, _13873_);
  or (_26974_, _26973_, _26972_);
  nand (_26975_, _26974_, _05916_);
  and (_26976_, _08867_, _07228_);
  nor (_26977_, _26976_, _06381_);
  nand (_26978_, _26977_, _26975_);
  and (_26980_, _26712_, _12954_);
  nor (_26981_, _12294_, _12954_);
  or (_26982_, _26981_, _06946_);
  or (_26983_, _26982_, _26980_);
  and (_26984_, _26983_, _12105_);
  and (_26985_, _26984_, _26978_);
  or (_26986_, _26985_, _26698_);
  nand (_26987_, _26986_, _12963_);
  nor (_26988_, _12963_, _12148_);
  nor (_26989_, _26988_, _10448_);
  nand (_26990_, _26989_, _26987_);
  and (_26991_, _26693_, _10448_);
  nor (_26992_, _26991_, _06260_);
  and (_26993_, _26992_, _26990_);
  nor (_26994_, _09113_, _06261_);
  or (_26995_, _26994_, _26993_);
  nand (_26996_, _26995_, _05924_);
  and (_26997_, _08867_, _12089_);
  nor (_26998_, _26997_, _06377_);
  nand (_26999_, _26998_, _26996_);
  and (_27001_, _12295_, _12954_);
  nor (_27002_, _26747_, _12954_);
  nor (_27003_, _27002_, _27001_);
  and (_27004_, _27003_, _06377_);
  nor (_27005_, _27004_, _12985_);
  nand (_27006_, _27005_, _26999_);
  nor (_27007_, _26693_, _12984_);
  nor (_27008_, _27007_, _06563_);
  and (_27009_, _27008_, _27006_);
  or (_27010_, _27009_, _26696_);
  nand (_27012_, _27010_, _12991_);
  nor (_27013_, _26706_, _12991_);
  nor (_27014_, _27013_, _07812_);
  nand (_27015_, _27014_, _27012_);
  and (_27016_, _08867_, _07812_);
  nor (_27017_, _27016_, _06199_);
  nand (_27018_, _27017_, _27015_);
  and (_27019_, _27003_, _06199_);
  nor (_27020_, _27019_, _13007_);
  nand (_27021_, _27020_, _27018_);
  nor (_27023_, _26693_, _13006_);
  nor (_27024_, _27023_, _06188_);
  and (_27025_, _27024_, _27021_);
  or (_27026_, _27025_, _26695_);
  nand (_27027_, _27026_, _13013_);
  nor (_27028_, _26706_, _13013_);
  nor (_27029_, _27028_, _25220_);
  nand (_27030_, _27029_, _27027_);
  and (_27031_, _25220_, _08867_);
  nor (_27032_, _27031_, _13025_);
  and (_27034_, _27032_, _27030_);
  or (_27035_, _27034_, _26694_);
  or (_27036_, _27035_, _01456_);
  or (_27037_, _01452_, \oc8051_golden_model_1.PC [5]);
  and (_27038_, _27037_, _43223_);
  and (_43860_, _27038_, _27036_);
  and (_27039_, _25220_, _08802_);
  and (_27040_, _08513_, _05571_);
  nor (_27041_, _27040_, \oc8051_golden_model_1.PC [6]);
  nor (_27042_, _27041_, _12091_);
  not (_27044_, _27042_);
  nor (_27045_, _27044_, _13013_);
  nand (_27046_, _08802_, _07812_);
  nand (_27047_, _27044_, _10448_);
  nand (_27048_, _27044_, _12245_);
  nand (_27049_, _12142_, _06483_);
  or (_27050_, _27042_, _12451_);
  nor (_27051_, _12331_, _12291_);
  nor (_27052_, _27051_, _12332_);
  or (_27053_, _27052_, _12402_);
  or (_27054_, _12404_, _12287_);
  and (_27055_, _27054_, _06251_);
  and (_27056_, _27055_, _27053_);
  and (_27057_, _12412_, _12141_);
  nor (_27058_, _12179_, _12145_);
  nor (_27059_, _27058_, _12180_);
  and (_27060_, _27059_, _12414_);
  or (_27061_, _27060_, _27057_);
  or (_27062_, _27061_, _08573_);
  and (_27063_, _08802_, _06705_);
  and (_27065_, _12142_, _07123_);
  or (_27066_, _27065_, _06808_);
  nand (_27067_, _12419_, \oc8051_golden_model_1.PC [6]);
  and (_27068_, _27067_, _07124_);
  or (_27069_, _27068_, _27066_);
  or (_27070_, _27044_, _12420_);
  and (_27071_, _27070_, _07272_);
  and (_27072_, _27071_, _27069_);
  or (_27073_, _27072_, _12432_);
  or (_27074_, _27073_, _27063_);
  or (_27076_, _27044_, _12427_);
  and (_27077_, _27076_, _08573_);
  and (_27078_, _27077_, _27074_);
  nor (_27079_, _27078_, _26411_);
  and (_27080_, _27079_, _27062_);
  or (_27081_, _27080_, _27056_);
  and (_27082_, _27081_, _12443_);
  and (_27083_, _27042_, _26383_);
  or (_27084_, _27083_, _06475_);
  or (_27085_, _27084_, _27082_);
  nand (_27087_, _12142_, _06475_);
  and (_27088_, _27087_, _05950_);
  and (_27089_, _27088_, _27085_);
  nor (_27090_, _08802_, _05950_);
  or (_27091_, _27090_, _06468_);
  or (_27092_, _27091_, _27089_);
  nand (_27093_, _12142_, _06468_);
  and (_27094_, _27093_, _27092_);
  or (_27095_, _27094_, _12452_);
  and (_27096_, _27095_, _27050_);
  or (_27098_, _27096_, _06466_);
  nand (_27099_, _12142_, _06466_);
  and (_27100_, _27099_, _12462_);
  and (_27101_, _27100_, _27098_);
  nor (_27102_, _27044_, _12462_);
  or (_27103_, _27102_, _06483_);
  or (_27104_, _27103_, _27101_);
  and (_27105_, _27104_, _27049_);
  or (_27106_, _27105_, _12466_);
  nand (_27107_, _08802_, _12466_);
  and (_27109_, _27107_, _07523_);
  and (_27110_, _27109_, _27106_);
  nand (_27111_, _12141_, _06247_);
  nand (_27112_, _27111_, _12478_);
  or (_27113_, _27112_, _27110_);
  or (_27114_, _27052_, _12513_);
  nand (_27115_, _12513_, _12288_);
  and (_27116_, _27115_, _27114_);
  or (_27117_, _27116_, _12478_);
  and (_27118_, _27117_, _27113_);
  or (_27120_, _27118_, _06344_);
  and (_27121_, _12392_, _12287_);
  not (_27122_, _12392_);
  and (_27123_, _27052_, _27122_);
  or (_27124_, _27123_, _06345_);
  or (_27125_, _27124_, _27121_);
  and (_27126_, _27125_, _12536_);
  and (_27127_, _27126_, _27120_);
  and (_27128_, _27052_, _12534_);
  and (_27129_, _12533_, _12287_);
  or (_27131_, _27129_, _27128_);
  and (_27132_, _27131_, _06338_);
  or (_27133_, _27132_, _27127_);
  and (_27134_, _27133_, _12522_);
  or (_27135_, _27052_, _12555_);
  nand (_27136_, _12555_, _12288_);
  and (_27137_, _27136_, _06373_);
  and (_27138_, _27137_, _27135_);
  or (_27139_, _27138_, _12245_);
  or (_27140_, _27139_, _27134_);
  and (_27142_, _27140_, _27048_);
  or (_27143_, _27142_, _06461_);
  nand (_27144_, _12142_, _06461_);
  and (_27145_, _27144_, _05947_);
  and (_27146_, _27145_, _27143_);
  nor (_27147_, _08802_, _05947_);
  or (_27148_, _27147_, _25366_);
  or (_27149_, _27148_, _27146_);
  or (_27150_, _25365_, _12141_);
  and (_27151_, _27150_, _27149_);
  or (_27153_, _27151_, _12243_);
  or (_27154_, _27042_, _12242_);
  and (_27155_, _27154_, _14007_);
  and (_27156_, _27155_, _27153_);
  and (_27157_, _12141_, _06505_);
  or (_27158_, _27157_, _25090_);
  or (_27159_, _27158_, _27156_);
  nand (_27160_, _08802_, _25090_);
  and (_27161_, _27160_, _14006_);
  and (_27162_, _27161_, _27159_);
  nand (_27164_, _12141_, _06504_);
  nand (_27165_, _27164_, _12237_);
  or (_27166_, _27165_, _27162_);
  or (_27167_, _27042_, _12237_);
  and (_27168_, _27167_, _12588_);
  and (_27169_, _27168_, _27166_);
  nor (_27170_, _12588_, _12142_);
  or (_27171_, _27170_, _05976_);
  or (_27172_, _27171_, _27169_);
  nand (_27173_, _27044_, _05976_);
  and (_27175_, _27173_, _27172_);
  or (_27176_, _27175_, _06241_);
  nand (_27177_, _12142_, _06241_);
  and (_27178_, _27177_, _08723_);
  and (_27179_, _27178_, _27176_);
  nor (_27180_, _08802_, _08723_);
  or (_27181_, _27180_, _06369_);
  or (_27182_, _27181_, _27179_);
  nand (_27183_, _12288_, _06369_);
  and (_27184_, _27183_, _12603_);
  and (_27186_, _27184_, _27182_);
  nor (_27187_, _12603_, _12142_);
  or (_27188_, _27187_, _05968_);
  or (_27189_, _27188_, _27186_);
  nand (_27190_, _12288_, _05968_);
  and (_27191_, _27190_, _12611_);
  and (_27192_, _27191_, _27189_);
  nor (_27193_, _27044_, _12611_);
  or (_27194_, _27193_, _06332_);
  or (_27195_, _27194_, _27192_);
  nand (_27197_, _12142_, _06332_);
  and (_27198_, _27197_, _25117_);
  and (_27199_, _27198_, _27195_);
  nor (_27200_, _08802_, _25117_);
  or (_27201_, _27200_, _12619_);
  or (_27202_, _27201_, _27199_);
  or (_27203_, _27059_, _12620_);
  and (_27204_, _27203_, _27202_);
  and (_27205_, _27204_, _08972_);
  nor (_27206_, _12142_, _08972_);
  or (_27208_, _27206_, _06371_);
  or (_27209_, _27208_, _27205_);
  nand (_27210_, _12288_, _06371_);
  and (_27211_, _27210_, _10905_);
  and (_27212_, _27211_, _27209_);
  and (_27213_, _12141_, _10904_);
  or (_27214_, _27213_, _12634_);
  or (_27215_, _27214_, _27212_);
  nor (_27216_, _12656_, _12642_);
  nor (_27217_, _27216_, _12657_);
  or (_27218_, _27217_, _12635_);
  and (_27219_, _27218_, _06921_);
  and (_27220_, _27219_, _27215_);
  and (_27221_, _12141_, _06331_);
  or (_27222_, _27221_, _05895_);
  or (_27223_, _27222_, _27220_);
  nand (_27224_, _08802_, _05895_);
  and (_27225_, _27224_, _12678_);
  and (_27226_, _27225_, _27223_);
  or (_27227_, _27059_, _11291_);
  nand (_27230_, _12142_, _11291_);
  and (_27231_, _27230_, _12677_);
  and (_27232_, _27231_, _27227_);
  or (_27233_, _27232_, _12682_);
  or (_27234_, _27233_, _27226_);
  or (_27235_, _27042_, _12232_);
  and (_27236_, _27235_, _12228_);
  and (_27237_, _27236_, _27234_);
  nor (_27238_, _12142_, _12228_);
  or (_27239_, _27238_, _06367_);
  or (_27241_, _27239_, _27237_);
  nand (_27242_, _12288_, _06367_);
  and (_27243_, _27242_, _27241_);
  or (_27244_, _27243_, _06533_);
  nand (_27245_, _12142_, _06533_);
  and (_27246_, _27245_, _05890_);
  and (_27247_, _27246_, _27244_);
  nor (_27248_, _08802_, _05890_);
  or (_27249_, _27248_, _27247_);
  and (_27250_, _27249_, _12702_);
  or (_27252_, _27059_, _12684_);
  or (_27253_, _12141_, _11291_);
  and (_27254_, _27253_, _12701_);
  and (_27255_, _27254_, _27252_);
  or (_27256_, _27255_, _12710_);
  or (_27257_, _27256_, _27250_);
  or (_27258_, _27042_, _12226_);
  and (_27259_, _27258_, _10967_);
  and (_27260_, _27259_, _27257_);
  nor (_27261_, _12142_, _10967_);
  or (_27263_, _27261_, _06366_);
  or (_27264_, _27263_, _27260_);
  nand (_27265_, _12288_, _06366_);
  and (_27266_, _27265_, _27264_);
  or (_27267_, _27266_, _06541_);
  nand (_27268_, _12142_, _06541_);
  and (_27269_, _27268_, _05919_);
  and (_27270_, _27269_, _27267_);
  nor (_27271_, _08802_, _05919_);
  or (_27272_, _27271_, _27270_);
  and (_27274_, _27272_, _12724_);
  or (_27275_, _27059_, \oc8051_golden_model_1.PSW [7]);
  or (_27276_, _12141_, _10854_);
  and (_27277_, _27276_, _12723_);
  and (_27278_, _27277_, _27275_);
  or (_27279_, _27278_, _12738_);
  or (_27280_, _27279_, _27274_);
  or (_27281_, _27042_, _12736_);
  and (_27282_, _27281_, _11005_);
  and (_27283_, _27282_, _27280_);
  nor (_27285_, _12142_, _11005_);
  or (_27286_, _27285_, _06383_);
  or (_27287_, _27286_, _27283_);
  nand (_27288_, _12288_, _06383_);
  and (_27289_, _27288_, _27287_);
  or (_27290_, _27289_, _06528_);
  nand (_27291_, _12142_, _06528_);
  and (_27292_, _27291_, _05922_);
  and (_27293_, _27292_, _27290_);
  nor (_27294_, _08802_, _05922_);
  or (_27296_, _27294_, _27293_);
  and (_27297_, _27296_, _12751_);
  or (_27298_, _27059_, _10854_);
  or (_27299_, _12141_, \oc8051_golden_model_1.PSW [7]);
  and (_27300_, _27299_, _12215_);
  and (_27301_, _27300_, _27298_);
  or (_27302_, _27301_, _12758_);
  or (_27303_, _27302_, _27297_);
  or (_27304_, _27042_, _12756_);
  and (_27305_, _27304_, _11051_);
  and (_27307_, _27305_, _27303_);
  nor (_27308_, _12142_, _11051_);
  or (_27309_, _27308_, _11080_);
  or (_27310_, _27309_, _27307_);
  nand (_27311_, _27044_, _11080_);
  and (_27312_, _27311_, _13873_);
  and (_27313_, _27312_, _27310_);
  and (_27314_, _09067_, _06547_);
  or (_27315_, _27314_, _07228_);
  or (_27316_, _27315_, _27313_);
  nand (_27318_, _08802_, _07228_);
  and (_27319_, _27318_, _06946_);
  and (_27320_, _27319_, _27316_);
  or (_27321_, _27052_, _12955_);
  or (_27322_, _12287_, _12954_);
  and (_27323_, _27322_, _06381_);
  and (_27324_, _27323_, _27321_);
  or (_27325_, _27324_, _12774_);
  or (_27326_, _27325_, _27320_);
  or (_27327_, _27042_, _12105_);
  and (_27329_, _27327_, _12963_);
  and (_27330_, _27329_, _27326_);
  nor (_27331_, _12963_, _12142_);
  or (_27332_, _27331_, _10448_);
  or (_27333_, _27332_, _27330_);
  and (_27334_, _27333_, _27047_);
  or (_27335_, _27334_, _06260_);
  or (_27336_, _09067_, _06261_);
  and (_27337_, _27336_, _05924_);
  and (_27338_, _27337_, _27335_);
  nor (_27340_, _08802_, _05924_);
  or (_27341_, _27340_, _06377_);
  or (_27342_, _27341_, _27338_);
  or (_27343_, _27052_, _12954_);
  nand (_27344_, _12288_, _12954_);
  and (_27345_, _27344_, _27343_);
  or (_27346_, _27345_, _06564_);
  and (_27347_, _27346_, _27342_);
  or (_27348_, _27347_, _12985_);
  or (_27349_, _27042_, _12984_);
  and (_27351_, _27349_, _27348_);
  or (_27352_, _27351_, _06563_);
  nand (_27353_, _12142_, _06563_);
  and (_27354_, _27353_, _12991_);
  and (_27355_, _27354_, _27352_);
  nor (_27356_, _27044_, _12991_);
  or (_27357_, _27356_, _07812_);
  or (_27358_, _27357_, _27355_);
  and (_27359_, _27358_, _27046_);
  or (_27360_, _27359_, _06199_);
  or (_27362_, _27345_, _06571_);
  and (_27363_, _27362_, _13006_);
  and (_27364_, _27363_, _27360_);
  nor (_27365_, _27044_, _13006_);
  nor (_27366_, _27365_, _06188_);
  not (_27367_, _27366_);
  nor (_27368_, _27367_, _27364_);
  and (_27369_, _12142_, _06188_);
  nor (_27370_, _27369_, _13014_);
  not (_27371_, _27370_);
  nor (_27373_, _27371_, _27368_);
  or (_27374_, _27373_, _25220_);
  nor (_27375_, _27374_, _27045_);
  or (_27376_, _27375_, _13025_);
  nor (_27377_, _27376_, _27039_);
  and (_27378_, _27042_, _13025_);
  nor (_27379_, _27378_, _27377_);
  nand (_27380_, _27379_, _01452_);
  or (_27381_, _01452_, \oc8051_golden_model_1.PC [6]);
  and (_27382_, _27381_, _43223_);
  and (_43861_, _27382_, _27380_);
  and (_27384_, _08518_, _06188_);
  nor (_27385_, _12091_, \oc8051_golden_model_1.PC [7]);
  nor (_27386_, _27385_, _12092_);
  nor (_27387_, _27386_, _12991_);
  nor (_27388_, _27386_, _12105_);
  nor (_27389_, _27386_, _12756_);
  nor (_27390_, _27386_, _12736_);
  nor (_27391_, _27386_, _12226_);
  nor (_27392_, _27386_, _12232_);
  nor (_27394_, _08972_, _08518_);
  and (_27395_, _08711_, _06241_);
  nor (_27396_, _27386_, _12237_);
  not (_27397_, _27386_);
  and (_27398_, _27397_, _12245_);
  nor (_27399_, _08769_, _07272_);
  and (_27400_, _08711_, _07123_);
  nor (_27401_, _27400_, _06808_);
  and (_27402_, _12419_, \oc8051_golden_model_1.PC [7]);
  or (_27403_, _27402_, _07123_);
  and (_27405_, _27403_, _27401_);
  or (_27406_, _27397_, _12420_);
  nand (_27407_, _27406_, _12427_);
  or (_27408_, _27407_, _27405_);
  and (_27409_, _27408_, _07272_);
  nor (_27410_, _27409_, _27399_);
  nor (_27411_, _27386_, _12427_);
  nor (_27412_, _27411_, _27410_);
  nor (_27413_, _27412_, _08572_);
  or (_27414_, _12137_, _12138_);
  and (_27416_, _27414_, _12181_);
  nor (_27417_, _27414_, _12181_);
  nor (_27418_, _27417_, _27416_);
  nand (_27419_, _27418_, _12414_);
  and (_27420_, _27419_, _08572_);
  or (_27421_, _12414_, _08711_);
  and (_27422_, _27421_, _27420_);
  or (_27423_, _27422_, _27413_);
  nand (_27424_, _27423_, _07338_);
  and (_27425_, _27397_, _07134_);
  nor (_27427_, _27425_, _06251_);
  nand (_27428_, _27427_, _27424_);
  or (_27429_, _12404_, _09363_);
  or (_27430_, _12283_, _12284_);
  and (_27431_, _27430_, _12333_);
  nor (_27432_, _27430_, _12333_);
  nor (_27433_, _27432_, _27431_);
  or (_27434_, _27433_, _12402_);
  and (_27435_, _27434_, _06251_);
  nand (_27436_, _27435_, _27429_);
  and (_27438_, _27436_, _12443_);
  nand (_27439_, _27438_, _27428_);
  nor (_27440_, _27386_, _12443_);
  nor (_27441_, _27440_, _06475_);
  nand (_27442_, _27441_, _27439_);
  and (_27443_, _08518_, _06475_);
  nor (_27444_, _27443_, _07474_);
  nand (_27445_, _27444_, _27442_);
  and (_27446_, _08769_, _07474_);
  nor (_27447_, _27446_, _06468_);
  nand (_27449_, _27447_, _27445_);
  and (_27450_, _08518_, _06468_);
  nor (_27451_, _27450_, _12452_);
  nand (_27452_, _27451_, _27449_);
  nor (_27453_, _27386_, _12451_);
  nor (_27454_, _27453_, _06466_);
  nand (_27455_, _27454_, _27452_);
  and (_27456_, _08518_, _06466_);
  nor (_27457_, _27456_, _12464_);
  nand (_27458_, _27457_, _27455_);
  nor (_27460_, _27386_, _12462_);
  nor (_27461_, _27460_, _06483_);
  nand (_27462_, _27461_, _27458_);
  and (_27463_, _08518_, _06483_);
  nor (_27464_, _27463_, _12466_);
  nand (_27465_, _27464_, _27462_);
  and (_27466_, _08769_, _12466_);
  nor (_27467_, _27466_, _06247_);
  nand (_27468_, _27467_, _27465_);
  and (_27469_, _08518_, _06247_);
  nor (_27471_, _27469_, _12479_);
  and (_27472_, _27471_, _27468_);
  and (_27473_, _12513_, _09363_);
  not (_27474_, _27433_);
  nor (_27475_, _27474_, _12513_);
  or (_27476_, _27475_, _12478_);
  nor (_27477_, _27476_, _27473_);
  nor (_27478_, _27477_, _27472_);
  or (_27479_, _27478_, _06344_);
  nor (_27480_, _27474_, _12392_);
  and (_27482_, _12392_, _09363_);
  or (_27483_, _27482_, _06345_);
  or (_27484_, _27483_, _27480_);
  and (_27485_, _27484_, _27479_);
  or (_27486_, _27485_, _06338_);
  nor (_27487_, _27474_, _12533_);
  and (_27488_, _12533_, _09363_);
  or (_27489_, _27488_, _12536_);
  or (_27490_, _27489_, _27487_);
  and (_27491_, _27490_, _12522_);
  nand (_27493_, _27491_, _27486_);
  nor (_27494_, _27433_, _12555_);
  and (_27495_, _12555_, _12282_);
  or (_27496_, _27495_, _12522_);
  or (_27497_, _27496_, _27494_);
  and (_27498_, _27497_, _12246_);
  and (_27499_, _27498_, _27493_);
  or (_27500_, _27499_, _27398_);
  nand (_27501_, _27500_, _07164_);
  and (_27502_, _08711_, _06461_);
  nor (_27504_, _27502_, _07471_);
  nand (_27505_, _27504_, _27501_);
  nor (_27506_, _08769_, _05947_);
  nor (_27507_, _27506_, _25366_);
  and (_27508_, _27507_, _27505_);
  nor (_27509_, _25365_, _08518_);
  or (_27510_, _27509_, _27508_);
  nand (_27511_, _27510_, _12242_);
  nor (_27512_, _27386_, _12242_);
  nor (_27513_, _27512_, _06505_);
  nand (_27515_, _27513_, _27511_);
  and (_27516_, _08518_, _06505_);
  nor (_27517_, _27516_, _25090_);
  nand (_27518_, _27517_, _27515_);
  and (_27519_, _08769_, _25090_);
  nor (_27520_, _27519_, _06504_);
  nand (_27521_, _27520_, _27518_);
  and (_27522_, _08518_, _06504_);
  nor (_27523_, _27522_, _12582_);
  and (_27524_, _27523_, _27521_);
  or (_27526_, _27524_, _27396_);
  nand (_27527_, _27526_, _12588_);
  nor (_27528_, _12588_, _08518_);
  nor (_27529_, _27528_, _05976_);
  nand (_27530_, _27529_, _27527_);
  and (_27531_, _27386_, _05976_);
  nor (_27532_, _27531_, _06241_);
  and (_27533_, _27532_, _27530_);
  or (_27534_, _27533_, _27395_);
  nand (_27535_, _27534_, _08723_);
  and (_27537_, _08769_, _05970_);
  nor (_27538_, _27537_, _06369_);
  nand (_27539_, _27538_, _27535_);
  and (_27540_, _09363_, _06369_);
  nor (_27541_, _27540_, _12604_);
  nand (_27542_, _27541_, _27539_);
  nor (_27543_, _12603_, _08518_);
  nor (_27544_, _27543_, _05968_);
  nand (_27545_, _27544_, _27542_);
  and (_27546_, _09363_, _05968_);
  nor (_27548_, _27546_, _12615_);
  nand (_27549_, _27548_, _27545_);
  nor (_27550_, _27386_, _12611_);
  nor (_27551_, _27550_, _06332_);
  and (_27552_, _27551_, _27549_);
  and (_27553_, _08518_, _06332_);
  or (_27554_, _27553_, _05900_);
  or (_27555_, _27554_, _27552_);
  and (_27556_, _08769_, _05900_);
  nor (_27557_, _27556_, _12619_);
  nand (_27559_, _27557_, _27555_);
  and (_27560_, _27418_, _12619_);
  nor (_27561_, _27560_, _08973_);
  and (_27562_, _27561_, _27559_);
  or (_27563_, _27562_, _27394_);
  nand (_27564_, _27563_, _07198_);
  and (_27565_, _12282_, _06371_);
  nor (_27566_, _27565_, _10904_);
  nand (_27567_, _27566_, _27564_);
  and (_27568_, _10904_, _08518_);
  nor (_27570_, _27568_, _12634_);
  nand (_27571_, _27570_, _27567_);
  or (_27572_, _12639_, _12638_);
  not (_27573_, _27572_);
  and (_27574_, _27573_, _12658_);
  nor (_27575_, _27573_, _12658_);
  nor (_27576_, _27575_, _27574_);
  and (_27577_, _27576_, _12634_);
  nor (_27578_, _27577_, _06331_);
  and (_27579_, _27578_, _27571_);
  and (_27581_, _08518_, _06331_);
  or (_27582_, _27581_, _05895_);
  or (_27583_, _27582_, _27579_);
  and (_27584_, _08769_, _05895_);
  nor (_27585_, _27584_, _12677_);
  nand (_27586_, _27585_, _27583_);
  and (_27587_, _11291_, _08518_);
  and (_27588_, _27418_, _12684_);
  or (_27589_, _27588_, _27587_);
  and (_27590_, _27589_, _12677_);
  nor (_27592_, _27590_, _12682_);
  and (_27593_, _27592_, _27586_);
  or (_27594_, _27593_, _27392_);
  nand (_27595_, _27594_, _12228_);
  nor (_27596_, _12228_, _08518_);
  nor (_27597_, _27596_, _06367_);
  and (_27598_, _27597_, _27595_);
  and (_27599_, _09363_, _06367_);
  or (_27600_, _27599_, _06533_);
  nor (_27601_, _27600_, _27598_);
  and (_27603_, _08711_, _06533_);
  or (_27604_, _27603_, _27601_);
  nand (_27605_, _27604_, _05890_);
  and (_27606_, _08769_, _05889_);
  nor (_27607_, _27606_, _12701_);
  nand (_27608_, _27607_, _27605_);
  nor (_27609_, _11291_, _08711_);
  and (_27610_, _27418_, _11291_);
  or (_27611_, _27610_, _27609_);
  and (_27612_, _27611_, _12701_);
  nor (_27614_, _27612_, _12710_);
  and (_27615_, _27614_, _27608_);
  or (_27616_, _27615_, _27391_);
  nand (_27617_, _27616_, _10967_);
  nor (_27618_, _10967_, _08518_);
  nor (_27619_, _27618_, _06366_);
  and (_27620_, _27619_, _27617_);
  and (_27621_, _09363_, _06366_);
  or (_27622_, _27621_, _06541_);
  nor (_27623_, _27622_, _27620_);
  and (_27625_, _08711_, _06541_);
  or (_27626_, _27625_, _27623_);
  nand (_27627_, _27626_, _05919_);
  and (_27628_, _08769_, _07209_);
  nor (_27629_, _27628_, _12723_);
  nand (_27630_, _27629_, _27627_);
  nor (_27631_, _27418_, \oc8051_golden_model_1.PSW [7]);
  nor (_27632_, _08518_, _10854_);
  nor (_27633_, _27632_, _12724_);
  not (_27634_, _27633_);
  nor (_27636_, _27634_, _27631_);
  nor (_27637_, _27636_, _12738_);
  and (_27638_, _27637_, _27630_);
  or (_27639_, _27638_, _27390_);
  nand (_27640_, _27639_, _11005_);
  nor (_27641_, _11005_, _08518_);
  nor (_27642_, _27641_, _06383_);
  and (_27643_, _27642_, _27640_);
  and (_27644_, _09363_, _06383_);
  or (_27645_, _27644_, _06528_);
  nor (_27647_, _27645_, _27643_);
  and (_27648_, _08711_, _06528_);
  or (_27649_, _27648_, _27647_);
  nand (_27650_, _27649_, _05922_);
  and (_27651_, _08769_, _12746_);
  nor (_27652_, _27651_, _12215_);
  nand (_27653_, _27652_, _27650_);
  and (_27654_, _08518_, _10854_);
  and (_27655_, _27418_, \oc8051_golden_model_1.PSW [7]);
  or (_27656_, _27655_, _27654_);
  and (_27658_, _27656_, _12215_);
  nor (_27659_, _27658_, _12758_);
  and (_27660_, _27659_, _27653_);
  or (_27661_, _27660_, _27389_);
  nand (_27662_, _27661_, _11051_);
  nor (_27663_, _11051_, _08518_);
  nor (_27664_, _27663_, _11080_);
  and (_27665_, _27664_, _27662_);
  and (_27666_, _27386_, _11080_);
  or (_27667_, _27666_, _06547_);
  nor (_27669_, _27667_, _27665_);
  nor (_27670_, _08671_, _13873_);
  or (_27671_, _27670_, _27669_);
  nand (_27672_, _27671_, _05916_);
  and (_27673_, _08769_, _07228_);
  nor (_27674_, _27673_, _06381_);
  nand (_27675_, _27674_, _27672_);
  and (_27676_, _27474_, _12954_);
  nor (_27677_, _12954_, _09363_);
  or (_27678_, _27677_, _06946_);
  or (_27680_, _27678_, _27676_);
  and (_27681_, _27680_, _12105_);
  and (_27682_, _27681_, _27675_);
  or (_27683_, _27682_, _27388_);
  nand (_27684_, _27683_, _12963_);
  nor (_27685_, _12963_, _08518_);
  nor (_27686_, _27685_, _10448_);
  nand (_27687_, _27686_, _27684_);
  and (_27688_, _27386_, _10448_);
  nor (_27689_, _27688_, _06260_);
  and (_27691_, _27689_, _27687_);
  nor (_27692_, _08671_, _06261_);
  or (_27693_, _27692_, _27691_);
  nand (_27694_, _27693_, _05924_);
  and (_27695_, _08769_, _12089_);
  nor (_27696_, _27695_, _06377_);
  nand (_27697_, _27696_, _27694_);
  and (_27698_, _12954_, _12282_);
  nor (_27699_, _27433_, _12954_);
  nor (_27700_, _27699_, _27698_);
  and (_27702_, _27700_, _06377_);
  nor (_27703_, _27702_, _12985_);
  nand (_27704_, _27703_, _27697_);
  nor (_27705_, _27386_, _12984_);
  nor (_27706_, _27705_, _06563_);
  nand (_27707_, _27706_, _27704_);
  and (_27708_, _08518_, _06563_);
  nor (_27709_, _27708_, _12992_);
  and (_27710_, _27709_, _27707_);
  or (_27711_, _27710_, _27387_);
  nand (_27713_, _27711_, _07250_);
  and (_27714_, _08769_, _07812_);
  nor (_27715_, _27714_, _06199_);
  nand (_27716_, _27715_, _27713_);
  and (_27717_, _27700_, _06199_);
  nor (_27718_, _27717_, _13007_);
  nand (_27719_, _27718_, _27716_);
  nor (_27720_, _27386_, _13006_);
  nor (_27721_, _27720_, _06188_);
  and (_27722_, _27721_, _27719_);
  or (_27724_, _27722_, _27384_);
  nand (_27725_, _27724_, _13013_);
  nor (_27726_, _27397_, _13013_);
  nor (_27727_, _27726_, _25220_);
  nand (_27728_, _27727_, _27725_);
  and (_27729_, _25220_, _08769_);
  nor (_27730_, _27729_, _13025_);
  and (_27731_, _27730_, _27728_);
  and (_27732_, _27386_, _13025_);
  or (_27733_, _27732_, _27731_);
  or (_27735_, _27733_, _01456_);
  or (_27736_, _01452_, \oc8051_golden_model_1.PC [7]);
  and (_27737_, _27736_, _43223_);
  and (_43862_, _27737_, _27735_);
  and (_27738_, _06799_, _06342_);
  and (_27739_, _06799_, _06378_);
  and (_27740_, _12280_, _06366_);
  nor (_27741_, _12185_, _08972_);
  nor (_27742_, _12619_, _05900_);
  not (_27743_, _27742_);
  and (_27745_, _12185_, _06332_);
  nor (_27746_, _12092_, \oc8051_golden_model_1.PC [8]);
  nor (_27747_, _27746_, _12093_);
  nor (_27748_, _27747_, _12611_);
  and (_27749_, _12279_, _05968_);
  and (_27750_, _12185_, _06483_);
  and (_27751_, _12185_, _06475_);
  and (_27752_, _12427_, _12419_);
  or (_27753_, _27752_, _27747_);
  not (_27754_, _12185_);
  nand (_27756_, _27754_, _07123_);
  and (_27757_, _27756_, _12418_);
  nor (_27758_, _07123_, \oc8051_golden_model_1.PC [8]);
  nand (_27759_, _27758_, _12419_);
  nand (_27760_, _27759_, _27757_);
  nand (_27761_, _27760_, _25018_);
  and (_27762_, _27761_, _27753_);
  and (_27763_, _27747_, _06808_);
  or (_27764_, _27763_, _08572_);
  or (_27765_, _27764_, _27762_);
  nor (_27767_, _12188_, _12183_);
  nor (_27768_, _27767_, _12189_);
  and (_27769_, _27768_, _12414_);
  or (_27770_, _27769_, _08573_);
  and (_27771_, _12412_, _12185_);
  or (_27772_, _27771_, _27770_);
  and (_27773_, _27772_, _27765_);
  or (_27774_, _27773_, _07134_);
  not (_27775_, _27747_);
  nand (_27776_, _27775_, _07134_);
  and (_27778_, _27776_, _06252_);
  and (_27779_, _27778_, _27774_);
  nor (_27780_, _12337_, _12335_);
  nor (_27781_, _27780_, _12338_);
  or (_27782_, _27781_, _12402_);
  and (_27783_, _27782_, _06251_);
  or (_27784_, _12404_, _12279_);
  and (_27785_, _27784_, _27783_);
  or (_27786_, _27785_, _12444_);
  or (_27787_, _27786_, _27779_);
  or (_27789_, _27747_, _12443_);
  and (_27790_, _27789_, _06476_);
  and (_27791_, _27790_, _27787_);
  or (_27792_, _27791_, _27751_);
  and (_27793_, _27792_, _12446_);
  nand (_27794_, _12185_, _06468_);
  nand (_27795_, _27794_, _12451_);
  or (_27796_, _27795_, _27793_);
  or (_27797_, _27747_, _12451_);
  and (_27798_, _27797_, _06801_);
  and (_27800_, _27798_, _27796_);
  nand (_27801_, _12185_, _06466_);
  nand (_27802_, _27801_, _12462_);
  or (_27803_, _27802_, _27800_);
  or (_27804_, _27747_, _12462_);
  and (_27805_, _27804_, _06484_);
  and (_27806_, _27805_, _27803_);
  or (_27807_, _27806_, _27750_);
  and (_27808_, _27807_, _12467_);
  nand (_27809_, _12185_, _06247_);
  nand (_27811_, _27809_, _12478_);
  or (_27812_, _27811_, _27808_);
  and (_27813_, _12513_, _12279_);
  not (_27814_, _27781_);
  nor (_27815_, _27814_, _12513_);
  or (_27816_, _27815_, _27813_);
  or (_27817_, _27816_, _12478_);
  and (_27818_, _27817_, _27812_);
  or (_27819_, _27818_, _06344_);
  nor (_27820_, _27814_, _12392_);
  and (_27822_, _12392_, _12279_);
  or (_27823_, _27822_, _06345_);
  or (_27824_, _27823_, _27820_);
  and (_27825_, _27824_, _27819_);
  or (_27826_, _27825_, _06338_);
  nor (_27827_, _27814_, _12533_);
  and (_27828_, _12533_, _12279_);
  or (_27829_, _27828_, _12536_);
  or (_27830_, _27829_, _27827_);
  and (_27831_, _27830_, _12522_);
  and (_27833_, _27831_, _27826_);
  or (_27834_, _27781_, _12555_);
  nand (_27835_, _12555_, _12280_);
  and (_27836_, _27835_, _06373_);
  and (_27837_, _27836_, _27834_);
  or (_27838_, _27837_, _12245_);
  or (_27839_, _27838_, _27833_);
  nand (_27840_, _27775_, _12245_);
  and (_27841_, _27840_, _07164_);
  and (_27842_, _27841_, _27839_);
  and (_27844_, _12185_, _06461_);
  or (_27845_, _27844_, _07471_);
  or (_27846_, _27845_, _27842_);
  and (_27847_, _27846_, _25365_);
  nor (_27848_, _25365_, _27754_);
  or (_27849_, _27848_, _12243_);
  or (_27850_, _27849_, _27847_);
  or (_27851_, _27747_, _12242_);
  and (_27852_, _27851_, _14007_);
  and (_27853_, _27852_, _27850_);
  and (_27854_, _12185_, _06505_);
  or (_27855_, _27854_, _25090_);
  or (_27856_, _27855_, _27853_);
  and (_27857_, _27856_, _14006_);
  nand (_27858_, _12185_, _06504_);
  nand (_27859_, _27858_, _12237_);
  or (_27860_, _27859_, _27857_);
  or (_27861_, _27747_, _12237_);
  and (_27862_, _27861_, _12588_);
  and (_27863_, _27862_, _27860_);
  nor (_27866_, _12588_, _27754_);
  or (_27867_, _27866_, _05976_);
  or (_27868_, _27867_, _27863_);
  nand (_27869_, _27775_, _05976_);
  and (_27870_, _27869_, _27868_);
  or (_27871_, _27870_, _06241_);
  nand (_27872_, _27754_, _06241_);
  nor (_27873_, _06369_, _05970_);
  and (_27874_, _27873_, _27872_);
  and (_27875_, _27874_, _27871_);
  and (_27877_, _12279_, _06369_);
  or (_27878_, _27877_, _12604_);
  nor (_27879_, _27878_, _27875_);
  nor (_27880_, _12603_, _12185_);
  nor (_27881_, _27880_, _05968_);
  not (_27882_, _27881_);
  nor (_27883_, _27882_, _27879_);
  or (_27884_, _27883_, _12615_);
  nor (_27885_, _27884_, _27749_);
  or (_27886_, _27885_, _06332_);
  nor (_27888_, _27886_, _27748_);
  nor (_27889_, _27888_, _27745_);
  nor (_27890_, _27889_, _27743_);
  and (_27891_, _27768_, _12619_);
  nor (_27892_, _27891_, _08973_);
  not (_27893_, _27892_);
  nor (_27894_, _27893_, _27890_);
  or (_27895_, _27894_, _27741_);
  nand (_27896_, _27895_, _07198_);
  and (_27897_, _12280_, _06371_);
  nor (_27899_, _27897_, _10904_);
  nand (_27900_, _27899_, _27896_);
  and (_27901_, _12185_, _10904_);
  nor (_27902_, _27901_, _12634_);
  nand (_27903_, _27902_, _27900_);
  and (_27904_, _12660_, _12637_);
  nor (_27905_, _27904_, _12661_);
  nor (_27906_, _27905_, _12635_);
  nor (_27907_, _27906_, _06331_);
  nand (_27908_, _27907_, _27903_);
  and (_27910_, _12185_, _06331_);
  nor (_27911_, _27910_, _05895_);
  nand (_27912_, _27911_, _27908_);
  nand (_27913_, _27912_, _12678_);
  and (_27914_, _12185_, _11291_);
  and (_27915_, _27768_, _12684_);
  or (_27916_, _27915_, _27914_);
  and (_27917_, _27916_, _12677_);
  nor (_27918_, _27917_, _12682_);
  nand (_27919_, _27918_, _27913_);
  nor (_27921_, _27747_, _12232_);
  nor (_27922_, _27921_, _12229_);
  nand (_27923_, _27922_, _27919_);
  nor (_27924_, _27754_, _12228_);
  nor (_27925_, _27924_, _06367_);
  nand (_27926_, _27925_, _27923_);
  and (_27927_, _12280_, _06367_);
  nor (_27928_, _27927_, _06533_);
  nand (_27929_, _27928_, _27926_);
  and (_27930_, _12185_, _06533_);
  nor (_27932_, _27930_, _05889_);
  nand (_27933_, _27932_, _27929_);
  nand (_27934_, _27933_, _12702_);
  nor (_27935_, _27754_, _11291_);
  and (_27936_, _27768_, _11291_);
  or (_27937_, _27936_, _27935_);
  and (_27938_, _27937_, _12701_);
  nor (_27939_, _27938_, _12710_);
  nand (_27940_, _27939_, _27934_);
  nor (_27941_, _27747_, _12226_);
  nor (_27943_, _27941_, _10968_);
  nand (_27944_, _27943_, _27940_);
  nor (_27945_, _27754_, _10967_);
  nor (_27946_, _27945_, _06366_);
  and (_27947_, _27946_, _27944_);
  or (_27948_, _27947_, _27740_);
  nand (_27949_, _27948_, _07210_);
  and (_27950_, _27754_, _06541_);
  not (_27951_, _27950_);
  nor (_27952_, _12723_, _07209_);
  and (_27954_, _27952_, _27951_);
  nand (_27955_, _27954_, _27949_);
  nor (_27956_, _27768_, \oc8051_golden_model_1.PSW [7]);
  nor (_27957_, _12185_, _10854_);
  nor (_27958_, _27957_, _12724_);
  not (_27959_, _27958_);
  nor (_27960_, _27959_, _27956_);
  nor (_27961_, _27960_, _12738_);
  nand (_27962_, _27961_, _27955_);
  nor (_27963_, _27747_, _12736_);
  nor (_27965_, _27963_, _11006_);
  and (_27966_, _27965_, _27962_);
  nor (_27967_, _27754_, _11005_);
  or (_27968_, _27967_, _27966_);
  and (_27969_, _27968_, _07231_);
  and (_27970_, _12279_, _06383_);
  or (_27971_, _27970_, _06528_);
  or (_27972_, _27971_, _27969_);
  and (_27973_, _27754_, _06528_);
  not (_27974_, _27973_);
  nor (_27976_, _12215_, _12746_);
  and (_27977_, _27976_, _27974_);
  nand (_27978_, _27977_, _27972_);
  and (_27979_, _12185_, _10854_);
  and (_27980_, _27768_, \oc8051_golden_model_1.PSW [7]);
  or (_27981_, _27980_, _27979_);
  and (_27982_, _27981_, _12215_);
  nor (_27983_, _27982_, _12758_);
  nand (_27984_, _27983_, _27978_);
  nor (_27985_, _27747_, _12756_);
  nor (_27987_, _27985_, _11052_);
  and (_27988_, _27987_, _27984_);
  nor (_27989_, _27754_, _11051_);
  or (_27990_, _27989_, _11080_);
  or (_27991_, _27990_, _27988_);
  and (_27992_, _27775_, _11080_);
  nor (_27993_, _27992_, _06547_);
  nand (_27994_, _27993_, _27991_);
  and (_27995_, _07325_, _06547_);
  nor (_27996_, _27995_, _07228_);
  nand (_27998_, _27996_, _27994_);
  nand (_27999_, _27998_, _06946_);
  and (_28000_, _27814_, _12954_);
  nor (_28001_, _12279_, _12954_);
  or (_28002_, _28001_, _06946_);
  or (_28003_, _28002_, _28000_);
  and (_28004_, _28003_, _12105_);
  nand (_28005_, _28004_, _27999_);
  nor (_28006_, _27747_, _12105_);
  nor (_28007_, _28006_, _12964_);
  and (_28009_, _28007_, _28005_);
  nor (_28010_, _12963_, _27754_);
  or (_28011_, _28010_, _10448_);
  or (_28012_, _28011_, _28009_);
  and (_28013_, _27775_, _10448_);
  nor (_28014_, _28013_, _06260_);
  nand (_28015_, _28014_, _28012_);
  and (_28016_, _07325_, _06260_);
  nor (_28017_, _28016_, _12089_);
  nand (_28018_, _28017_, _28015_);
  nand (_28020_, _28018_, _06564_);
  and (_28021_, _12280_, _12954_);
  nor (_28022_, _27781_, _12954_);
  nor (_28023_, _28022_, _28021_);
  and (_28024_, _28023_, _06377_);
  nor (_28025_, _28024_, _12985_);
  nand (_28026_, _28025_, _28020_);
  nor (_28027_, _27747_, _12984_);
  nor (_28028_, _28027_, _06563_);
  nand (_28029_, _28028_, _28026_);
  and (_28031_, _12185_, _06563_);
  nor (_28032_, _28031_, _12992_);
  nand (_28033_, _28032_, _28029_);
  nor (_28034_, _27747_, _12991_);
  nor (_28035_, _28034_, _06378_);
  and (_28036_, _28035_, _28033_);
  or (_28037_, _28036_, _27739_);
  nor (_28038_, _05912_, _06199_);
  nand (_28039_, _28038_, _28037_);
  and (_28040_, _28023_, _06199_);
  nor (_28042_, _28040_, _13007_);
  nand (_28043_, _28042_, _28039_);
  nor (_28044_, _27747_, _13006_);
  nor (_28045_, _28044_, _06188_);
  nand (_28046_, _28045_, _28043_);
  and (_28047_, _12185_, _06188_);
  nor (_28048_, _28047_, _13014_);
  nand (_28049_, _28048_, _28046_);
  nor (_28050_, _27747_, _13013_);
  nor (_28051_, _28050_, _06342_);
  and (_28053_, _28051_, _28049_);
  or (_28054_, _28053_, _27738_);
  nor (_28055_, _13025_, _05907_);
  and (_28056_, _28055_, _28054_);
  and (_28057_, _27747_, _13025_);
  or (_28058_, _28057_, _28056_);
  or (_28059_, _28058_, _01456_);
  or (_28060_, _01452_, \oc8051_golden_model_1.PC [8]);
  and (_28061_, _28060_, _43223_);
  and (_43863_, _28061_, _28059_);
  nor (_28063_, _06155_, _13018_);
  nor (_28064_, _06155_, _08505_);
  nor (_28065_, _12093_, \oc8051_golden_model_1.PC [9]);
  nor (_28066_, _28065_, _12094_);
  nor (_28067_, _28066_, _12105_);
  nor (_28068_, _28066_, _12756_);
  and (_28069_, _12274_, _06383_);
  nor (_28070_, _28066_, _12736_);
  and (_28071_, _12274_, _06366_);
  nor (_28072_, _28066_, _12226_);
  and (_28074_, _12274_, _06367_);
  nor (_28075_, _28066_, _12232_);
  nor (_28076_, _12133_, _08972_);
  and (_28077_, _12133_, _06332_);
  and (_28078_, _12133_, _06504_);
  nor (_28079_, _06504_, _25090_);
  not (_28080_, _28066_);
  and (_28081_, _28080_, _12245_);
  or (_28082_, _12277_, _12276_);
  not (_28083_, _28082_);
  nor (_28085_, _28083_, _12339_);
  and (_28086_, _28083_, _12339_);
  nor (_28087_, _28086_, _28085_);
  nor (_28088_, _28087_, _12533_);
  and (_28089_, _12533_, _12274_);
  nor (_28090_, _28089_, _28088_);
  or (_28091_, _28090_, _12536_);
  and (_28092_, _12392_, _12274_);
  nor (_28093_, _28087_, _12392_);
  or (_28094_, _28093_, _28092_);
  nor (_28096_, _28094_, _06345_);
  and (_28097_, _28087_, _12404_);
  and (_28098_, _12402_, _12275_);
  nor (_28099_, _28098_, _28097_);
  or (_28100_, _28099_, _06252_);
  and (_28101_, _12412_, _12133_);
  not (_28102_, _28101_);
  nor (_28103_, _12189_, _12186_);
  and (_28104_, _28103_, _12136_);
  nor (_28105_, _28103_, _12136_);
  nor (_28107_, _28105_, _28104_);
  nor (_28108_, _28107_, _12412_);
  nor (_28109_, _28108_, _08573_);
  and (_28110_, _28109_, _28102_);
  and (_28111_, _28066_, _06808_);
  or (_28112_, _28066_, _27752_);
  not (_28113_, _12133_);
  and (_28114_, _28113_, _07123_);
  nor (_28115_, _28114_, _06808_);
  nor (_28116_, _07123_, \oc8051_golden_model_1.PC [9]);
  nand (_28118_, _28116_, _12419_);
  nand (_28119_, _28118_, _28115_);
  nand (_28120_, _28119_, _25018_);
  and (_28121_, _28120_, _28112_);
  or (_28122_, _28121_, _08572_);
  nor (_28123_, _28122_, _28111_);
  or (_28124_, _28123_, _07134_);
  nor (_28125_, _28124_, _28110_);
  and (_28126_, _28066_, _07134_);
  or (_28127_, _28126_, _06251_);
  or (_28129_, _28127_, _28125_);
  and (_28130_, _28129_, _28100_);
  nor (_28131_, _28130_, _12444_);
  nor (_28132_, _28066_, _12443_);
  nor (_28133_, _28132_, _06475_);
  not (_28134_, _28133_);
  or (_28135_, _28134_, _28131_);
  and (_28136_, _12133_, _06475_);
  nor (_28137_, _28136_, _07474_);
  nand (_28138_, _28137_, _28135_);
  nand (_28140_, _28138_, _07142_);
  and (_28141_, _12133_, _06468_);
  nor (_28142_, _28141_, _12452_);
  nand (_28143_, _28142_, _28140_);
  nor (_28144_, _28066_, _12451_);
  nor (_28145_, _28144_, _06466_);
  nand (_28146_, _28145_, _28143_);
  and (_28147_, _12133_, _06466_);
  nor (_28148_, _28147_, _12464_);
  nand (_28149_, _28148_, _28146_);
  nor (_28151_, _28066_, _12462_);
  nor (_28152_, _28151_, _06483_);
  nand (_28153_, _28152_, _28149_);
  and (_28154_, _12133_, _06483_);
  nor (_28155_, _28154_, _12466_);
  nand (_28156_, _28155_, _28153_);
  nand (_28157_, _28156_, _07523_);
  and (_28158_, _12133_, _06247_);
  nor (_28159_, _28158_, _12479_);
  and (_28160_, _28159_, _28157_);
  and (_28161_, _12513_, _12274_);
  nor (_28162_, _28087_, _12513_);
  or (_28163_, _28162_, _28161_);
  nor (_28164_, _28163_, _12478_);
  or (_28165_, _28164_, _28160_);
  and (_28166_, _28165_, _06345_);
  or (_28167_, _28166_, _28096_);
  or (_28168_, _28167_, _06338_);
  and (_28169_, _28168_, _28091_);
  or (_28170_, _28169_, _06373_);
  and (_28173_, _12555_, _12274_);
  nor (_28174_, _28087_, _12555_);
  or (_28175_, _28174_, _28173_);
  and (_28176_, _28175_, _06373_);
  nor (_28177_, _28176_, _12245_);
  and (_28178_, _28177_, _28170_);
  or (_28179_, _28178_, _28081_);
  nand (_28180_, _28179_, _07164_);
  and (_28181_, _28113_, _06461_);
  and (_28182_, _25365_, _05947_);
  not (_28184_, _28182_);
  nor (_28185_, _28184_, _28181_);
  nand (_28186_, _28185_, _28180_);
  nor (_28187_, _25365_, _28113_);
  nor (_28188_, _28187_, _12243_);
  nand (_28189_, _28188_, _28186_);
  nor (_28190_, _28066_, _12242_);
  nor (_28191_, _28190_, _06505_);
  and (_28192_, _28191_, _28189_);
  and (_28193_, _12133_, _06505_);
  or (_28195_, _28193_, _28192_);
  and (_28196_, _28195_, _28079_);
  or (_28197_, _28196_, _28078_);
  nand (_28198_, _28197_, _12237_);
  nor (_28199_, _28080_, _12237_);
  nor (_28200_, _28199_, _12589_);
  nand (_28201_, _28200_, _28198_);
  nor (_28202_, _12588_, _12133_);
  nor (_28203_, _28202_, _05976_);
  nand (_28204_, _28203_, _28201_);
  and (_28206_, _28066_, _05976_);
  nor (_28207_, _28206_, _06241_);
  nand (_28208_, _28207_, _28204_);
  not (_28209_, _27873_);
  and (_28210_, _28113_, _06241_);
  nor (_28211_, _28210_, _28209_);
  nand (_28212_, _28211_, _28208_);
  and (_28213_, _12274_, _06369_);
  nor (_28214_, _28213_, _12604_);
  nand (_28215_, _28214_, _28212_);
  nor (_28217_, _12603_, _12133_);
  nor (_28218_, _28217_, _05968_);
  nand (_28219_, _28218_, _28215_);
  and (_28220_, _12274_, _05968_);
  nor (_28221_, _28220_, _12615_);
  nand (_28222_, _28221_, _28219_);
  nor (_28223_, _28066_, _12611_);
  nor (_28224_, _28223_, _06332_);
  and (_28225_, _28224_, _28222_);
  or (_28226_, _28225_, _28077_);
  nand (_28228_, _28226_, _27742_);
  nor (_28229_, _28107_, _12620_);
  nor (_28230_, _28229_, _08973_);
  and (_28231_, _28230_, _28228_);
  or (_28232_, _28231_, _28076_);
  nand (_28233_, _28232_, _07198_);
  and (_28234_, _12275_, _06371_);
  nor (_28235_, _28234_, _10904_);
  nand (_28236_, _28235_, _28233_);
  and (_28237_, _12133_, _10904_);
  nor (_28239_, _28237_, _12634_);
  nand (_28240_, _28239_, _28236_);
  nor (_28241_, _12661_, \oc8051_golden_model_1.DPH [1]);
  nor (_28242_, _28241_, _12662_);
  nor (_28243_, _28242_, _12635_);
  nor (_28244_, _28243_, _06331_);
  nand (_28245_, _28244_, _28240_);
  and (_28246_, _12133_, _06331_);
  nor (_28247_, _28246_, _05895_);
  nand (_28248_, _28247_, _28245_);
  nand (_28250_, _28248_, _12678_);
  and (_28251_, _12133_, _11291_);
  nor (_28252_, _28107_, _11291_);
  or (_28253_, _28252_, _28251_);
  and (_28254_, _28253_, _12677_);
  nor (_28255_, _28254_, _12682_);
  and (_28256_, _28255_, _28250_);
  or (_28257_, _28256_, _28075_);
  nand (_28258_, _28257_, _12228_);
  nor (_28259_, _12133_, _12228_);
  nor (_28261_, _28259_, _06367_);
  and (_28262_, _28261_, _28258_);
  or (_28263_, _28262_, _28074_);
  nand (_28264_, _28263_, _07216_);
  and (_28265_, _12133_, _06533_);
  nor (_28266_, _28265_, _05889_);
  nand (_28267_, _28266_, _28264_);
  nand (_28268_, _28267_, _12702_);
  and (_28269_, _28107_, _11291_);
  nor (_28270_, _12133_, _11291_);
  nor (_28272_, _28270_, _12702_);
  not (_28273_, _28272_);
  nor (_28274_, _28273_, _28269_);
  nor (_28275_, _28274_, _12710_);
  and (_28276_, _28275_, _28268_);
  or (_28277_, _28276_, _28072_);
  nand (_28278_, _28277_, _10967_);
  nor (_28279_, _12133_, _10967_);
  nor (_28280_, _28279_, _06366_);
  and (_28281_, _28280_, _28278_);
  or (_28283_, _28281_, _28071_);
  nand (_28284_, _28283_, _07210_);
  and (_28285_, _12133_, _06541_);
  nor (_28286_, _28285_, _07209_);
  nand (_28287_, _28286_, _28284_);
  nand (_28288_, _28287_, _12724_);
  and (_28289_, _12133_, \oc8051_golden_model_1.PSW [7]);
  nor (_28290_, _28107_, \oc8051_golden_model_1.PSW [7]);
  or (_28291_, _28290_, _28289_);
  and (_28292_, _28291_, _12723_);
  nor (_28294_, _28292_, _12738_);
  and (_28295_, _28294_, _28288_);
  or (_28296_, _28295_, _28070_);
  nand (_28297_, _28296_, _11005_);
  nor (_28298_, _12133_, _11005_);
  nor (_28299_, _28298_, _06383_);
  and (_28300_, _28299_, _28297_);
  or (_28301_, _28300_, _28069_);
  nand (_28302_, _28301_, _07229_);
  and (_28303_, _12133_, _06528_);
  nor (_28305_, _28303_, _12746_);
  nand (_28306_, _28305_, _28302_);
  nand (_28307_, _28306_, _12751_);
  and (_28308_, _12133_, _10854_);
  nor (_28309_, _28107_, _10854_);
  or (_28310_, _28309_, _28308_);
  and (_28311_, _28310_, _12215_);
  nor (_28312_, _28311_, _12758_);
  and (_28313_, _28312_, _28307_);
  or (_28314_, _28313_, _28068_);
  nand (_28316_, _28314_, _11051_);
  nor (_28317_, _12133_, _11051_);
  nor (_28318_, _28317_, _11080_);
  nand (_28319_, _28318_, _28316_);
  and (_28320_, _28066_, _11080_);
  nor (_28321_, _28320_, _06547_);
  nand (_28322_, _28321_, _28319_);
  nor (_28323_, _06381_, _07228_);
  not (_28324_, _28323_);
  and (_28325_, _07120_, _06547_);
  nor (_28327_, _28325_, _28324_);
  nand (_28328_, _28327_, _28322_);
  and (_28329_, _28087_, _12954_);
  nor (_28330_, _12274_, _12954_);
  or (_28331_, _28330_, _06946_);
  or (_28332_, _28331_, _28329_);
  and (_28333_, _28332_, _12105_);
  and (_28334_, _28333_, _28328_);
  or (_28335_, _28334_, _28067_);
  nand (_28336_, _28335_, _12963_);
  nor (_28338_, _12963_, _12133_);
  nor (_28339_, _28338_, _10448_);
  nand (_28340_, _28339_, _28336_);
  and (_28341_, _28066_, _10448_);
  nor (_28342_, _28341_, _06260_);
  nand (_28343_, _28342_, _28340_);
  nor (_28344_, _06377_, _12089_);
  not (_28345_, _28344_);
  and (_28346_, _07120_, _06260_);
  nor (_28347_, _28346_, _28345_);
  nand (_28349_, _28347_, _28343_);
  and (_28350_, _12274_, _12954_);
  nor (_28351_, _28087_, _12954_);
  or (_28352_, _28351_, _28350_);
  and (_28353_, _28352_, _06377_);
  nor (_28354_, _28353_, _12985_);
  nand (_28355_, _28354_, _28349_);
  nor (_28356_, _28066_, _12984_);
  nor (_28357_, _28356_, _06563_);
  nand (_28358_, _28357_, _28355_);
  and (_28360_, _12133_, _06563_);
  nor (_28361_, _28360_, _12992_);
  nand (_28362_, _28361_, _28358_);
  nor (_28363_, _28066_, _12991_);
  nor (_28364_, _28363_, _06378_);
  and (_28365_, _28364_, _28362_);
  or (_28366_, _28365_, _28064_);
  nand (_28367_, _28366_, _28038_);
  and (_28368_, _28352_, _06199_);
  nor (_28369_, _28368_, _13007_);
  nand (_28371_, _28369_, _28367_);
  nor (_28372_, _28066_, _13006_);
  nor (_28373_, _28372_, _06188_);
  nand (_28374_, _28373_, _28371_);
  and (_28375_, _12133_, _06188_);
  nor (_28376_, _28375_, _13014_);
  nand (_28377_, _28376_, _28374_);
  nor (_28378_, _28066_, _13013_);
  nor (_28379_, _28378_, _06342_);
  and (_28380_, _28379_, _28377_);
  or (_28382_, _28380_, _28063_);
  and (_28383_, _28382_, _28055_);
  and (_28384_, _28066_, _13025_);
  or (_28385_, _28384_, _28383_);
  or (_28386_, _28385_, _01456_);
  or (_28387_, _01452_, \oc8051_golden_model_1.PC [9]);
  and (_28388_, _28387_, _43223_);
  and (_43864_, _28388_, _28386_);
  nor (_28389_, _12094_, \oc8051_golden_model_1.PC [10]);
  nor (_28390_, _28389_, _12095_);
  or (_28392_, _28390_, _12984_);
  or (_28393_, _28390_, _12966_);
  or (_28394_, _28390_, _11081_);
  nand (_28395_, _12269_, _06383_);
  nand (_28396_, _12269_, _06366_);
  or (_28397_, _25365_, _12127_);
  nor (_28398_, _12342_, _12272_);
  nor (_28399_, _28398_, _12343_);
  or (_28400_, _28399_, _12392_);
  nand (_28401_, _12392_, _12269_);
  and (_28403_, _28401_, _28400_);
  or (_28404_, _28403_, _06345_);
  not (_28405_, _12127_);
  nand (_28406_, _28405_, _06466_);
  and (_28407_, _12127_, _07123_);
  and (_28408_, _07124_, \oc8051_golden_model_1.PC [10]);
  and (_28409_, _28408_, _12419_);
  or (_28410_, _28409_, _28407_);
  and (_28411_, _28410_, _12418_);
  or (_28412_, _28411_, _06705_);
  and (_28414_, _28412_, _12427_);
  and (_28415_, _12427_, _12420_);
  not (_28416_, _28415_);
  and (_28417_, _28416_, _28390_);
  or (_28418_, _28417_, _08572_);
  or (_28419_, _28418_, _28414_);
  nor (_28420_, _12193_, _12190_);
  not (_28421_, _28420_);
  and (_28422_, _28421_, _12130_);
  nor (_28423_, _28421_, _12130_);
  nor (_28425_, _28423_, _28422_);
  and (_28426_, _28425_, _12414_);
  and (_28427_, _12412_, _12127_);
  or (_28428_, _28427_, _28426_);
  or (_28429_, _28428_, _08573_);
  and (_28430_, _28429_, _28419_);
  or (_28431_, _28430_, _07134_);
  or (_28432_, _28390_, _07338_);
  and (_28433_, _28432_, _06252_);
  and (_28434_, _28433_, _28431_);
  or (_28436_, _28399_, _12402_);
  or (_28437_, _12404_, _12268_);
  and (_28438_, _28437_, _06251_);
  and (_28439_, _28438_, _28436_);
  or (_28440_, _28439_, _12444_);
  or (_28441_, _28440_, _28434_);
  or (_28442_, _28390_, _12443_);
  and (_28443_, _28442_, _06476_);
  and (_28444_, _28443_, _28441_);
  and (_28445_, _12446_, _28405_);
  nor (_28447_, _28445_, _12447_);
  or (_28448_, _28447_, _28444_);
  nand (_28449_, _28405_, _06468_);
  and (_28450_, _28449_, _12451_);
  and (_28451_, _28450_, _28448_);
  and (_28452_, _28390_, _12452_);
  or (_28453_, _28452_, _06466_);
  or (_28454_, _28453_, _28451_);
  and (_28455_, _28454_, _28406_);
  or (_28456_, _28455_, _12464_);
  or (_28458_, _28390_, _12462_);
  and (_28459_, _28458_, _06484_);
  and (_28460_, _28459_, _28456_);
  and (_28461_, _12127_, _06483_);
  or (_28462_, _28461_, _12466_);
  or (_28463_, _28462_, _28460_);
  and (_28464_, _28463_, _07523_);
  nand (_28465_, _12127_, _06247_);
  nand (_28466_, _28465_, _12478_);
  or (_28467_, _28466_, _28464_);
  or (_28469_, _28399_, _12513_);
  nand (_28470_, _12513_, _12269_);
  and (_28471_, _28470_, _28469_);
  or (_28472_, _28471_, _12478_);
  and (_28473_, _28472_, _28467_);
  or (_28474_, _28473_, _06344_);
  and (_28475_, _28474_, _28404_);
  or (_28476_, _28475_, _06338_);
  and (_28477_, _12533_, _12268_);
  and (_28478_, _28399_, _12534_);
  or (_28480_, _28478_, _12536_);
  or (_28481_, _28480_, _28477_);
  and (_28482_, _28481_, _12522_);
  and (_28483_, _28482_, _28476_);
  or (_28484_, _28399_, _12555_);
  nand (_28485_, _12555_, _12269_);
  and (_28486_, _28485_, _06373_);
  and (_28487_, _28486_, _28484_);
  or (_28488_, _28487_, _12245_);
  or (_28489_, _28488_, _28483_);
  or (_28491_, _28390_, _12246_);
  and (_28492_, _28491_, _07164_);
  and (_28493_, _28492_, _28489_);
  or (_28494_, _28493_, _28184_);
  and (_28495_, _28494_, _28397_);
  nand (_28496_, _12127_, _06461_);
  nand (_28497_, _28496_, _12242_);
  or (_28498_, _28497_, _28495_);
  or (_28499_, _28390_, _12242_);
  and (_28500_, _28499_, _14007_);
  and (_28502_, _28500_, _28498_);
  or (_28503_, _28502_, _25090_);
  and (_28504_, _28503_, _14006_);
  or (_28505_, _28405_, _06506_);
  nand (_28506_, _28505_, _12237_);
  or (_28507_, _28506_, _28504_);
  or (_28508_, _28390_, _12237_);
  and (_28509_, _28508_, _12588_);
  and (_28510_, _28509_, _28507_);
  nor (_28511_, _12588_, _28405_);
  or (_28512_, _28511_, _05976_);
  or (_28513_, _28512_, _28510_);
  or (_28514_, _28390_, _05977_);
  and (_28515_, _28514_, _06242_);
  and (_28516_, _28515_, _28513_);
  nand (_28517_, _12127_, _06241_);
  nand (_28518_, _28517_, _27873_);
  or (_28519_, _28518_, _28516_);
  nand (_28520_, _12269_, _06369_);
  and (_28521_, _28520_, _12603_);
  and (_28524_, _28521_, _28519_);
  nor (_28525_, _12603_, _28405_);
  or (_28526_, _28525_, _05968_);
  or (_28527_, _28526_, _28524_);
  nand (_28528_, _12269_, _05968_);
  and (_28529_, _28528_, _12611_);
  and (_28530_, _28529_, _28527_);
  and (_28531_, _28390_, _12615_);
  nor (_28532_, _28531_, _28530_);
  nor (_28533_, _28532_, _06332_);
  nand (_28535_, _12127_, _06332_);
  nand (_28536_, _28535_, _27742_);
  or (_28537_, _28536_, _28533_);
  or (_28538_, _28425_, _12620_);
  and (_28539_, _28538_, _08972_);
  and (_28540_, _28539_, _28537_);
  nor (_28541_, _28405_, _08972_);
  or (_28542_, _28541_, _06371_);
  or (_28543_, _28542_, _28540_);
  nand (_28544_, _12269_, _06371_);
  and (_28546_, _28544_, _10905_);
  and (_28547_, _28546_, _28543_);
  and (_28548_, _12127_, _10904_);
  or (_28549_, _28548_, _12634_);
  or (_28550_, _28549_, _28547_);
  nor (_28551_, _12662_, \oc8051_golden_model_1.DPH [2]);
  nor (_28552_, _28551_, _12663_);
  or (_28553_, _28552_, _12635_);
  and (_28554_, _28553_, _06921_);
  and (_28555_, _28554_, _28550_);
  and (_28557_, _12127_, _06331_);
  or (_28558_, _28557_, _28555_);
  nor (_28559_, _12677_, _05895_);
  and (_28560_, _28559_, _28558_);
  or (_28561_, _28425_, _11291_);
  or (_28562_, _12127_, _12684_);
  and (_28563_, _28562_, _12677_);
  and (_28564_, _28563_, _28561_);
  or (_28565_, _28564_, _12682_);
  or (_28566_, _28565_, _28560_);
  or (_28568_, _28390_, _12232_);
  and (_28569_, _28568_, _12228_);
  and (_28570_, _28569_, _28566_);
  nor (_28571_, _28405_, _12228_);
  or (_28572_, _28571_, _06367_);
  or (_28573_, _28572_, _28570_);
  nand (_28574_, _12269_, _06367_);
  and (_28575_, _28574_, _28573_);
  or (_28576_, _28575_, _06533_);
  nand (_28577_, _28405_, _06533_);
  nor (_28579_, _12701_, _05889_);
  and (_28580_, _28579_, _28577_);
  and (_28581_, _28580_, _28576_);
  or (_28582_, _28425_, _12684_);
  or (_28583_, _12127_, _11291_);
  and (_28584_, _28583_, _12701_);
  and (_28585_, _28584_, _28582_);
  or (_28586_, _28585_, _12710_);
  or (_28587_, _28586_, _28581_);
  or (_28588_, _28390_, _12226_);
  and (_28590_, _28588_, _10967_);
  and (_28591_, _28590_, _28587_);
  nor (_28592_, _28405_, _10967_);
  or (_28593_, _28592_, _06366_);
  or (_28594_, _28593_, _28591_);
  and (_28595_, _28594_, _28396_);
  or (_28596_, _28595_, _06541_);
  nand (_28597_, _28405_, _06541_);
  and (_28598_, _28597_, _27952_);
  and (_28599_, _28598_, _28596_);
  or (_28601_, _28425_, \oc8051_golden_model_1.PSW [7]);
  or (_28602_, _12127_, _10854_);
  and (_28603_, _28602_, _12723_);
  and (_28604_, _28603_, _28601_);
  or (_28605_, _28604_, _12738_);
  or (_28606_, _28605_, _28599_);
  or (_28607_, _28390_, _12736_);
  and (_28608_, _28607_, _11005_);
  and (_28609_, _28608_, _28606_);
  nor (_28610_, _28405_, _11005_);
  or (_28612_, _28610_, _06383_);
  or (_28613_, _28612_, _28609_);
  and (_28614_, _28613_, _28395_);
  or (_28615_, _28614_, _06528_);
  nand (_28616_, _28405_, _06528_);
  and (_28617_, _28616_, _27976_);
  and (_28618_, _28617_, _28615_);
  or (_28619_, _28425_, _10854_);
  or (_28620_, _12127_, \oc8051_golden_model_1.PSW [7]);
  and (_28621_, _28620_, _12215_);
  and (_28623_, _28621_, _28619_);
  or (_28624_, _28623_, _12758_);
  or (_28625_, _28624_, _28618_);
  or (_28626_, _28390_, _12756_);
  and (_28627_, _28626_, _11051_);
  and (_28628_, _28627_, _28625_);
  nor (_28629_, _28405_, _11051_);
  or (_28630_, _28629_, _11080_);
  or (_28631_, _28630_, _28628_);
  and (_28632_, _28631_, _28394_);
  or (_28634_, _28632_, _06547_);
  nand (_28635_, _07578_, _06547_);
  and (_28636_, _28635_, _28323_);
  and (_28637_, _28636_, _28634_);
  or (_28638_, _28399_, _12955_);
  or (_28639_, _12268_, _12954_);
  and (_28640_, _28639_, _06381_);
  and (_28641_, _28640_, _28638_);
  or (_28642_, _28641_, _12774_);
  or (_28643_, _28642_, _28637_);
  or (_28645_, _28390_, _12105_);
  and (_28646_, _28645_, _12963_);
  and (_28647_, _28646_, _28643_);
  nor (_28648_, _12963_, _28405_);
  or (_28649_, _28648_, _10448_);
  or (_28650_, _28649_, _28647_);
  and (_28651_, _28650_, _28393_);
  or (_28652_, _28651_, _06260_);
  nand (_28653_, _07578_, _06260_);
  and (_28654_, _28653_, _28344_);
  and (_28656_, _28654_, _28652_);
  or (_28657_, _28399_, _12954_);
  nand (_28658_, _12269_, _12954_);
  and (_28659_, _28658_, _28657_);
  and (_28660_, _28659_, _06377_);
  or (_28661_, _28660_, _12985_);
  or (_28662_, _28661_, _28656_);
  and (_28663_, _28662_, _28392_);
  or (_28664_, _28663_, _06563_);
  nand (_28665_, _28405_, _06563_);
  and (_28667_, _28665_, _12991_);
  and (_28668_, _28667_, _28664_);
  and (_28669_, _28390_, _12992_);
  or (_28670_, _28669_, _06378_);
  or (_28671_, _28670_, _28668_);
  nand (_28672_, _06750_, _06378_);
  and (_28673_, _28672_, _28038_);
  and (_28674_, _28673_, _28671_);
  and (_28675_, _28659_, _06199_);
  or (_28676_, _28675_, _13007_);
  or (_28678_, _28676_, _28674_);
  or (_28679_, _28390_, _13006_);
  and (_28680_, _28679_, _28678_);
  or (_28681_, _28680_, _06188_);
  nand (_28682_, _28405_, _06188_);
  and (_28683_, _28682_, _13013_);
  and (_28684_, _28683_, _28681_);
  and (_28685_, _28390_, _13014_);
  or (_28686_, _28685_, _06342_);
  or (_28687_, _28686_, _28684_);
  nand (_28689_, _06750_, _06342_);
  and (_28690_, _28689_, _28055_);
  and (_28691_, _28690_, _28687_);
  and (_28692_, _28390_, _13025_);
  or (_28693_, _28692_, _28691_);
  or (_28694_, _28693_, _01456_);
  or (_28695_, _01452_, \oc8051_golden_model_1.PC [10]);
  and (_28696_, _28695_, _43223_);
  and (_43865_, _28696_, _28694_);
  and (_28697_, _12092_, _09412_);
  nor (_28699_, _28697_, _12119_);
  and (_28700_, _28697_, _12119_);
  or (_28701_, _28700_, _28699_);
  nor (_28702_, _28701_, _12105_);
  and (_28703_, _12122_, \oc8051_golden_model_1.PSW [7]);
  nor (_28704_, _28422_, _12128_);
  and (_28705_, _28704_, _12125_);
  nor (_28706_, _28704_, _12125_);
  nor (_28707_, _28706_, _28705_);
  nor (_28708_, _28707_, \oc8051_golden_model_1.PSW [7]);
  or (_28710_, _28708_, _28703_);
  and (_28711_, _28710_, _12723_);
  nor (_28712_, _28701_, _12226_);
  nor (_28713_, _28701_, _12232_);
  nor (_28714_, _12122_, _08972_);
  and (_28715_, _12263_, _05968_);
  and (_28716_, _12392_, _12263_);
  or (_28717_, _12265_, _12266_);
  and (_28718_, _28717_, _12344_);
  nor (_28719_, _28717_, _12344_);
  nor (_28721_, _28719_, _28718_);
  not (_28722_, _28721_);
  nor (_28723_, _28722_, _12392_);
  or (_28724_, _28723_, _28716_);
  nor (_28725_, _28724_, _06345_);
  and (_28726_, _12513_, _12263_);
  nor (_28727_, _28722_, _12513_);
  or (_28728_, _28727_, _28726_);
  nor (_28729_, _28728_, _12478_);
  and (_28730_, _12122_, _06466_);
  and (_28732_, _12419_, _12119_);
  nor (_28733_, _28732_, _07123_);
  and (_28734_, _12122_, _07123_);
  or (_28735_, _28734_, _06808_);
  or (_28736_, _28735_, _28733_);
  or (_28737_, _28701_, _12420_);
  and (_28738_, _28737_, _25018_);
  and (_28739_, _28738_, _28736_);
  and (_28740_, _12122_, _06705_);
  not (_28741_, _28701_);
  nor (_28743_, _28741_, _12427_);
  or (_28744_, _28743_, _08572_);
  or (_28745_, _28744_, _28740_);
  nor (_28746_, _28745_, _28739_);
  and (_28747_, _12412_, _12122_);
  not (_28748_, _28747_);
  nor (_28749_, _28707_, _12412_);
  nor (_28750_, _28749_, _08573_);
  and (_28751_, _28750_, _28748_);
  nor (_28752_, _28751_, _28746_);
  nor (_28754_, _28752_, _07134_);
  and (_28755_, _28741_, _07134_);
  nor (_28756_, _28755_, _28754_);
  and (_28757_, _28756_, _06252_);
  and (_28758_, _12402_, _12263_);
  and (_28759_, _28721_, _12404_);
  or (_28760_, _28759_, _28758_);
  and (_28761_, _28760_, _06251_);
  or (_28762_, _28761_, _12444_);
  nor (_28763_, _28762_, _28757_);
  nor (_28765_, _28701_, _12443_);
  or (_28766_, _28765_, _28763_);
  nor (_28767_, _28766_, _12453_);
  not (_28768_, _12122_);
  nor (_28769_, _12447_, _28768_);
  nor (_28770_, _28769_, _12452_);
  not (_28771_, _28770_);
  nor (_28772_, _28771_, _28767_);
  nor (_28773_, _28701_, _12451_);
  nor (_28774_, _28773_, _06466_);
  not (_28776_, _28774_);
  nor (_28777_, _28776_, _28772_);
  nor (_28778_, _28777_, _28730_);
  nor (_28779_, _28778_, _12464_);
  nor (_28780_, _28741_, _12462_);
  nor (_28781_, _28780_, _12469_);
  not (_28782_, _28781_);
  nor (_28783_, _28782_, _28779_);
  nor (_28784_, _12468_, _12122_);
  nor (_28785_, _28784_, _28783_);
  nor (_28787_, _28785_, _12479_);
  nor (_28788_, _28787_, _28729_);
  nor (_28789_, _28788_, _06344_);
  nor (_28790_, _28789_, _28725_);
  nand (_28791_, _28790_, _12536_);
  and (_28792_, _12533_, _12263_);
  nor (_28793_, _28722_, _12533_);
  nor (_28794_, _28793_, _28792_);
  or (_28795_, _28794_, _12536_);
  and (_28796_, _28795_, _28791_);
  or (_28798_, _28796_, _06373_);
  nand (_28799_, _12555_, _12263_);
  not (_28800_, _12555_);
  nand (_28801_, _28721_, _28800_);
  and (_28802_, _28801_, _28799_);
  or (_28803_, _28802_, _12522_);
  nand (_28804_, _28803_, _28798_);
  nand (_28805_, _28804_, _12246_);
  not (_28806_, _12573_);
  and (_28807_, _28701_, _12245_);
  nor (_28809_, _28807_, _28806_);
  nand (_28810_, _28809_, _28805_);
  nor (_28811_, _12573_, _12122_);
  nor (_28812_, _28811_, _12243_);
  nand (_28813_, _28812_, _28810_);
  nor (_28814_, _28741_, _12242_);
  nor (_28815_, _28814_, _12583_);
  and (_28816_, _28815_, _28813_);
  nor (_28817_, _12580_, _12122_);
  or (_28818_, _28817_, _12582_);
  or (_28820_, _28818_, _28816_);
  nor (_28821_, _28741_, _12237_);
  nor (_28822_, _28821_, _12589_);
  nand (_28823_, _28822_, _28820_);
  nor (_28824_, _12588_, _12122_);
  nor (_28825_, _28824_, _05976_);
  nand (_28826_, _28825_, _28823_);
  and (_28827_, _28701_, _05976_);
  nor (_28828_, _28827_, _12596_);
  nand (_28829_, _28828_, _28826_);
  nor (_28831_, _12595_, _12122_);
  nor (_28832_, _28831_, _06369_);
  nand (_28833_, _28832_, _28829_);
  and (_28834_, _12263_, _06369_);
  nor (_28835_, _28834_, _12604_);
  nand (_28836_, _28835_, _28833_);
  nor (_28837_, _12603_, _12122_);
  nor (_28838_, _28837_, _05968_);
  and (_28839_, _28838_, _28836_);
  or (_28840_, _28839_, _28715_);
  nand (_28842_, _28840_, _12611_);
  nor (_28843_, _28741_, _12611_);
  nor (_28844_, _28843_, _12614_);
  nand (_28845_, _28844_, _28842_);
  nor (_28846_, _12613_, _12122_);
  nor (_28847_, _28846_, _12619_);
  nand (_28848_, _28847_, _28845_);
  nor (_28849_, _28707_, _12620_);
  nor (_28850_, _28849_, _08973_);
  and (_28851_, _28850_, _28848_);
  or (_28853_, _28851_, _28714_);
  nand (_28854_, _28853_, _07198_);
  and (_28855_, _12264_, _06371_);
  nor (_28856_, _28855_, _10904_);
  and (_28857_, _28856_, _28854_);
  and (_28858_, _12122_, _10904_);
  or (_28859_, _28858_, _28857_);
  nand (_28860_, _28859_, _12635_);
  nor (_28861_, _12663_, \oc8051_golden_model_1.DPH [3]);
  not (_28862_, _28861_);
  nor (_28864_, _12665_, _12635_);
  and (_28865_, _28864_, _28862_);
  nor (_28866_, _28865_, _12674_);
  nand (_28867_, _28866_, _28860_);
  nor (_28868_, _12673_, _12122_);
  nor (_28869_, _28868_, _12677_);
  nand (_28870_, _28869_, _28867_);
  and (_28871_, _12122_, _11291_);
  nor (_28872_, _28707_, _11291_);
  or (_28873_, _28872_, _28871_);
  and (_28875_, _28873_, _12677_);
  nor (_28876_, _28875_, _12682_);
  and (_28877_, _28876_, _28870_);
  or (_28878_, _28877_, _28713_);
  nand (_28879_, _28878_, _12228_);
  nor (_28880_, _12122_, _12228_);
  nor (_28881_, _28880_, _06367_);
  nand (_28882_, _28881_, _28879_);
  and (_28883_, _12263_, _06367_);
  nor (_28884_, _28883_, _12698_);
  nand (_28885_, _28884_, _28882_);
  nor (_28886_, _12697_, _12122_);
  nor (_28887_, _28886_, _12701_);
  nand (_28888_, _28887_, _28885_);
  and (_28889_, _12122_, _12684_);
  nor (_28890_, _28707_, _12684_);
  or (_28891_, _28890_, _28889_);
  and (_28892_, _28891_, _12701_);
  nor (_28893_, _28892_, _12710_);
  and (_28894_, _28893_, _28888_);
  or (_28897_, _28894_, _28712_);
  nand (_28898_, _28897_, _10967_);
  nor (_28899_, _12122_, _10967_);
  nor (_28900_, _28899_, _06366_);
  nand (_28901_, _28900_, _28898_);
  and (_28902_, _12263_, _06366_);
  nor (_28903_, _28902_, _12720_);
  nand (_28904_, _28903_, _28901_);
  nor (_28905_, _12719_, _12122_);
  nor (_28906_, _28905_, _12723_);
  and (_28908_, _28906_, _28904_);
  or (_28909_, _28908_, _28711_);
  nand (_28910_, _28909_, _12736_);
  nor (_28911_, _28741_, _12736_);
  nor (_28912_, _28911_, _11006_);
  nand (_28913_, _28912_, _28910_);
  nor (_28914_, _12122_, _11005_);
  nor (_28915_, _28914_, _06383_);
  nand (_28916_, _28915_, _28913_);
  and (_28917_, _12263_, _06383_);
  nor (_28919_, _28917_, _12748_);
  nand (_28920_, _28919_, _28916_);
  nor (_28921_, _12747_, _12122_);
  nor (_28922_, _28921_, _12215_);
  nand (_28923_, _28922_, _28920_);
  nand (_28924_, _12122_, _10854_);
  or (_28925_, _28707_, _10854_);
  and (_28926_, _28925_, _28924_);
  or (_28927_, _28926_, _12751_);
  nand (_28928_, _28927_, _28923_);
  nand (_28930_, _28928_, _12756_);
  nor (_28931_, _28741_, _12756_);
  nor (_28932_, _28931_, _11052_);
  nand (_28933_, _28932_, _28930_);
  nor (_28934_, _12122_, _11051_);
  nor (_28935_, _28934_, _11080_);
  and (_28936_, _28935_, _28933_);
  and (_28937_, _28701_, _11080_);
  or (_28938_, _28937_, _06547_);
  nor (_28939_, _28938_, _28936_);
  and (_28941_, _07713_, _06547_);
  or (_28942_, _28941_, _28939_);
  nand (_28943_, _28942_, _05916_);
  nor (_28944_, _12122_, _05916_);
  nor (_28945_, _28944_, _06381_);
  nand (_28946_, _28945_, _28943_);
  nor (_28947_, _12263_, _12954_);
  and (_28948_, _28722_, _12954_);
  or (_28949_, _28948_, _06946_);
  or (_28950_, _28949_, _28947_);
  and (_28952_, _28950_, _12105_);
  and (_28953_, _28952_, _28946_);
  or (_28954_, _28953_, _28702_);
  nand (_28955_, _28954_, _12963_);
  nor (_28956_, _12963_, _12122_);
  nor (_28957_, _28956_, _10448_);
  nand (_28958_, _28957_, _28955_);
  and (_28959_, _28701_, _10448_);
  nor (_28960_, _28959_, _06260_);
  and (_28961_, _28960_, _28958_);
  and (_28963_, _07713_, _06260_);
  or (_28964_, _28963_, _28961_);
  nand (_28965_, _28964_, _05924_);
  nor (_28966_, _12122_, _05924_);
  nor (_28967_, _28966_, _06377_);
  nand (_28968_, _28967_, _28965_);
  nor (_28969_, _28721_, _12954_);
  and (_28970_, _12264_, _12954_);
  nor (_28971_, _28970_, _28969_);
  and (_28972_, _28971_, _06377_);
  nor (_28974_, _28972_, _12985_);
  nand (_28975_, _28974_, _28968_);
  nor (_28976_, _28701_, _12984_);
  nor (_28977_, _28976_, _06563_);
  nand (_28978_, _28977_, _28975_);
  and (_28979_, _12122_, _06563_);
  nor (_28980_, _28979_, _12992_);
  nand (_28981_, _28980_, _28978_);
  nor (_28982_, _28701_, _12991_);
  nor (_28983_, _28982_, _06378_);
  nand (_28985_, _28983_, _28981_);
  nor (_28986_, _08505_, _06292_);
  nor (_28987_, _28986_, _05912_);
  nand (_28988_, _28987_, _28985_);
  and (_28989_, _28768_, _05912_);
  nor (_28990_, _28989_, _06199_);
  nand (_28991_, _28990_, _28988_);
  and (_28992_, _28971_, _06199_);
  nor (_28993_, _28992_, _13007_);
  nand (_28994_, _28993_, _28991_);
  nor (_28996_, _28701_, _13006_);
  nor (_28997_, _28996_, _06188_);
  nand (_28998_, _28997_, _28994_);
  and (_28999_, _12122_, _06188_);
  nor (_29000_, _28999_, _13014_);
  nand (_29001_, _29000_, _28998_);
  nor (_29002_, _28701_, _13013_);
  nor (_29003_, _29002_, _06342_);
  nand (_29004_, _29003_, _29001_);
  nor (_29005_, _13018_, _06292_);
  nor (_29007_, _29005_, _05907_);
  and (_29008_, _29007_, _29004_);
  and (_29009_, _28768_, _05907_);
  nor (_29010_, _29009_, _29008_);
  and (_29011_, _29010_, _13026_);
  and (_29012_, _28701_, _13025_);
  or (_29013_, _29012_, _29011_);
  or (_29014_, _29013_, _01456_);
  or (_29015_, _01452_, \oc8051_golden_model_1.PC [11]);
  and (_29016_, _29015_, _43223_);
  and (_43866_, _29016_, _29014_);
  and (_29018_, _06230_, _06342_);
  or (_29019_, _29018_, _05907_);
  and (_29020_, _28697_, \oc8051_golden_model_1.PC [11]);
  and (_29021_, _29020_, \oc8051_golden_model_1.PC [12]);
  nor (_29022_, _29020_, \oc8051_golden_model_1.PC [12]);
  nor (_29023_, _29022_, _29021_);
  not (_29024_, _29023_);
  and (_29025_, _29024_, _10448_);
  not (_29026_, _12117_);
  nor (_29028_, _12747_, _29026_);
  nor (_29029_, _12719_, _29026_);
  nor (_29030_, _12697_, _29026_);
  nor (_29031_, _29023_, _12237_);
  and (_29032_, _12392_, _12259_);
  nor (_29033_, _12348_, _12346_);
  nor (_29034_, _29033_, _12349_);
  nor (_29035_, _29034_, _12392_);
  or (_29036_, _29035_, _06345_);
  nor (_29037_, _29036_, _29032_);
  nor (_29039_, _12468_, _29026_);
  nor (_29040_, _29023_, _12451_);
  and (_29041_, _29023_, _07134_);
  and (_29042_, _12412_, _12117_);
  and (_29043_, _12200_, _12197_);
  nor (_29044_, _29043_, _12201_);
  and (_29045_, _29044_, _12414_);
  or (_29046_, _29045_, _29042_);
  nor (_29047_, _29046_, _08573_);
  nor (_29048_, _29024_, _28415_);
  not (_29050_, _29048_);
  and (_29051_, _12117_, _07123_);
  and (_29052_, _07124_, \oc8051_golden_model_1.PC [12]);
  and (_29053_, _29052_, _12419_);
  nor (_29054_, _29053_, _29051_);
  not (_29055_, _29054_);
  and (_29056_, _25018_, _12418_);
  and (_29057_, _29056_, _29055_);
  and (_29058_, _12117_, _06705_);
  nor (_29059_, _29058_, _08572_);
  not (_29061_, _29059_);
  nor (_29062_, _29061_, _29057_);
  and (_29063_, _29062_, _29050_);
  or (_29064_, _29063_, _07134_);
  nor (_29065_, _29064_, _29047_);
  or (_29066_, _29065_, _29041_);
  nor (_29067_, _29066_, _06251_);
  not (_29068_, _29034_);
  and (_29069_, _29068_, _12404_);
  nor (_29070_, _12404_, _12258_);
  nor (_29072_, _29070_, _29069_);
  nor (_29073_, _29072_, _06252_);
  nor (_29074_, _29073_, _29067_);
  nor (_29075_, _29074_, _12444_);
  nor (_29076_, _29023_, _12443_);
  nor (_29077_, _29076_, _12453_);
  not (_29078_, _29077_);
  nor (_29079_, _29078_, _29075_);
  nor (_29080_, _12447_, _29026_);
  or (_29081_, _29080_, _12452_);
  nor (_29083_, _29081_, _29079_);
  nor (_29084_, _29083_, _29040_);
  nor (_29085_, _29084_, _06466_);
  and (_29086_, _29026_, _06466_);
  nor (_29087_, _29086_, _12464_);
  not (_29088_, _29087_);
  nor (_29089_, _29088_, _29085_);
  nor (_29090_, _29024_, _12462_);
  nor (_29091_, _29090_, _29089_);
  nor (_29092_, _29091_, _12469_);
  or (_29094_, _29092_, _12479_);
  nor (_29095_, _29094_, _29039_);
  and (_29096_, _12513_, _12258_);
  nor (_29097_, _29068_, _12513_);
  or (_29098_, _29097_, _12478_);
  nor (_29099_, _29098_, _29096_);
  or (_29100_, _29099_, _06344_);
  nor (_29101_, _29100_, _29095_);
  or (_29102_, _29101_, _29037_);
  or (_29103_, _29102_, _06338_);
  nor (_29105_, _29068_, _12533_);
  and (_29106_, _12533_, _12258_);
  or (_29107_, _29106_, _12536_);
  or (_29108_, _29107_, _29105_);
  and (_29109_, _29108_, _12522_);
  and (_29110_, _29109_, _29103_);
  and (_29111_, _12555_, _12258_);
  and (_29112_, _29034_, _28800_);
  or (_29113_, _29112_, _29111_);
  and (_29114_, _29113_, _06373_);
  or (_29116_, _29114_, _29110_);
  and (_29117_, _29116_, _12246_);
  and (_29118_, _29023_, _12245_);
  or (_29119_, _29118_, _29117_);
  nor (_29120_, _29119_, _28806_);
  nor (_29121_, _12573_, _12117_);
  nor (_29122_, _29121_, _29120_);
  nor (_29123_, _29122_, _12243_);
  nor (_29124_, _29023_, _12242_);
  nor (_29125_, _29124_, _12583_);
  not (_29127_, _29125_);
  nor (_29128_, _29127_, _29123_);
  nor (_29129_, _12580_, _29026_);
  nor (_29130_, _29129_, _12582_);
  not (_29131_, _29130_);
  nor (_29132_, _29131_, _29128_);
  or (_29133_, _29132_, _12589_);
  nor (_29134_, _29133_, _29031_);
  nor (_29135_, _12588_, _29026_);
  nor (_29136_, _29135_, _05976_);
  not (_29138_, _29136_);
  or (_29139_, _29138_, _29134_);
  and (_29140_, _29024_, _05976_);
  nor (_29141_, _29140_, _12596_);
  nand (_29142_, _29141_, _29139_);
  nor (_29143_, _12595_, _29026_);
  nor (_29144_, _29143_, _06369_);
  nand (_29145_, _29144_, _29142_);
  and (_29146_, _12259_, _06369_);
  nor (_29147_, _29146_, _12604_);
  nand (_29149_, _29147_, _29145_);
  nor (_29150_, _12603_, _29026_);
  nor (_29151_, _29150_, _05968_);
  nand (_29152_, _29151_, _29149_);
  and (_29153_, _12259_, _05968_);
  nor (_29154_, _29153_, _12615_);
  nand (_29155_, _29154_, _29152_);
  nor (_29156_, _29024_, _12611_);
  nor (_29157_, _29156_, _12614_);
  nand (_29158_, _29157_, _29155_);
  nor (_29160_, _12613_, _12117_);
  nor (_29161_, _29160_, _12619_);
  nand (_29162_, _29161_, _29158_);
  and (_29163_, _29044_, _12619_);
  nor (_29164_, _29163_, _08973_);
  and (_29165_, _29164_, _29162_);
  nor (_29166_, _12117_, _08972_);
  or (_29167_, _29166_, _29165_);
  nand (_29168_, _29167_, _07198_);
  and (_29169_, _12259_, _06371_);
  nor (_29171_, _29169_, _10904_);
  nand (_29172_, _29171_, _29168_);
  and (_29173_, _12117_, _10904_);
  nor (_29174_, _29173_, _12634_);
  nand (_29175_, _29174_, _29172_);
  nor (_29176_, _12665_, \oc8051_golden_model_1.DPH [4]);
  nor (_29177_, _29176_, _12666_);
  nor (_29178_, _29177_, _12635_);
  nor (_29179_, _29178_, _12674_);
  and (_29180_, _29179_, _29175_);
  nor (_29182_, _12673_, _29026_);
  or (_29183_, _29182_, _29180_);
  nand (_29184_, _29183_, _12678_);
  nor (_29185_, _29044_, _11291_);
  nor (_29186_, _12117_, _12684_);
  nor (_29187_, _29186_, _12678_);
  not (_29188_, _29187_);
  nor (_29189_, _29188_, _29185_);
  nor (_29190_, _29189_, _12682_);
  nand (_29191_, _29190_, _29184_);
  nor (_29193_, _29023_, _12232_);
  nor (_29194_, _29193_, _12229_);
  nand (_29195_, _29194_, _29191_);
  nor (_29196_, _29026_, _12228_);
  nor (_29197_, _29196_, _06367_);
  nand (_29198_, _29197_, _29195_);
  and (_29199_, _12259_, _06367_);
  nor (_29200_, _29199_, _12698_);
  and (_29201_, _29200_, _29198_);
  or (_29202_, _29201_, _29030_);
  nand (_29204_, _29202_, _12702_);
  and (_29205_, _12117_, _12684_);
  and (_29206_, _29044_, _11291_);
  or (_29207_, _29206_, _29205_);
  and (_29208_, _29207_, _12701_);
  nor (_29209_, _29208_, _12710_);
  nand (_29210_, _29209_, _29204_);
  nor (_29211_, _29023_, _12226_);
  nor (_29212_, _29211_, _10968_);
  nand (_29213_, _29212_, _29210_);
  nor (_29215_, _29026_, _10967_);
  nor (_29216_, _29215_, _06366_);
  nand (_29217_, _29216_, _29213_);
  and (_29218_, _12259_, _06366_);
  nor (_29219_, _29218_, _12720_);
  and (_29220_, _29219_, _29217_);
  or (_29221_, _29220_, _29029_);
  nand (_29222_, _29221_, _12724_);
  and (_29223_, _12117_, \oc8051_golden_model_1.PSW [7]);
  and (_29224_, _29044_, _10854_);
  or (_29226_, _29224_, _29223_);
  and (_29227_, _29226_, _12723_);
  nor (_29228_, _29227_, _12738_);
  nand (_29229_, _29228_, _29222_);
  nor (_29230_, _29023_, _12736_);
  nor (_29231_, _29230_, _11006_);
  nand (_29232_, _29231_, _29229_);
  nor (_29233_, _29026_, _11005_);
  nor (_29234_, _29233_, _06383_);
  nand (_29235_, _29234_, _29232_);
  and (_29237_, _12259_, _06383_);
  nor (_29238_, _29237_, _12748_);
  and (_29239_, _29238_, _29235_);
  or (_29240_, _29239_, _29028_);
  nand (_29241_, _29240_, _12751_);
  and (_29242_, _12117_, _10854_);
  and (_29243_, _29044_, \oc8051_golden_model_1.PSW [7]);
  or (_29244_, _29243_, _29242_);
  and (_29245_, _29244_, _12215_);
  nor (_29246_, _29245_, _12758_);
  nand (_29248_, _29246_, _29241_);
  nor (_29249_, _29023_, _12756_);
  nor (_29250_, _29249_, _11052_);
  nand (_29251_, _29250_, _29248_);
  nor (_29252_, _29026_, _11051_);
  nor (_29253_, _29252_, _11080_);
  nand (_29254_, _29253_, _29251_);
  and (_29255_, _29024_, _11080_);
  nor (_29256_, _29255_, _06547_);
  and (_29257_, _29256_, _29254_);
  nor (_29259_, _08494_, _13873_);
  or (_29260_, _29259_, _07228_);
  or (_29261_, _29260_, _29257_);
  nor (_29262_, _12117_, _05916_);
  nor (_29263_, _29262_, _06381_);
  nand (_29264_, _29263_, _29261_);
  nor (_29265_, _12258_, _12954_);
  and (_29266_, _29068_, _12954_);
  or (_29267_, _29266_, _06946_);
  or (_29268_, _29267_, _29265_);
  and (_29270_, _29268_, _12105_);
  nand (_29271_, _29270_, _29264_);
  nor (_29272_, _29023_, _12105_);
  nor (_29273_, _29272_, _12964_);
  nand (_29274_, _29273_, _29271_);
  nor (_29275_, _12963_, _29026_);
  nor (_29276_, _29275_, _10448_);
  and (_29277_, _29276_, _29274_);
  or (_29278_, _29277_, _29025_);
  nand (_29279_, _29278_, _06261_);
  and (_29281_, _08494_, _06260_);
  nor (_29282_, _29281_, _12089_);
  and (_29283_, _29282_, _29279_);
  nor (_29284_, _29026_, _05924_);
  or (_29285_, _29284_, _06377_);
  nor (_29286_, _29285_, _29283_);
  nor (_29287_, _29034_, _12954_);
  and (_29288_, _12259_, _12954_);
  nor (_29289_, _29288_, _29287_);
  nor (_29290_, _29289_, _06564_);
  or (_29292_, _29290_, _29286_);
  and (_29293_, _29292_, _12984_);
  nor (_29294_, _29023_, _12984_);
  or (_29295_, _29294_, _29293_);
  nand (_29296_, _29295_, _07241_);
  nand (_29297_, _29026_, _06563_);
  and (_29298_, _29297_, _12991_);
  nand (_29299_, _29298_, _29296_);
  nor (_29300_, _29024_, _12991_);
  nor (_29301_, _29300_, _06378_);
  nand (_29303_, _29301_, _29299_);
  and (_29304_, _06230_, _06378_);
  nor (_29305_, _29304_, _05912_);
  and (_29306_, _29305_, _29303_);
  and (_29307_, _12117_, _05912_);
  or (_29308_, _29307_, _06199_);
  or (_29309_, _29308_, _29306_);
  nor (_29310_, _29289_, _06571_);
  nor (_29311_, _29310_, _13007_);
  nand (_29312_, _29311_, _29309_);
  nor (_29314_, _29024_, _13006_);
  nor (_29315_, _29314_, _06188_);
  nand (_29316_, _29315_, _29312_);
  and (_29317_, _29026_, _06188_);
  nor (_29318_, _29317_, _13014_);
  nand (_29319_, _29318_, _29316_);
  nor (_29320_, _29024_, _13013_);
  nor (_29321_, _29320_, _06342_);
  and (_29322_, _29321_, _29319_);
  or (_29323_, _29322_, _29019_);
  and (_29325_, _12117_, _05907_);
  nor (_29326_, _29325_, _13025_);
  and (_29327_, _29326_, _29323_);
  and (_29328_, _29024_, _13025_);
  nor (_29329_, _29328_, _29327_);
  or (_29330_, _29329_, _01456_);
  or (_29331_, _01452_, \oc8051_golden_model_1.PC [12]);
  and (_29332_, _29331_, _43223_);
  and (_43867_, _29332_, _29330_);
  and (_29333_, _29021_, \oc8051_golden_model_1.PC [13]);
  nor (_29335_, _29021_, \oc8051_golden_model_1.PC [13]);
  nor (_29336_, _29335_, _29333_);
  or (_29337_, _29336_, _12105_);
  or (_29338_, _12115_, _12114_);
  not (_29339_, _29338_);
  nor (_29340_, _29339_, _12202_);
  and (_29341_, _29339_, _12202_);
  or (_29342_, _29341_, _29340_);
  or (_29343_, _29342_, _10854_);
  or (_29344_, _12113_, \oc8051_golden_model_1.PSW [7]);
  and (_29346_, _29344_, _12215_);
  and (_29347_, _29346_, _29343_);
  or (_29348_, _29336_, _12226_);
  or (_29349_, _29336_, _12232_);
  and (_29350_, _12253_, _05968_);
  or (_29351_, _12254_, _12255_);
  not (_29352_, _29351_);
  nor (_29353_, _29352_, _12350_);
  and (_29354_, _29352_, _12350_);
  nor (_29355_, _29354_, _29353_);
  not (_29357_, _29355_);
  or (_29358_, _29357_, _12392_);
  or (_29359_, _27122_, _12253_);
  and (_29360_, _29359_, _06344_);
  and (_29361_, _29360_, _29358_);
  and (_29362_, _12113_, _06466_);
  or (_29363_, _12404_, _12253_);
  or (_29364_, _29357_, _12402_);
  and (_29365_, _29364_, _29363_);
  or (_29366_, _29365_, _06252_);
  and (_29368_, _12412_, _12113_);
  and (_29369_, _29342_, _12414_);
  or (_29370_, _29369_, _29368_);
  or (_29371_, _29370_, _08573_);
  or (_29372_, _29336_, _28415_);
  or (_29373_, _12428_, _12113_);
  nor (_29374_, _07123_, \oc8051_golden_model_1.PC [13]);
  and (_29375_, _29374_, _12420_);
  nand (_29376_, _29375_, _25018_);
  and (_29377_, _29376_, _29373_);
  and (_29379_, _29377_, _29372_);
  or (_29380_, _29379_, _08572_);
  and (_29381_, _29380_, _07338_);
  and (_29382_, _29381_, _29371_);
  and (_29383_, _29336_, _07134_);
  or (_29384_, _29383_, _06251_);
  or (_29385_, _29384_, _29382_);
  and (_29386_, _29385_, _29366_);
  or (_29387_, _29386_, _12444_);
  or (_29388_, _29336_, _12443_);
  and (_29390_, _29388_, _12447_);
  and (_29391_, _29390_, _29387_);
  nor (_29392_, _12447_, _15483_);
  or (_29393_, _29392_, _12452_);
  or (_29394_, _29393_, _29391_);
  or (_29395_, _29336_, _12451_);
  and (_29396_, _29395_, _06801_);
  and (_29397_, _29396_, _29394_);
  or (_29398_, _29397_, _29362_);
  and (_29399_, _29398_, _12462_);
  not (_29401_, _29336_);
  or (_29402_, _29401_, _12462_);
  nand (_29403_, _29402_, _12468_);
  or (_29404_, _29403_, _29399_);
  or (_29405_, _12468_, _12113_);
  and (_29406_, _29405_, _29404_);
  or (_29407_, _29406_, _12479_);
  and (_29408_, _12513_, _12253_);
  nor (_29409_, _29355_, _12513_);
  or (_29410_, _29409_, _29408_);
  or (_29411_, _29410_, _12478_);
  and (_29412_, _29411_, _06345_);
  and (_29413_, _29412_, _29407_);
  or (_29414_, _29413_, _06338_);
  or (_29415_, _29414_, _29361_);
  nor (_29416_, _29355_, _12533_);
  and (_29417_, _12533_, _12253_);
  or (_29418_, _29417_, _12536_);
  or (_29419_, _29418_, _29416_);
  and (_29420_, _29419_, _12522_);
  and (_29423_, _29420_, _29415_);
  nand (_29424_, _29355_, _28800_);
  or (_29425_, _28800_, _12253_);
  and (_29426_, _29425_, _06373_);
  and (_29427_, _29426_, _29424_);
  or (_29428_, _29427_, _29423_);
  and (_29429_, _29428_, _12246_);
  nand (_29430_, _29336_, _12245_);
  nand (_29431_, _29430_, _12573_);
  or (_29432_, _29431_, _29429_);
  or (_29434_, _12573_, _12113_);
  and (_29435_, _29434_, _12242_);
  and (_29436_, _29435_, _29432_);
  nor (_29437_, _29401_, _12242_);
  or (_29438_, _29437_, _12583_);
  or (_29439_, _29438_, _29436_);
  or (_29440_, _12580_, _12113_);
  and (_29441_, _29440_, _12237_);
  and (_29442_, _29441_, _29439_);
  nor (_29443_, _29401_, _12237_);
  or (_29445_, _29443_, _12589_);
  or (_29446_, _29445_, _29442_);
  or (_29447_, _12588_, _12113_);
  and (_29448_, _29447_, _05977_);
  and (_29449_, _29448_, _29446_);
  nand (_29450_, _29336_, _05976_);
  nand (_29451_, _29450_, _12595_);
  or (_29452_, _29451_, _29449_);
  or (_29453_, _12595_, _12113_);
  and (_29454_, _29453_, _06370_);
  and (_29456_, _29454_, _29452_);
  nand (_29457_, _12253_, _06369_);
  nand (_29458_, _29457_, _12603_);
  or (_29459_, _29458_, _29456_);
  or (_29460_, _12603_, _12113_);
  and (_29461_, _29460_, _06336_);
  and (_29462_, _29461_, _29459_);
  or (_29463_, _29462_, _29350_);
  and (_29464_, _29463_, _12611_);
  nor (_29465_, _29401_, _12611_);
  or (_29467_, _29465_, _12614_);
  or (_29468_, _29467_, _29464_);
  or (_29469_, _12613_, _12113_);
  and (_29470_, _29469_, _12620_);
  and (_29471_, _29470_, _29468_);
  and (_29472_, _29342_, _12619_);
  or (_29473_, _29472_, _08973_);
  or (_29474_, _29473_, _29471_);
  or (_29475_, _12113_, _08972_);
  and (_29476_, _29475_, _07198_);
  and (_29478_, _29476_, _29474_);
  and (_29479_, _12253_, _06371_);
  or (_29480_, _29479_, _10904_);
  or (_29481_, _29480_, _29478_);
  nand (_29482_, _15483_, _10904_);
  and (_29483_, _29482_, _12635_);
  and (_29484_, _29483_, _29481_);
  nor (_29485_, _12666_, \oc8051_golden_model_1.DPH [5]);
  nor (_29486_, _29485_, _12667_);
  and (_29487_, _29486_, _12634_);
  or (_29489_, _29487_, _12674_);
  or (_29490_, _29489_, _29484_);
  or (_29491_, _12673_, _12113_);
  and (_29492_, _29491_, _12678_);
  and (_29493_, _29492_, _29490_);
  or (_29494_, _29342_, _11291_);
  or (_29495_, _12113_, _12684_);
  and (_29496_, _29495_, _12677_);
  and (_29497_, _29496_, _29494_);
  or (_29498_, _29497_, _12682_);
  or (_29500_, _29498_, _29493_);
  and (_29501_, _29500_, _29349_);
  or (_29502_, _29501_, _12229_);
  or (_29503_, _12113_, _12228_);
  and (_29504_, _29503_, _07218_);
  and (_29505_, _29504_, _29502_);
  nand (_29506_, _12253_, _06367_);
  nand (_29507_, _29506_, _12697_);
  or (_29508_, _29507_, _29505_);
  or (_29509_, _12697_, _12113_);
  and (_29511_, _29509_, _12702_);
  and (_29512_, _29511_, _29508_);
  or (_29513_, _29342_, _12684_);
  or (_29514_, _12113_, _11291_);
  and (_29515_, _29514_, _12701_);
  and (_29516_, _29515_, _29513_);
  or (_29517_, _29516_, _12710_);
  or (_29518_, _29517_, _29512_);
  and (_29519_, _29518_, _29348_);
  or (_29520_, _29519_, _10968_);
  or (_29522_, _12113_, _10967_);
  and (_29523_, _29522_, _07213_);
  and (_29524_, _29523_, _29520_);
  nand (_29525_, _12253_, _06366_);
  nand (_29526_, _29525_, _12719_);
  or (_29527_, _29526_, _29524_);
  or (_29528_, _12719_, _12113_);
  and (_29529_, _29528_, _12724_);
  and (_29530_, _29529_, _29527_);
  or (_29531_, _29342_, \oc8051_golden_model_1.PSW [7]);
  or (_29533_, _12113_, _10854_);
  and (_29534_, _29533_, _12723_);
  and (_29535_, _29534_, _29531_);
  or (_29536_, _29535_, _29530_);
  and (_29537_, _29536_, _12736_);
  nor (_29538_, _29401_, _12736_);
  or (_29539_, _29538_, _11006_);
  or (_29540_, _29539_, _29537_);
  or (_29541_, _12113_, _11005_);
  and (_29542_, _29541_, _07231_);
  and (_29544_, _29542_, _29540_);
  nand (_29545_, _12253_, _06383_);
  nand (_29546_, _29545_, _12747_);
  or (_29547_, _29546_, _29544_);
  or (_29548_, _12747_, _12113_);
  and (_29549_, _29548_, _12751_);
  and (_29550_, _29549_, _29547_);
  or (_29551_, _29550_, _29347_);
  and (_29552_, _29551_, _12756_);
  nor (_29553_, _29401_, _12756_);
  or (_29555_, _29553_, _11052_);
  or (_29556_, _29555_, _29552_);
  or (_29557_, _12113_, _11051_);
  and (_29558_, _29557_, _11081_);
  and (_29559_, _29558_, _29556_);
  and (_29560_, _29336_, _11080_);
  or (_29561_, _29560_, _06547_);
  or (_29562_, _29561_, _29559_);
  nand (_29563_, _08209_, _06547_);
  and (_29564_, _29563_, _29562_);
  or (_29566_, _29564_, _07228_);
  nor (_29567_, _12113_, _05916_);
  nor (_29568_, _29567_, _06381_);
  and (_29569_, _29568_, _29566_);
  or (_29570_, _12253_, _12954_);
  nand (_29571_, _29355_, _12954_);
  and (_29572_, _29571_, _06381_);
  and (_29573_, _29572_, _29570_);
  or (_29574_, _29573_, _12774_);
  or (_29575_, _29574_, _29569_);
  and (_29577_, _29575_, _29337_);
  or (_29578_, _29577_, _12964_);
  or (_29579_, _12963_, _12113_);
  and (_29580_, _29579_, _12966_);
  and (_29581_, _29580_, _29578_);
  and (_29582_, _29336_, _10448_);
  or (_29583_, _29582_, _06260_);
  or (_29584_, _29583_, _29581_);
  nand (_29585_, _08209_, _06260_);
  and (_29586_, _29585_, _29584_);
  or (_29588_, _29586_, _12089_);
  nor (_29589_, _12113_, _05924_);
  nor (_29590_, _29589_, _06377_);
  and (_29591_, _29590_, _29588_);
  and (_29592_, _12253_, _12954_);
  nor (_29593_, _29355_, _12954_);
  or (_29594_, _29593_, _29592_);
  and (_29595_, _29594_, _06377_);
  or (_29596_, _29595_, _12985_);
  or (_29597_, _29596_, _29591_);
  or (_29599_, _29336_, _12984_);
  and (_29600_, _29599_, _07241_);
  and (_29601_, _29600_, _29597_);
  nand (_29602_, _12113_, _06563_);
  nand (_29603_, _29602_, _12991_);
  or (_29604_, _29603_, _29601_);
  or (_29605_, _29336_, _12991_);
  and (_29606_, _29605_, _08505_);
  and (_29607_, _29606_, _29604_);
  nor (_29608_, _06608_, _08505_);
  or (_29610_, _29608_, _05912_);
  or (_29611_, _29610_, _29607_);
  nand (_29612_, _15483_, _05912_);
  and (_29613_, _29612_, _06571_);
  and (_29614_, _29613_, _29611_);
  and (_29615_, _29594_, _06199_);
  or (_29616_, _29615_, _13007_);
  or (_29617_, _29616_, _29614_);
  or (_29618_, _29336_, _13006_);
  and (_29619_, _29618_, _06189_);
  and (_29621_, _29619_, _29617_);
  nand (_29622_, _12113_, _06188_);
  nand (_29623_, _29622_, _13013_);
  or (_29624_, _29623_, _29621_);
  or (_29625_, _29336_, _13013_);
  and (_29626_, _29625_, _13018_);
  and (_29627_, _29626_, _29624_);
  nor (_29628_, _06608_, _13018_);
  or (_29629_, _29628_, _05907_);
  or (_29630_, _29629_, _29627_);
  nand (_29632_, _15483_, _05907_);
  and (_29633_, _29632_, _13026_);
  and (_29634_, _29633_, _29630_);
  and (_29635_, _29336_, _13025_);
  or (_29636_, _29635_, _29634_);
  or (_29637_, _29636_, _01456_);
  or (_29638_, _01452_, \oc8051_golden_model_1.PC [13]);
  and (_29639_, _29638_, _43223_);
  and (_43869_, _29639_, _29637_);
  nand (_29640_, _06342_, _06326_);
  or (_29642_, _29333_, \oc8051_golden_model_1.PC [14]);
  and (_29643_, _29642_, _12099_);
  or (_29644_, _29643_, _12966_);
  nor (_29645_, _12747_, _15682_);
  nor (_29646_, _12719_, _15682_);
  nor (_29647_, _12697_, _15682_);
  nor (_29648_, _12673_, _15682_);
  or (_29649_, _12108_, _08972_);
  and (_29650_, _12392_, _12248_);
  nor (_29651_, _12353_, _12251_);
  nor (_29653_, _29651_, _12354_);
  and (_29654_, _29653_, _27122_);
  or (_29655_, _29654_, _29650_);
  or (_29656_, _29655_, _06345_);
  or (_29657_, _29643_, _12451_);
  and (_29658_, _29643_, _07134_);
  and (_29659_, _12412_, _12108_);
  nor (_29660_, _12205_, _12111_);
  nor (_29661_, _29660_, _12206_);
  and (_29662_, _29661_, _12414_);
  or (_29664_, _29662_, _29659_);
  or (_29665_, _29664_, _08573_);
  or (_29666_, _29643_, _12427_);
  nand (_29667_, _12427_, _15682_);
  and (_29668_, _29667_, _29666_);
  or (_29669_, _29668_, _25018_);
  and (_29670_, _29643_, _28416_);
  nand (_29671_, _15682_, _07123_);
  and (_29672_, _29671_, _12418_);
  and (_29673_, _12419_, \oc8051_golden_model_1.PC [14]);
  or (_29675_, _29673_, _07123_);
  and (_29676_, _29675_, _29672_);
  or (_29677_, _29676_, _06705_);
  or (_29678_, _29677_, _29670_);
  and (_29679_, _29678_, _29669_);
  or (_29680_, _29679_, _08572_);
  and (_29681_, _29680_, _07338_);
  and (_29682_, _29681_, _29665_);
  or (_29683_, _29682_, _29658_);
  or (_29684_, _29683_, _06251_);
  or (_29685_, _12404_, _12248_);
  or (_29686_, _29653_, _12402_);
  and (_29687_, _29686_, _29685_);
  or (_29688_, _29687_, _06252_);
  and (_29689_, _29688_, _29684_);
  or (_29690_, _29689_, _12444_);
  or (_29691_, _29643_, _12443_);
  and (_29692_, _29691_, _12447_);
  and (_29693_, _29692_, _29690_);
  nor (_29694_, _12447_, _15682_);
  or (_29697_, _29694_, _12452_);
  or (_29698_, _29697_, _29693_);
  and (_29699_, _29698_, _29657_);
  or (_29700_, _29699_, _06466_);
  nand (_29701_, _15682_, _06466_);
  and (_29702_, _29701_, _12462_);
  and (_29703_, _29702_, _29700_);
  and (_29704_, _29643_, _12464_);
  or (_29705_, _29704_, _29703_);
  and (_29706_, _29705_, _12468_);
  or (_29708_, _12468_, _15682_);
  nand (_29709_, _29708_, _12478_);
  or (_29710_, _29709_, _29706_);
  and (_29711_, _12513_, _12248_);
  and (_29712_, _29653_, _14042_);
  or (_29713_, _29712_, _29711_);
  or (_29714_, _29713_, _12478_);
  and (_29715_, _29714_, _29710_);
  or (_29716_, _29715_, _06344_);
  and (_29717_, _29716_, _29656_);
  or (_29719_, _29717_, _06338_);
  and (_29720_, _29653_, _12534_);
  and (_29721_, _12533_, _12248_);
  or (_29722_, _29721_, _12536_);
  or (_29723_, _29722_, _29720_);
  and (_29724_, _29723_, _12522_);
  and (_29725_, _29724_, _29719_);
  or (_29726_, _29653_, _12555_);
  or (_29727_, _28800_, _12248_);
  and (_29728_, _29727_, _06373_);
  and (_29730_, _29728_, _29726_);
  or (_29731_, _29730_, _12245_);
  or (_29732_, _29731_, _29725_);
  or (_29733_, _29643_, _12246_);
  and (_29734_, _29733_, _12573_);
  and (_29735_, _29734_, _29732_);
  nor (_29736_, _12573_, _15682_);
  or (_29737_, _29736_, _12243_);
  or (_29738_, _29737_, _29735_);
  or (_29739_, _29643_, _12242_);
  and (_29741_, _29739_, _12580_);
  and (_29742_, _29741_, _29738_);
  nor (_29743_, _12580_, _15682_);
  or (_29744_, _29743_, _12582_);
  or (_29745_, _29744_, _29742_);
  or (_29746_, _29643_, _12237_);
  and (_29747_, _29746_, _12588_);
  and (_29748_, _29747_, _29745_);
  nor (_29749_, _12588_, _15682_);
  or (_29750_, _29749_, _05976_);
  or (_29752_, _29750_, _29748_);
  or (_29753_, _29643_, _05977_);
  and (_29754_, _29753_, _12595_);
  and (_29755_, _29754_, _29752_);
  nor (_29756_, _12595_, _15682_);
  or (_29757_, _29756_, _06369_);
  or (_29758_, _29757_, _29755_);
  or (_29759_, _12248_, _06370_);
  and (_29760_, _29759_, _12603_);
  and (_29761_, _29760_, _29758_);
  nor (_29763_, _12603_, _15682_);
  or (_29764_, _29763_, _05968_);
  or (_29765_, _29764_, _29761_);
  or (_29766_, _12248_, _06336_);
  and (_29767_, _29766_, _12611_);
  and (_29768_, _29767_, _29765_);
  and (_29769_, _29643_, _12615_);
  or (_29770_, _29769_, _12614_);
  or (_29771_, _29770_, _29768_);
  or (_29772_, _12613_, _12108_);
  and (_29774_, _29772_, _12620_);
  and (_29775_, _29774_, _29771_);
  and (_29776_, _29661_, _12619_);
  or (_29777_, _29776_, _08973_);
  or (_29778_, _29777_, _29775_);
  and (_29779_, _29778_, _29649_);
  or (_29780_, _29779_, _06371_);
  or (_29781_, _12248_, _07198_);
  and (_29782_, _29781_, _10905_);
  and (_29783_, _29782_, _29780_);
  and (_29785_, _12108_, _10904_);
  or (_29786_, _29785_, _12634_);
  or (_29787_, _29786_, _29783_);
  nor (_29788_, _12667_, \oc8051_golden_model_1.DPH [6]);
  nor (_29789_, _29788_, _12668_);
  or (_29790_, _29789_, _12635_);
  and (_29791_, _29790_, _12673_);
  and (_29792_, _29791_, _29787_);
  or (_29793_, _29792_, _29648_);
  and (_29794_, _29793_, _12678_);
  or (_29796_, _29661_, _11291_);
  or (_29797_, _12108_, _12684_);
  and (_29798_, _29797_, _12677_);
  and (_29799_, _29798_, _29796_);
  or (_29800_, _29799_, _12682_);
  or (_29801_, _29800_, _29794_);
  or (_29802_, _29643_, _12232_);
  and (_29803_, _29802_, _12228_);
  and (_29804_, _29803_, _29801_);
  nor (_29805_, _15682_, _12228_);
  or (_29807_, _29805_, _06367_);
  or (_29808_, _29807_, _29804_);
  or (_29809_, _12248_, _07218_);
  and (_29810_, _29809_, _12697_);
  and (_29811_, _29810_, _29808_);
  or (_29812_, _29811_, _29647_);
  and (_29813_, _29812_, _12702_);
  or (_29814_, _29661_, _12684_);
  or (_29815_, _12108_, _11291_);
  and (_29816_, _29815_, _12701_);
  and (_29818_, _29816_, _29814_);
  or (_29819_, _29818_, _12710_);
  or (_29820_, _29819_, _29813_);
  or (_29821_, _29643_, _12226_);
  and (_29822_, _29821_, _10967_);
  and (_29823_, _29822_, _29820_);
  nor (_29824_, _15682_, _10967_);
  or (_29825_, _29824_, _06366_);
  or (_29826_, _29825_, _29823_);
  or (_29827_, _12248_, _07213_);
  and (_29829_, _29827_, _12719_);
  and (_29830_, _29829_, _29826_);
  or (_29831_, _29830_, _29646_);
  and (_29832_, _29831_, _12724_);
  or (_29833_, _29661_, \oc8051_golden_model_1.PSW [7]);
  or (_29834_, _12108_, _10854_);
  and (_29835_, _29834_, _12723_);
  and (_29836_, _29835_, _29833_);
  or (_29837_, _29836_, _12738_);
  or (_29838_, _29837_, _29832_);
  or (_29840_, _29643_, _12736_);
  and (_29841_, _29840_, _11005_);
  and (_29842_, _29841_, _29838_);
  nor (_29843_, _15682_, _11005_);
  or (_29844_, _29843_, _06383_);
  or (_29845_, _29844_, _29842_);
  or (_29846_, _12248_, _07231_);
  and (_29847_, _29846_, _12747_);
  and (_29848_, _29847_, _29845_);
  or (_29849_, _29848_, _29645_);
  and (_29851_, _29849_, _12751_);
  or (_29852_, _29661_, _10854_);
  or (_29853_, _12108_, \oc8051_golden_model_1.PSW [7]);
  and (_29854_, _29853_, _12215_);
  and (_29855_, _29854_, _29852_);
  or (_29856_, _29855_, _12758_);
  or (_29857_, _29856_, _29851_);
  or (_29858_, _29643_, _12756_);
  and (_29859_, _29858_, _11051_);
  and (_29860_, _29859_, _29857_);
  nor (_29862_, _15682_, _11051_);
  or (_29863_, _29862_, _11080_);
  or (_29864_, _29863_, _29860_);
  or (_29865_, _29643_, _11081_);
  and (_29866_, _29865_, _13873_);
  and (_29867_, _29866_, _29864_);
  nor (_29868_, _08106_, _13873_);
  or (_29869_, _29868_, _07228_);
  or (_29870_, _29869_, _29867_);
  nor (_29871_, _12108_, _05916_);
  nor (_29873_, _29871_, _06381_);
  and (_29874_, _29873_, _29870_);
  or (_29875_, _29653_, _12955_);
  or (_29876_, _12248_, _12954_);
  and (_29877_, _29876_, _06381_);
  and (_29878_, _29877_, _29875_);
  or (_29879_, _29878_, _12774_);
  or (_29880_, _29879_, _29874_);
  or (_29881_, _29643_, _12105_);
  and (_29882_, _29881_, _12963_);
  and (_29884_, _29882_, _29880_);
  nor (_29885_, _12963_, _15682_);
  or (_29886_, _29885_, _10448_);
  or (_29887_, _29886_, _29884_);
  and (_29888_, _29887_, _29644_);
  or (_29889_, _29888_, _06260_);
  nand (_29890_, _08106_, _06260_);
  and (_29891_, _29890_, _05924_);
  and (_29892_, _29891_, _29889_);
  nor (_29893_, _15682_, _05924_);
  or (_29895_, _29893_, _06377_);
  or (_29896_, _29895_, _29892_);
  or (_29897_, _12248_, _12955_);
  or (_29898_, _29653_, _12954_);
  and (_29899_, _29898_, _29897_);
  or (_29900_, _29899_, _06564_);
  and (_29901_, _29900_, _29896_);
  or (_29902_, _29901_, _12985_);
  or (_29903_, _29643_, _12984_);
  and (_29904_, _29903_, _29902_);
  or (_29906_, _29904_, _06563_);
  nand (_29907_, _15682_, _06563_);
  and (_29908_, _29907_, _12991_);
  and (_29909_, _29908_, _29906_);
  and (_29910_, _29643_, _12992_);
  or (_29911_, _29910_, _06378_);
  or (_29912_, _29911_, _29909_);
  nand (_29913_, _06378_, _06326_);
  and (_29914_, _29913_, _05913_);
  and (_29915_, _29914_, _29912_);
  and (_29917_, _12108_, _05912_);
  or (_29918_, _29917_, _06199_);
  or (_29919_, _29918_, _29915_);
  or (_29920_, _29899_, _06571_);
  and (_29921_, _29920_, _13006_);
  and (_29922_, _29921_, _29919_);
  and (_29923_, _29643_, _13007_);
  or (_29924_, _29923_, _06188_);
  or (_29925_, _29924_, _29922_);
  nand (_29926_, _15682_, _06188_);
  and (_29928_, _29926_, _13013_);
  and (_29929_, _29928_, _29925_);
  and (_29930_, _29643_, _13014_);
  or (_29931_, _29930_, _06342_);
  or (_29932_, _29931_, _29929_);
  and (_29933_, _29932_, _29640_);
  or (_29934_, _29933_, _05907_);
  nand (_29935_, _15682_, _05907_);
  and (_29936_, _29935_, _13026_);
  and (_29937_, _29936_, _29934_);
  and (_29939_, _29643_, _13025_);
  or (_29940_, _29939_, _29937_);
  or (_29941_, _29940_, _01456_);
  or (_29942_, _01452_, \oc8051_golden_model_1.PC [14]);
  and (_29943_, _29942_, _43223_);
  and (_43870_, _29943_, _29941_);
  nand (_29944_, _11218_, _07881_);
  and (_29945_, _13035_, \oc8051_golden_model_1.P2 [0]);
  nor (_29946_, _29945_, _07210_);
  nand (_29947_, _29946_, _29944_);
  and (_29949_, _07881_, _07325_);
  or (_29950_, _29949_, _29945_);
  or (_29951_, _29950_, _07188_);
  and (_29952_, _13043_, \oc8051_golden_model_1.P2 [0]);
  and (_29953_, _14341_, _08535_);
  or (_29954_, _29953_, _29952_);
  and (_29955_, _29954_, _06475_);
  nor (_29956_, _08351_, _13035_);
  or (_29957_, _29956_, _29945_);
  or (_29958_, _29957_, _06252_);
  and (_29960_, _07881_, \oc8051_golden_model_1.ACC [0]);
  or (_29961_, _29960_, _29945_);
  and (_29962_, _29961_, _07123_);
  and (_29963_, _07124_, \oc8051_golden_model_1.P2 [0]);
  or (_29964_, _29963_, _06251_);
  or (_29965_, _29964_, _29962_);
  and (_29966_, _29965_, _06476_);
  and (_29967_, _29966_, _29958_);
  or (_29968_, _29967_, _29955_);
  and (_29969_, _29968_, _07142_);
  and (_29971_, _29950_, _06468_);
  or (_29972_, _29971_, _06466_);
  or (_29973_, _29972_, _29969_);
  or (_29974_, _29961_, _06801_);
  and (_29975_, _29974_, _06484_);
  and (_29976_, _29975_, _29973_);
  and (_29977_, _29945_, _06483_);
  or (_29978_, _29977_, _06461_);
  or (_29979_, _29978_, _29976_);
  or (_29980_, _29957_, _07164_);
  and (_29982_, _29980_, _06242_);
  and (_29983_, _29982_, _29979_);
  or (_29984_, _29952_, _14371_);
  and (_29985_, _29984_, _06241_);
  and (_29986_, _29985_, _29954_);
  or (_29987_, _29986_, _07187_);
  or (_29988_, _29987_, _29983_);
  and (_29989_, _29988_, _29951_);
  or (_29990_, _29989_, _07182_);
  and (_29991_, _09342_, _07881_);
  or (_29993_, _29945_, _07183_);
  or (_29994_, _29993_, _29991_);
  and (_29995_, _29994_, _29990_);
  or (_29996_, _29995_, _05968_);
  and (_29997_, _14427_, _07881_);
  or (_29998_, _29945_, _06336_);
  or (_29999_, _29998_, _29997_);
  and (_30000_, _29999_, _07198_);
  and (_30001_, _30000_, _29996_);
  and (_30002_, _07881_, _08908_);
  or (_30004_, _30002_, _29945_);
  and (_30005_, _30004_, _06371_);
  or (_30006_, _30005_, _06367_);
  or (_30007_, _30006_, _30001_);
  and (_30008_, _14442_, _07881_);
  or (_30009_, _30008_, _29945_);
  or (_30010_, _30009_, _07218_);
  and (_30011_, _30010_, _07216_);
  and (_30012_, _30011_, _30007_);
  nor (_30013_, _12526_, _13035_);
  or (_30015_, _30013_, _29945_);
  and (_30016_, _29944_, _06533_);
  and (_30017_, _30016_, _30015_);
  or (_30018_, _30017_, _30012_);
  and (_30019_, _30018_, _07213_);
  nand (_30020_, _30004_, _06366_);
  nor (_30021_, _30020_, _29956_);
  or (_30022_, _30021_, _06541_);
  or (_30023_, _30022_, _30019_);
  and (_30024_, _30023_, _29947_);
  or (_30026_, _30024_, _06383_);
  and (_30027_, _14325_, _07881_);
  or (_30028_, _29945_, _07231_);
  or (_30029_, _30028_, _30027_);
  and (_30030_, _30029_, _07229_);
  and (_30031_, _30030_, _30026_);
  and (_30032_, _30015_, _06528_);
  or (_30033_, _30032_, _06563_);
  or (_30034_, _30033_, _30031_);
  or (_30035_, _29957_, _07241_);
  and (_30037_, _30035_, _30034_);
  or (_30038_, _30037_, _06199_);
  or (_30039_, _29945_, _06571_);
  and (_30040_, _30039_, _30038_);
  or (_30041_, _30040_, _06188_);
  or (_30042_, _29957_, _06189_);
  and (_30043_, _30042_, _01452_);
  and (_30044_, _30043_, _30041_);
  nor (_30045_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_30046_, _30045_, _00000_);
  or (_43871_, _30046_, _30044_);
  nor (_30048_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_30049_, _30048_, _00000_);
  and (_30050_, _13035_, \oc8051_golden_model_1.P2 [1]);
  nor (_30051_, _11216_, _13035_);
  or (_30052_, _30051_, _30050_);
  or (_30053_, _30052_, _07229_);
  nand (_30054_, _07881_, _07018_);
  or (_30055_, _07881_, \oc8051_golden_model_1.P2 [1]);
  and (_30056_, _30055_, _06371_);
  and (_30058_, _30056_, _30054_);
  and (_30059_, _14503_, _07881_);
  not (_30060_, _30059_);
  and (_30061_, _30060_, _30055_);
  and (_30062_, _30061_, _06251_);
  and (_30063_, _07124_, \oc8051_golden_model_1.P2 [1]);
  and (_30064_, _07881_, \oc8051_golden_model_1.ACC [1]);
  or (_30065_, _30064_, _30050_);
  and (_30066_, _30065_, _07123_);
  or (_30067_, _30066_, _30063_);
  and (_30069_, _30067_, _06252_);
  or (_30070_, _30069_, _06475_);
  or (_30071_, _30070_, _30062_);
  and (_30072_, _13043_, \oc8051_golden_model_1.P2 [1]);
  and (_30073_, _14510_, _08535_);
  or (_30074_, _30073_, _30072_);
  or (_30075_, _30074_, _06476_);
  and (_30076_, _30075_, _30071_);
  or (_30077_, _30076_, _06468_);
  nor (_30078_, _13035_, _07120_);
  or (_30080_, _30078_, _30050_);
  or (_30081_, _30080_, _07142_);
  and (_30082_, _30081_, _30077_);
  or (_30083_, _30082_, _06466_);
  or (_30084_, _30065_, _06801_);
  and (_30085_, _30084_, _06484_);
  and (_30086_, _30085_, _30083_);
  and (_30087_, _14513_, _08535_);
  or (_30088_, _30087_, _30072_);
  and (_30089_, _30088_, _06483_);
  or (_30091_, _30089_, _06461_);
  or (_30092_, _30091_, _30086_);
  or (_30093_, _30072_, _14509_);
  and (_30094_, _30093_, _30074_);
  or (_30095_, _30094_, _07164_);
  and (_30096_, _30095_, _06242_);
  and (_30097_, _30096_, _30092_);
  or (_30098_, _30072_, _14553_);
  and (_30099_, _30098_, _06241_);
  and (_30100_, _30099_, _30074_);
  or (_30102_, _30100_, _07187_);
  or (_30103_, _30102_, _30097_);
  or (_30104_, _30080_, _07188_);
  and (_30105_, _30104_, _30103_);
  or (_30106_, _30105_, _07182_);
  and (_30107_, _09297_, _07881_);
  or (_30108_, _30050_, _07183_);
  or (_30109_, _30108_, _30107_);
  and (_30110_, _30109_, _06336_);
  and (_30111_, _30110_, _30106_);
  and (_30113_, _14609_, _07881_);
  or (_30114_, _30113_, _30050_);
  and (_30115_, _30114_, _05968_);
  or (_30116_, _30115_, _30111_);
  and (_30117_, _30116_, _07198_);
  or (_30118_, _30117_, _30058_);
  and (_30119_, _30118_, _07218_);
  or (_30120_, _14625_, _13035_);
  and (_30121_, _30055_, _06367_);
  and (_30122_, _30121_, _30120_);
  or (_30124_, _30122_, _06533_);
  or (_30125_, _30124_, _30119_);
  nand (_30126_, _11215_, _07881_);
  and (_30127_, _30126_, _30052_);
  or (_30128_, _30127_, _07216_);
  and (_30129_, _30128_, _07213_);
  and (_30130_, _30129_, _30125_);
  or (_30131_, _14623_, _13035_);
  and (_30132_, _30055_, _06366_);
  and (_30133_, _30132_, _30131_);
  or (_30135_, _30133_, _06541_);
  or (_30136_, _30135_, _30130_);
  nor (_30137_, _30050_, _07210_);
  nand (_30138_, _30137_, _30126_);
  and (_30139_, _30138_, _07231_);
  and (_30140_, _30139_, _30136_);
  or (_30141_, _30054_, _08302_);
  and (_30142_, _30055_, _06383_);
  and (_30143_, _30142_, _30141_);
  or (_30144_, _30143_, _06528_);
  or (_30146_, _30144_, _30140_);
  and (_30147_, _30146_, _30053_);
  or (_30148_, _30147_, _06563_);
  or (_30149_, _30061_, _07241_);
  and (_30150_, _30149_, _06571_);
  and (_30151_, _30150_, _30148_);
  and (_30152_, _30088_, _06199_);
  or (_30153_, _30152_, _06188_);
  or (_30154_, _30153_, _30151_);
  or (_30155_, _30050_, _06189_);
  or (_30157_, _30155_, _30059_);
  and (_30158_, _30157_, _01452_);
  and (_30159_, _30158_, _30154_);
  or (_43873_, _30159_, _30049_);
  and (_30160_, _13035_, \oc8051_golden_model_1.P2 [2]);
  nor (_30161_, _13035_, _07578_);
  or (_30162_, _30161_, _30160_);
  or (_30163_, _30162_, _07188_);
  and (_30164_, _14712_, _07881_);
  or (_30165_, _30164_, _30160_);
  or (_30167_, _30165_, _06252_);
  and (_30168_, _07881_, \oc8051_golden_model_1.ACC [2]);
  or (_30169_, _30168_, _30160_);
  and (_30170_, _30169_, _07123_);
  and (_30171_, _07124_, \oc8051_golden_model_1.P2 [2]);
  or (_30172_, _30171_, _06251_);
  or (_30173_, _30172_, _30170_);
  and (_30174_, _30173_, _06476_);
  and (_30175_, _30174_, _30167_);
  and (_30176_, _13043_, \oc8051_golden_model_1.P2 [2]);
  and (_30178_, _14702_, _08535_);
  or (_30179_, _30178_, _30176_);
  and (_30180_, _30179_, _06475_);
  or (_30181_, _30180_, _06468_);
  or (_30182_, _30181_, _30175_);
  or (_30183_, _30162_, _07142_);
  and (_30184_, _30183_, _30182_);
  or (_30185_, _30184_, _06466_);
  or (_30186_, _30169_, _06801_);
  and (_30187_, _30186_, _06484_);
  and (_30189_, _30187_, _30185_);
  and (_30190_, _14706_, _08535_);
  or (_30191_, _30190_, _30176_);
  and (_30192_, _30191_, _06483_);
  or (_30193_, _30192_, _06461_);
  or (_30194_, _30193_, _30189_);
  or (_30195_, _30176_, _14739_);
  and (_30196_, _30195_, _30179_);
  or (_30197_, _30196_, _07164_);
  and (_30198_, _30197_, _06242_);
  and (_30200_, _30198_, _30194_);
  or (_30201_, _30176_, _14703_);
  and (_30202_, _30201_, _06241_);
  and (_30203_, _30202_, _30179_);
  or (_30204_, _30203_, _07187_);
  or (_30205_, _30204_, _30200_);
  and (_30206_, _30205_, _30163_);
  or (_30207_, _30206_, _07182_);
  and (_30208_, _09251_, _07881_);
  or (_30209_, _30160_, _07183_);
  or (_30211_, _30209_, _30208_);
  and (_30212_, _30211_, _06336_);
  and (_30213_, _30212_, _30207_);
  and (_30214_, _14808_, _07881_);
  or (_30215_, _30214_, _30160_);
  and (_30216_, _30215_, _05968_);
  or (_30217_, _30216_, _06371_);
  or (_30218_, _30217_, _30213_);
  and (_30219_, _07881_, _08945_);
  or (_30220_, _30219_, _30160_);
  or (_30222_, _30220_, _07198_);
  and (_30223_, _30222_, _30218_);
  or (_30224_, _30223_, _06367_);
  and (_30225_, _14824_, _07881_);
  or (_30226_, _30225_, _30160_);
  or (_30227_, _30226_, _07218_);
  and (_30228_, _30227_, _07216_);
  and (_30229_, _30228_, _30224_);
  and (_30230_, _11214_, _07881_);
  or (_30231_, _30230_, _30160_);
  and (_30233_, _30231_, _06533_);
  or (_30234_, _30233_, _30229_);
  and (_30235_, _30234_, _07213_);
  or (_30236_, _30160_, _08397_);
  and (_30237_, _30220_, _06366_);
  and (_30238_, _30237_, _30236_);
  or (_30239_, _30238_, _30235_);
  and (_30240_, _30239_, _07210_);
  and (_30241_, _30169_, _06541_);
  and (_30242_, _30241_, _30236_);
  or (_30244_, _30242_, _06383_);
  or (_30245_, _30244_, _30240_);
  and (_30246_, _14821_, _07881_);
  or (_30247_, _30160_, _07231_);
  or (_30248_, _30247_, _30246_);
  and (_30249_, _30248_, _07229_);
  and (_30250_, _30249_, _30245_);
  nor (_30251_, _11213_, _13035_);
  or (_30252_, _30251_, _30160_);
  and (_30253_, _30252_, _06528_);
  or (_30255_, _30253_, _06563_);
  or (_30256_, _30255_, _30250_);
  or (_30257_, _30165_, _07241_);
  and (_30258_, _30257_, _06571_);
  and (_30259_, _30258_, _30256_);
  and (_30260_, _30191_, _06199_);
  or (_30261_, _30260_, _06188_);
  or (_30262_, _30261_, _30259_);
  and (_30263_, _14884_, _07881_);
  or (_30264_, _30160_, _06189_);
  or (_30266_, _30264_, _30263_);
  and (_30267_, _30266_, _01452_);
  and (_30268_, _30267_, _30262_);
  nor (_30269_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_30270_, _30269_, _00000_);
  or (_43874_, _30270_, _30268_);
  and (_30271_, _13035_, \oc8051_golden_model_1.P2 [3]);
  nor (_30272_, _13035_, _07713_);
  or (_30273_, _30272_, _30271_);
  or (_30274_, _30273_, _07188_);
  or (_30276_, _30273_, _07142_);
  and (_30277_, _14898_, _07881_);
  or (_30278_, _30277_, _30271_);
  or (_30279_, _30278_, _06252_);
  and (_30280_, _07881_, \oc8051_golden_model_1.ACC [3]);
  or (_30281_, _30280_, _30271_);
  and (_30282_, _30281_, _07123_);
  and (_30283_, _07124_, \oc8051_golden_model_1.P2 [3]);
  or (_30284_, _30283_, _06251_);
  or (_30285_, _30284_, _30282_);
  and (_30287_, _30285_, _06476_);
  and (_30288_, _30287_, _30279_);
  and (_30289_, _13043_, \oc8051_golden_model_1.P2 [3]);
  and (_30290_, _14906_, _08535_);
  or (_30291_, _30290_, _30289_);
  and (_30292_, _30291_, _06475_);
  or (_30293_, _30292_, _06468_);
  or (_30294_, _30293_, _30288_);
  and (_30295_, _30294_, _30276_);
  or (_30296_, _30295_, _06466_);
  or (_30298_, _30281_, _06801_);
  and (_30299_, _30298_, _06484_);
  and (_30300_, _30299_, _30296_);
  and (_30301_, _14904_, _08535_);
  or (_30302_, _30301_, _30289_);
  and (_30303_, _30302_, _06483_);
  or (_30304_, _30303_, _06461_);
  or (_30305_, _30304_, _30300_);
  or (_30306_, _30289_, _14931_);
  and (_30307_, _30306_, _30291_);
  or (_30308_, _30307_, _07164_);
  and (_30309_, _30308_, _06242_);
  and (_30310_, _30309_, _30305_);
  or (_30311_, _30289_, _14947_);
  and (_30312_, _30311_, _06241_);
  and (_30313_, _30312_, _30291_);
  or (_30314_, _30313_, _07187_);
  or (_30315_, _30314_, _30310_);
  and (_30316_, _30315_, _30274_);
  or (_30317_, _30316_, _07182_);
  and (_30320_, _09205_, _07881_);
  or (_30321_, _30271_, _07183_);
  or (_30322_, _30321_, _30320_);
  and (_30323_, _30322_, _06336_);
  and (_30324_, _30323_, _30317_);
  and (_30325_, _15003_, _07881_);
  or (_30326_, _30325_, _30271_);
  and (_30327_, _30326_, _05968_);
  or (_30328_, _30327_, _06371_);
  or (_30329_, _30328_, _30324_);
  and (_30331_, _07881_, _08872_);
  or (_30332_, _30331_, _30271_);
  or (_30333_, _30332_, _07198_);
  and (_30334_, _30333_, _30329_);
  or (_30335_, _30334_, _06367_);
  and (_30336_, _15018_, _07881_);
  or (_30337_, _30336_, _30271_);
  or (_30338_, _30337_, _07218_);
  and (_30339_, _30338_, _07216_);
  and (_30340_, _30339_, _30335_);
  and (_30342_, _12523_, _07881_);
  or (_30343_, _30342_, _30271_);
  and (_30344_, _30343_, _06533_);
  or (_30345_, _30344_, _30340_);
  and (_30346_, _30345_, _07213_);
  or (_30347_, _30271_, _08257_);
  and (_30348_, _30332_, _06366_);
  and (_30349_, _30348_, _30347_);
  or (_30350_, _30349_, _30346_);
  and (_30351_, _30350_, _07210_);
  and (_30353_, _30281_, _06541_);
  and (_30354_, _30353_, _30347_);
  or (_30355_, _30354_, _06383_);
  or (_30356_, _30355_, _30351_);
  and (_30357_, _15015_, _07881_);
  or (_30358_, _30271_, _07231_);
  or (_30359_, _30358_, _30357_);
  and (_30360_, _30359_, _07229_);
  and (_30361_, _30360_, _30356_);
  nor (_30362_, _11211_, _13035_);
  or (_30364_, _30362_, _30271_);
  and (_30365_, _30364_, _06528_);
  or (_30366_, _30365_, _06563_);
  or (_30367_, _30366_, _30361_);
  or (_30368_, _30278_, _07241_);
  and (_30369_, _30368_, _06571_);
  and (_30370_, _30369_, _30367_);
  and (_30371_, _30302_, _06199_);
  or (_30372_, _30371_, _06188_);
  or (_30373_, _30372_, _30370_);
  and (_30375_, _15075_, _07881_);
  or (_30376_, _30271_, _06189_);
  or (_30377_, _30376_, _30375_);
  and (_30378_, _30377_, _01452_);
  and (_30379_, _30378_, _30373_);
  nor (_30380_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_30381_, _30380_, _00000_);
  or (_43875_, _30381_, _30379_);
  nor (_30382_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_30383_, _30382_, _00000_);
  and (_30385_, _13035_, \oc8051_golden_model_1.P2 [4]);
  nor (_30386_, _08494_, _13035_);
  or (_30387_, _30386_, _30385_);
  or (_30388_, _30387_, _07188_);
  and (_30389_, _13043_, \oc8051_golden_model_1.P2 [4]);
  and (_30390_, _15089_, _08535_);
  or (_30391_, _30390_, _30389_);
  and (_30392_, _30391_, _06483_);
  or (_30393_, _30387_, _07142_);
  and (_30394_, _15108_, _07881_);
  or (_30396_, _30394_, _30385_);
  or (_30397_, _30396_, _06252_);
  and (_30398_, _07881_, \oc8051_golden_model_1.ACC [4]);
  or (_30399_, _30398_, _30385_);
  and (_30400_, _30399_, _07123_);
  and (_30401_, _07124_, \oc8051_golden_model_1.P2 [4]);
  or (_30402_, _30401_, _06251_);
  or (_30403_, _30402_, _30400_);
  and (_30404_, _30403_, _06476_);
  and (_30405_, _30404_, _30397_);
  and (_30407_, _15091_, _08535_);
  or (_30408_, _30407_, _30389_);
  and (_30409_, _30408_, _06475_);
  or (_30410_, _30409_, _06468_);
  or (_30411_, _30410_, _30405_);
  and (_30412_, _30411_, _30393_);
  or (_30413_, _30412_, _06466_);
  or (_30414_, _30399_, _06801_);
  and (_30415_, _30414_, _06484_);
  and (_30416_, _30415_, _30413_);
  or (_30418_, _30416_, _30392_);
  and (_30419_, _30418_, _07164_);
  or (_30420_, _30389_, _15125_);
  and (_30421_, _30408_, _06461_);
  and (_30422_, _30421_, _30420_);
  or (_30423_, _30422_, _30419_);
  and (_30424_, _30423_, _06242_);
  or (_30425_, _30389_, _15141_);
  and (_30426_, _30425_, _06241_);
  and (_30427_, _30426_, _30408_);
  or (_30429_, _30427_, _07187_);
  or (_30430_, _30429_, _30424_);
  and (_30431_, _30430_, _30388_);
  or (_30432_, _30431_, _07182_);
  and (_30433_, _09159_, _07881_);
  or (_30434_, _30385_, _07183_);
  or (_30435_, _30434_, _30433_);
  and (_30436_, _30435_, _06336_);
  and (_30437_, _30436_, _30432_);
  and (_30438_, _15198_, _07881_);
  or (_30440_, _30438_, _30385_);
  and (_30441_, _30440_, _05968_);
  or (_30442_, _30441_, _06371_);
  or (_30443_, _30442_, _30437_);
  and (_30444_, _08892_, _07881_);
  or (_30445_, _30444_, _30385_);
  or (_30446_, _30445_, _07198_);
  and (_30447_, _30446_, _30443_);
  or (_30448_, _30447_, _06367_);
  and (_30449_, _15214_, _07881_);
  or (_30451_, _30449_, _30385_);
  or (_30452_, _30451_, _07218_);
  and (_30453_, _30452_, _07216_);
  and (_30454_, _30453_, _30448_);
  and (_30455_, _11209_, _07881_);
  or (_30456_, _30455_, _30385_);
  and (_30457_, _30456_, _06533_);
  or (_30458_, _30457_, _30454_);
  and (_30459_, _30458_, _07213_);
  or (_30460_, _30385_, _08497_);
  and (_30462_, _30445_, _06366_);
  and (_30463_, _30462_, _30460_);
  or (_30464_, _30463_, _30459_);
  and (_30465_, _30464_, _07210_);
  and (_30466_, _30399_, _06541_);
  and (_30467_, _30466_, _30460_);
  or (_30468_, _30467_, _06383_);
  or (_30469_, _30468_, _30465_);
  and (_30470_, _15211_, _07881_);
  or (_30471_, _30385_, _07231_);
  or (_30473_, _30471_, _30470_);
  and (_30474_, _30473_, _07229_);
  and (_30475_, _30474_, _30469_);
  nor (_30476_, _11208_, _13035_);
  or (_30477_, _30476_, _30385_);
  and (_30478_, _30477_, _06528_);
  or (_30479_, _30478_, _06563_);
  or (_30480_, _30479_, _30475_);
  or (_30481_, _30396_, _07241_);
  and (_30482_, _30481_, _06571_);
  and (_30484_, _30482_, _30480_);
  and (_30485_, _30391_, _06199_);
  or (_30486_, _30485_, _06188_);
  or (_30487_, _30486_, _30484_);
  and (_30488_, _15280_, _07881_);
  or (_30489_, _30385_, _06189_);
  or (_30490_, _30489_, _30488_);
  and (_30491_, _30490_, _01452_);
  and (_30492_, _30491_, _30487_);
  or (_43876_, _30492_, _30383_);
  and (_30494_, _13035_, \oc8051_golden_model_1.P2 [5]);
  nor (_30495_, _08209_, _13035_);
  or (_30496_, _30495_, _30494_);
  or (_30497_, _30496_, _07142_);
  and (_30498_, _15311_, _07881_);
  or (_30499_, _30498_, _30494_);
  or (_30500_, _30499_, _06252_);
  and (_30501_, _07881_, \oc8051_golden_model_1.ACC [5]);
  or (_30502_, _30501_, _30494_);
  and (_30503_, _30502_, _07123_);
  and (_30505_, _07124_, \oc8051_golden_model_1.P2 [5]);
  or (_30506_, _30505_, _06251_);
  or (_30507_, _30506_, _30503_);
  and (_30508_, _30507_, _06476_);
  and (_30509_, _30508_, _30500_);
  and (_30510_, _13043_, \oc8051_golden_model_1.P2 [5]);
  and (_30511_, _15296_, _08535_);
  or (_30512_, _30511_, _30510_);
  and (_30513_, _30512_, _06475_);
  or (_30514_, _30513_, _06468_);
  or (_30516_, _30514_, _30509_);
  and (_30517_, _30516_, _30497_);
  or (_30518_, _30517_, _06466_);
  or (_30519_, _30502_, _06801_);
  and (_30520_, _30519_, _06484_);
  and (_30521_, _30520_, _30518_);
  and (_30522_, _15294_, _08535_);
  or (_30523_, _30522_, _30510_);
  and (_30524_, _30523_, _06483_);
  or (_30525_, _30524_, _06461_);
  or (_30527_, _30525_, _30521_);
  or (_30528_, _30510_, _15328_);
  and (_30529_, _30528_, _30512_);
  or (_30530_, _30529_, _07164_);
  and (_30531_, _30530_, _06242_);
  and (_30532_, _30531_, _30527_);
  or (_30533_, _30510_, _15344_);
  and (_30534_, _30533_, _06241_);
  and (_30535_, _30534_, _30512_);
  or (_30536_, _30535_, _07187_);
  or (_30538_, _30536_, _30532_);
  or (_30539_, _30496_, _07188_);
  and (_30540_, _30539_, _30538_);
  or (_30541_, _30540_, _07182_);
  and (_30542_, _09113_, _07881_);
  or (_30543_, _30494_, _07183_);
  or (_30544_, _30543_, _30542_);
  and (_30545_, _30544_, _06336_);
  and (_30546_, _30545_, _30541_);
  and (_30547_, _15400_, _07881_);
  or (_30549_, _30547_, _30494_);
  and (_30550_, _30549_, _05968_);
  or (_30551_, _30550_, _06371_);
  or (_30552_, _30551_, _30546_);
  and (_30553_, _08888_, _07881_);
  or (_30554_, _30553_, _30494_);
  or (_30555_, _30554_, _07198_);
  and (_30556_, _30555_, _30552_);
  or (_30557_, _30556_, _06367_);
  and (_30558_, _15416_, _07881_);
  or (_30560_, _30558_, _30494_);
  or (_30561_, _30560_, _07218_);
  and (_30562_, _30561_, _07216_);
  and (_30563_, _30562_, _30557_);
  and (_30564_, _11205_, _07881_);
  or (_30565_, _30564_, _30494_);
  and (_30566_, _30565_, _06533_);
  or (_30567_, _30566_, _30563_);
  and (_30568_, _30567_, _07213_);
  or (_30569_, _30494_, _08212_);
  and (_30571_, _30554_, _06366_);
  and (_30572_, _30571_, _30569_);
  or (_30573_, _30572_, _30568_);
  and (_30574_, _30573_, _07210_);
  and (_30575_, _30502_, _06541_);
  and (_30576_, _30575_, _30569_);
  or (_30577_, _30576_, _06383_);
  or (_30578_, _30577_, _30574_);
  and (_30579_, _15413_, _07881_);
  or (_30580_, _30494_, _07231_);
  or (_30582_, _30580_, _30579_);
  and (_30583_, _30582_, _07229_);
  and (_30584_, _30583_, _30578_);
  nor (_30585_, _11204_, _13035_);
  or (_30586_, _30585_, _30494_);
  and (_30587_, _30586_, _06528_);
  or (_30588_, _30587_, _06563_);
  or (_30589_, _30588_, _30584_);
  or (_30590_, _30499_, _07241_);
  and (_30591_, _30590_, _06571_);
  and (_30593_, _30591_, _30589_);
  and (_30594_, _30523_, _06199_);
  or (_30595_, _30594_, _06188_);
  or (_30596_, _30595_, _30593_);
  and (_30597_, _15477_, _07881_);
  or (_30598_, _30494_, _06189_);
  or (_30599_, _30598_, _30597_);
  and (_30600_, _30599_, _01452_);
  and (_30601_, _30600_, _30596_);
  nor (_30602_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_30604_, _30602_, _00000_);
  or (_43877_, _30604_, _30601_);
  nor (_30605_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_30606_, _30605_, _00000_);
  and (_30607_, _13035_, \oc8051_golden_model_1.P2 [6]);
  nor (_30608_, _08106_, _13035_);
  or (_30609_, _30608_, _30607_);
  or (_30610_, _30609_, _07142_);
  and (_30611_, _15512_, _07881_);
  or (_30612_, _30611_, _30607_);
  or (_30614_, _30612_, _06252_);
  and (_30615_, _07881_, \oc8051_golden_model_1.ACC [6]);
  or (_30616_, _30615_, _30607_);
  and (_30617_, _30616_, _07123_);
  and (_30618_, _07124_, \oc8051_golden_model_1.P2 [6]);
  or (_30619_, _30618_, _06251_);
  or (_30620_, _30619_, _30617_);
  and (_30621_, _30620_, _06476_);
  and (_30622_, _30621_, _30614_);
  and (_30623_, _13043_, \oc8051_golden_model_1.P2 [6]);
  and (_30625_, _15499_, _08535_);
  or (_30626_, _30625_, _30623_);
  and (_30627_, _30626_, _06475_);
  or (_30628_, _30627_, _06468_);
  or (_30629_, _30628_, _30622_);
  and (_30630_, _30629_, _30610_);
  or (_30631_, _30630_, _06466_);
  or (_30632_, _30616_, _06801_);
  and (_30633_, _30632_, _06484_);
  and (_30634_, _30633_, _30631_);
  and (_30636_, _15497_, _08535_);
  or (_30637_, _30636_, _30623_);
  and (_30638_, _30637_, _06483_);
  or (_30639_, _30638_, _06461_);
  or (_30640_, _30639_, _30634_);
  or (_30641_, _30623_, _15529_);
  and (_30642_, _30641_, _30626_);
  or (_30643_, _30642_, _07164_);
  and (_30644_, _30643_, _06242_);
  and (_30645_, _30644_, _30640_);
  or (_30647_, _30623_, _15545_);
  and (_30648_, _30647_, _06241_);
  and (_30649_, _30648_, _30626_);
  or (_30650_, _30649_, _07187_);
  or (_30651_, _30650_, _30645_);
  or (_30652_, _30609_, _07188_);
  and (_30653_, _30652_, _30651_);
  or (_30654_, _30653_, _07182_);
  and (_30655_, _09067_, _07881_);
  or (_30656_, _30607_, _07183_);
  or (_30658_, _30656_, _30655_);
  and (_30659_, _30658_, _06336_);
  and (_30660_, _30659_, _30654_);
  and (_30661_, _15601_, _07881_);
  or (_30662_, _30661_, _30607_);
  and (_30663_, _30662_, _05968_);
  or (_30664_, _30663_, _06371_);
  or (_30665_, _30664_, _30660_);
  and (_30666_, _15608_, _07881_);
  or (_30667_, _30666_, _30607_);
  or (_30669_, _30667_, _07198_);
  and (_30670_, _30669_, _30665_);
  or (_30671_, _30670_, _06367_);
  and (_30672_, _15618_, _07881_);
  or (_30673_, _30672_, _30607_);
  or (_30674_, _30673_, _07218_);
  and (_30675_, _30674_, _07216_);
  and (_30676_, _30675_, _30671_);
  and (_30677_, _11202_, _07881_);
  or (_30678_, _30677_, _30607_);
  and (_30680_, _30678_, _06533_);
  or (_30681_, _30680_, _30676_);
  and (_30682_, _30681_, _07213_);
  or (_30683_, _30607_, _08109_);
  and (_30684_, _30667_, _06366_);
  and (_30685_, _30684_, _30683_);
  or (_30686_, _30685_, _30682_);
  and (_30687_, _30686_, _07210_);
  and (_30688_, _30616_, _06541_);
  and (_30689_, _30688_, _30683_);
  or (_30691_, _30689_, _06383_);
  or (_30692_, _30691_, _30687_);
  and (_30693_, _15615_, _07881_);
  or (_30694_, _30607_, _07231_);
  or (_30695_, _30694_, _30693_);
  and (_30696_, _30695_, _07229_);
  and (_30697_, _30696_, _30692_);
  nor (_30698_, _11201_, _13035_);
  or (_30699_, _30698_, _30607_);
  and (_30700_, _30699_, _06528_);
  or (_30702_, _30700_, _06563_);
  or (_30703_, _30702_, _30697_);
  or (_30704_, _30612_, _07241_);
  and (_30705_, _30704_, _06571_);
  and (_30706_, _30705_, _30703_);
  and (_30707_, _30637_, _06199_);
  or (_30708_, _30707_, _06188_);
  or (_30709_, _30708_, _30706_);
  and (_30710_, _15676_, _07881_);
  or (_30711_, _30607_, _06189_);
  or (_30713_, _30711_, _30710_);
  and (_30714_, _30713_, _01452_);
  and (_30715_, _30714_, _30709_);
  or (_43878_, _30715_, _30606_);
  and (_30716_, _07871_, \oc8051_golden_model_1.ACC [0]);
  and (_30717_, _30716_, _08351_);
  and (_30718_, _13138_, \oc8051_golden_model_1.P3 [0]);
  or (_30719_, _30718_, _07210_);
  or (_30720_, _30719_, _30717_);
  and (_30721_, _07871_, _07325_);
  or (_30723_, _30721_, _30718_);
  or (_30724_, _30723_, _07188_);
  and (_30725_, _13146_, \oc8051_golden_model_1.P3 [0]);
  and (_30726_, _14341_, _08539_);
  or (_30727_, _30726_, _30725_);
  and (_30728_, _30727_, _06475_);
  nor (_30729_, _08351_, _13138_);
  or (_30730_, _30729_, _30718_);
  or (_30731_, _30730_, _06252_);
  or (_30732_, _30716_, _30718_);
  and (_30734_, _30732_, _07123_);
  and (_30735_, _07124_, \oc8051_golden_model_1.P3 [0]);
  or (_30736_, _30735_, _06251_);
  or (_30737_, _30736_, _30734_);
  and (_30738_, _30737_, _06476_);
  and (_30739_, _30738_, _30731_);
  or (_30740_, _30739_, _30728_);
  and (_30741_, _30740_, _07142_);
  and (_30742_, _30723_, _06468_);
  or (_30743_, _30742_, _06466_);
  or (_30745_, _30743_, _30741_);
  or (_30746_, _30732_, _06801_);
  and (_30747_, _30746_, _06484_);
  and (_30748_, _30747_, _30745_);
  and (_30749_, _30718_, _06483_);
  or (_30750_, _30749_, _06461_);
  or (_30751_, _30750_, _30748_);
  or (_30752_, _30730_, _07164_);
  and (_30753_, _30752_, _06242_);
  and (_30754_, _30753_, _30751_);
  or (_30756_, _30725_, _14371_);
  and (_30757_, _30756_, _06241_);
  and (_30758_, _30757_, _30727_);
  or (_30759_, _30758_, _07187_);
  or (_30760_, _30759_, _30754_);
  and (_30761_, _30760_, _30724_);
  or (_30762_, _30761_, _07182_);
  and (_30763_, _09342_, _07871_);
  or (_30764_, _30718_, _07183_);
  or (_30765_, _30764_, _30763_);
  and (_30767_, _30765_, _30762_);
  or (_30768_, _30767_, _05968_);
  and (_30769_, _14427_, _07871_);
  or (_30770_, _30718_, _06336_);
  or (_30771_, _30770_, _30769_);
  and (_30772_, _30771_, _07198_);
  and (_30773_, _30772_, _30768_);
  and (_30774_, _07871_, _08908_);
  or (_30775_, _30774_, _30718_);
  and (_30776_, _30775_, _06371_);
  or (_30778_, _30776_, _06367_);
  or (_30779_, _30778_, _30773_);
  and (_30780_, _14442_, _07871_);
  or (_30781_, _30780_, _30718_);
  or (_30782_, _30781_, _07218_);
  and (_30783_, _30782_, _07216_);
  and (_30784_, _30783_, _30779_);
  nor (_30785_, _12526_, _13138_);
  or (_30786_, _30785_, _30718_);
  nor (_30787_, _30717_, _07216_);
  and (_30789_, _30787_, _30786_);
  or (_30790_, _30789_, _30784_);
  and (_30791_, _30790_, _07213_);
  nand (_30792_, _30775_, _06366_);
  nor (_30793_, _30792_, _30729_);
  or (_30794_, _30793_, _06541_);
  or (_30795_, _30794_, _30791_);
  and (_30796_, _30795_, _30720_);
  or (_30797_, _30796_, _06383_);
  and (_30798_, _14325_, _07871_);
  or (_30800_, _30798_, _30718_);
  or (_30801_, _30800_, _07231_);
  and (_30802_, _30801_, _07229_);
  and (_30803_, _30802_, _30797_);
  and (_30804_, _30786_, _06528_);
  or (_30805_, _30804_, _06563_);
  or (_30806_, _30805_, _30803_);
  or (_30807_, _30730_, _07241_);
  and (_30808_, _30807_, _30806_);
  or (_30809_, _30808_, _06199_);
  or (_30811_, _30718_, _06571_);
  and (_30812_, _30811_, _30809_);
  or (_30813_, _30812_, _06188_);
  or (_30814_, _30730_, _06189_);
  and (_30815_, _30814_, _01452_);
  and (_30816_, _30815_, _30813_);
  nor (_30817_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_30818_, _30817_, _00000_);
  or (_43880_, _30818_, _30816_);
  and (_30819_, _13138_, \oc8051_golden_model_1.P3 [1]);
  nor (_30821_, _11216_, _13138_);
  or (_30822_, _30821_, _30819_);
  or (_30823_, _30822_, _07229_);
  nand (_30824_, _07871_, _07018_);
  or (_30825_, _07871_, \oc8051_golden_model_1.P3 [1]);
  and (_30826_, _30825_, _06371_);
  and (_30827_, _30826_, _30824_);
  nor (_30828_, _13138_, _07120_);
  or (_30829_, _30828_, _30819_);
  or (_30830_, _30829_, _07142_);
  and (_30832_, _14503_, _07871_);
  not (_30833_, _30832_);
  and (_30834_, _30833_, _30825_);
  or (_30835_, _30834_, _06252_);
  and (_30836_, _07871_, \oc8051_golden_model_1.ACC [1]);
  or (_30837_, _30836_, _30819_);
  and (_30838_, _30837_, _07123_);
  and (_30839_, _07124_, \oc8051_golden_model_1.P3 [1]);
  or (_30840_, _30839_, _06251_);
  or (_30841_, _30840_, _30838_);
  and (_30843_, _30841_, _06476_);
  and (_30844_, _30843_, _30835_);
  and (_30845_, _13146_, \oc8051_golden_model_1.P3 [1]);
  and (_30846_, _14510_, _08539_);
  or (_30847_, _30846_, _30845_);
  and (_30848_, _30847_, _06475_);
  or (_30849_, _30848_, _06468_);
  or (_30850_, _30849_, _30844_);
  and (_30851_, _30850_, _30830_);
  or (_30852_, _30851_, _06466_);
  or (_30854_, _30837_, _06801_);
  and (_30855_, _30854_, _06484_);
  and (_30856_, _30855_, _30852_);
  and (_30857_, _14513_, _08539_);
  or (_30858_, _30857_, _30845_);
  and (_30859_, _30858_, _06483_);
  or (_30860_, _30859_, _06461_);
  or (_30861_, _30860_, _30856_);
  or (_30862_, _30845_, _14509_);
  and (_30863_, _30862_, _30847_);
  or (_30865_, _30863_, _07164_);
  and (_30866_, _30865_, _06242_);
  and (_30867_, _30866_, _30861_);
  or (_30868_, _30845_, _14553_);
  and (_30869_, _30868_, _06241_);
  and (_30870_, _30869_, _30847_);
  or (_30871_, _30870_, _07187_);
  or (_30872_, _30871_, _30867_);
  or (_30873_, _30829_, _07188_);
  and (_30874_, _30873_, _30872_);
  or (_30876_, _30874_, _07182_);
  and (_30877_, _09297_, _07871_);
  or (_30878_, _30819_, _07183_);
  or (_30879_, _30878_, _30877_);
  and (_30880_, _30879_, _06336_);
  and (_30881_, _30880_, _30876_);
  and (_30882_, _14609_, _07871_);
  or (_30883_, _30882_, _30819_);
  and (_30884_, _30883_, _05968_);
  or (_30885_, _30884_, _30881_);
  and (_30887_, _30885_, _07198_);
  or (_30888_, _30887_, _30827_);
  and (_30889_, _30888_, _07218_);
  or (_30890_, _14625_, _13138_);
  and (_30891_, _30825_, _06367_);
  and (_30892_, _30891_, _30890_);
  or (_30893_, _30892_, _06533_);
  or (_30894_, _30893_, _30889_);
  and (_30895_, _11217_, _07871_);
  or (_30896_, _30895_, _30819_);
  or (_30898_, _30896_, _07216_);
  and (_30899_, _30898_, _07213_);
  and (_30900_, _30899_, _30894_);
  or (_30901_, _14623_, _13138_);
  and (_30902_, _30825_, _06366_);
  and (_30903_, _30902_, _30901_);
  or (_30904_, _30903_, _06541_);
  or (_30905_, _30904_, _30900_);
  and (_30906_, _30836_, _08302_);
  or (_30907_, _30819_, _07210_);
  or (_30909_, _30907_, _30906_);
  and (_30910_, _30909_, _07231_);
  and (_30911_, _30910_, _30905_);
  or (_30912_, _30824_, _08302_);
  and (_30913_, _30825_, _06383_);
  and (_30914_, _30913_, _30912_);
  or (_30915_, _30914_, _06528_);
  or (_30916_, _30915_, _30911_);
  and (_30917_, _30916_, _30823_);
  or (_30918_, _30917_, _06563_);
  or (_30920_, _30834_, _07241_);
  and (_30921_, _30920_, _06571_);
  and (_30922_, _30921_, _30918_);
  and (_30923_, _30858_, _06199_);
  or (_30924_, _30923_, _06188_);
  or (_30925_, _30924_, _30922_);
  or (_30926_, _30819_, _06189_);
  or (_30927_, _30926_, _30832_);
  and (_30928_, _30927_, _01452_);
  and (_30929_, _30928_, _30925_);
  nor (_30931_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_30932_, _30931_, _00000_);
  or (_43881_, _30932_, _30929_);
  and (_30933_, _13138_, \oc8051_golden_model_1.P3 [2]);
  nor (_30934_, _13138_, _07578_);
  or (_30935_, _30934_, _30933_);
  or (_30936_, _30935_, _07188_);
  and (_30937_, _14712_, _07871_);
  or (_30938_, _30937_, _30933_);
  or (_30939_, _30938_, _06252_);
  and (_30941_, _07871_, \oc8051_golden_model_1.ACC [2]);
  or (_30942_, _30941_, _30933_);
  and (_30943_, _30942_, _07123_);
  and (_30944_, _07124_, \oc8051_golden_model_1.P3 [2]);
  or (_30945_, _30944_, _06251_);
  or (_30946_, _30945_, _30943_);
  and (_30947_, _30946_, _06476_);
  and (_30948_, _30947_, _30939_);
  and (_30949_, _13146_, \oc8051_golden_model_1.P3 [2]);
  and (_30950_, _14702_, _08539_);
  or (_30952_, _30950_, _30949_);
  and (_30953_, _30952_, _06475_);
  or (_30954_, _30953_, _06468_);
  or (_30955_, _30954_, _30948_);
  or (_30956_, _30935_, _07142_);
  and (_30957_, _30956_, _30955_);
  or (_30958_, _30957_, _06466_);
  or (_30959_, _30942_, _06801_);
  and (_30960_, _30959_, _06484_);
  and (_30961_, _30960_, _30958_);
  and (_30963_, _14706_, _08539_);
  or (_30964_, _30963_, _30949_);
  and (_30965_, _30964_, _06483_);
  or (_30966_, _30965_, _06461_);
  or (_30967_, _30966_, _30961_);
  or (_30968_, _30949_, _14739_);
  and (_30969_, _30968_, _30952_);
  or (_30970_, _30969_, _07164_);
  and (_30971_, _30970_, _06242_);
  and (_30972_, _30971_, _30967_);
  or (_30974_, _30949_, _14703_);
  and (_30975_, _30974_, _06241_);
  and (_30976_, _30975_, _30952_);
  or (_30977_, _30976_, _07187_);
  or (_30978_, _30977_, _30972_);
  and (_30979_, _30978_, _30936_);
  or (_30980_, _30979_, _07182_);
  and (_30981_, _09251_, _07871_);
  or (_30982_, _30933_, _07183_);
  or (_30983_, _30982_, _30981_);
  and (_30985_, _30983_, _06336_);
  and (_30986_, _30985_, _30980_);
  and (_30987_, _14808_, _07871_);
  or (_30988_, _30987_, _30933_);
  and (_30989_, _30988_, _05968_);
  or (_30990_, _30989_, _06371_);
  or (_30991_, _30990_, _30986_);
  and (_30992_, _07871_, _08945_);
  or (_30993_, _30992_, _30933_);
  or (_30994_, _30993_, _07198_);
  and (_30996_, _30994_, _30991_);
  or (_30997_, _30996_, _06367_);
  and (_30998_, _14824_, _07871_);
  or (_30999_, _30998_, _30933_);
  or (_31000_, _30999_, _07218_);
  and (_31001_, _31000_, _07216_);
  and (_31002_, _31001_, _30997_);
  and (_31003_, _11214_, _07871_);
  or (_31004_, _31003_, _30933_);
  and (_31005_, _31004_, _06533_);
  or (_31007_, _31005_, _31002_);
  and (_31008_, _31007_, _07213_);
  or (_31009_, _30933_, _08397_);
  and (_31010_, _30993_, _06366_);
  and (_31011_, _31010_, _31009_);
  or (_31012_, _31011_, _31008_);
  and (_31013_, _31012_, _07210_);
  and (_31014_, _30942_, _06541_);
  and (_31015_, _31014_, _31009_);
  or (_31016_, _31015_, _06383_);
  or (_31018_, _31016_, _31013_);
  and (_31019_, _14821_, _07871_);
  or (_31020_, _30933_, _07231_);
  or (_31021_, _31020_, _31019_);
  and (_31022_, _31021_, _07229_);
  and (_31023_, _31022_, _31018_);
  nor (_31024_, _11213_, _13138_);
  or (_31025_, _31024_, _30933_);
  and (_31026_, _31025_, _06528_);
  or (_31027_, _31026_, _06563_);
  or (_31030_, _31027_, _31023_);
  or (_31031_, _30938_, _07241_);
  and (_31032_, _31031_, _06571_);
  and (_31033_, _31032_, _31030_);
  and (_31034_, _30964_, _06199_);
  or (_31035_, _31034_, _06188_);
  or (_31036_, _31035_, _31033_);
  and (_31037_, _14884_, _07871_);
  or (_31038_, _30933_, _06189_);
  or (_31039_, _31038_, _31037_);
  and (_31041_, _31039_, _01452_);
  and (_31042_, _31041_, _31036_);
  nor (_31043_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_31044_, _31043_, _00000_);
  or (_43882_, _31044_, _31042_);
  nor (_31045_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_31046_, _31045_, _00000_);
  and (_31047_, _13138_, \oc8051_golden_model_1.P3 [3]);
  nor (_31048_, _13138_, _07713_);
  or (_31049_, _31048_, _31047_);
  or (_31052_, _31049_, _07188_);
  or (_31053_, _31049_, _07142_);
  and (_31054_, _14898_, _07871_);
  or (_31055_, _31054_, _31047_);
  or (_31056_, _31055_, _06252_);
  and (_31057_, _07871_, \oc8051_golden_model_1.ACC [3]);
  or (_31058_, _31057_, _31047_);
  and (_31059_, _31058_, _07123_);
  and (_31060_, _07124_, \oc8051_golden_model_1.P3 [3]);
  or (_31061_, _31060_, _06251_);
  or (_31063_, _31061_, _31059_);
  and (_31064_, _31063_, _06476_);
  and (_31065_, _31064_, _31056_);
  and (_31066_, _13146_, \oc8051_golden_model_1.P3 [3]);
  and (_31067_, _14906_, _08539_);
  or (_31068_, _31067_, _31066_);
  and (_31069_, _31068_, _06475_);
  or (_31070_, _31069_, _06468_);
  or (_31071_, _31070_, _31065_);
  and (_31072_, _31071_, _31053_);
  or (_31075_, _31072_, _06466_);
  or (_31076_, _31058_, _06801_);
  and (_31077_, _31076_, _06484_);
  and (_31078_, _31077_, _31075_);
  and (_31079_, _14904_, _08539_);
  or (_31080_, _31079_, _31066_);
  and (_31081_, _31080_, _06483_);
  or (_31082_, _31081_, _06461_);
  or (_31083_, _31082_, _31078_);
  or (_31084_, _31066_, _14931_);
  and (_31086_, _31084_, _31068_);
  or (_31087_, _31086_, _07164_);
  and (_31088_, _31087_, _06242_);
  and (_31089_, _31088_, _31083_);
  or (_31090_, _31066_, _14947_);
  and (_31091_, _31090_, _06241_);
  and (_31092_, _31091_, _31068_);
  or (_31093_, _31092_, _07187_);
  or (_31094_, _31093_, _31089_);
  and (_31095_, _31094_, _31052_);
  or (_31098_, _31095_, _07182_);
  and (_31099_, _09205_, _07871_);
  or (_31100_, _31047_, _07183_);
  or (_31101_, _31100_, _31099_);
  and (_31102_, _31101_, _06336_);
  and (_31103_, _31102_, _31098_);
  and (_31104_, _15003_, _07871_);
  or (_31105_, _31104_, _31047_);
  and (_31106_, _31105_, _05968_);
  or (_31107_, _31106_, _06371_);
  or (_31109_, _31107_, _31103_);
  and (_31110_, _07871_, _08872_);
  or (_31111_, _31110_, _31047_);
  or (_31112_, _31111_, _07198_);
  and (_31113_, _31112_, _31109_);
  or (_31114_, _31113_, _06367_);
  and (_31115_, _15018_, _07871_);
  or (_31116_, _31115_, _31047_);
  or (_31117_, _31116_, _07218_);
  and (_31118_, _31117_, _07216_);
  and (_31120_, _31118_, _31114_);
  and (_31121_, _12523_, _07871_);
  or (_31122_, _31121_, _31047_);
  and (_31123_, _31122_, _06533_);
  or (_31124_, _31123_, _31120_);
  and (_31125_, _31124_, _07213_);
  or (_31126_, _31047_, _08257_);
  and (_31127_, _31111_, _06366_);
  and (_31128_, _31127_, _31126_);
  or (_31129_, _31128_, _31125_);
  and (_31131_, _31129_, _07210_);
  and (_31132_, _31058_, _06541_);
  and (_31133_, _31132_, _31126_);
  or (_31134_, _31133_, _06383_);
  or (_31135_, _31134_, _31131_);
  and (_31136_, _15015_, _07871_);
  or (_31137_, _31047_, _07231_);
  or (_31138_, _31137_, _31136_);
  and (_31139_, _31138_, _07229_);
  and (_31140_, _31139_, _31135_);
  nor (_31141_, _11211_, _13138_);
  or (_31142_, _31141_, _31047_);
  and (_31143_, _31142_, _06528_);
  or (_31144_, _31143_, _06563_);
  or (_31145_, _31144_, _31140_);
  or (_31146_, _31055_, _07241_);
  and (_31147_, _31146_, _06571_);
  and (_31148_, _31147_, _31145_);
  and (_31149_, _31080_, _06199_);
  or (_31150_, _31149_, _06188_);
  or (_31153_, _31150_, _31148_);
  and (_31154_, _15075_, _07871_);
  or (_31155_, _31047_, _06189_);
  or (_31156_, _31155_, _31154_);
  and (_31157_, _31156_, _01452_);
  and (_31158_, _31157_, _31153_);
  or (_43883_, _31158_, _31046_);
  and (_31159_, _13138_, \oc8051_golden_model_1.P3 [4]);
  nor (_31160_, _08494_, _13138_);
  or (_31161_, _31160_, _31159_);
  or (_31162_, _31161_, _07188_);
  and (_31163_, _13146_, \oc8051_golden_model_1.P3 [4]);
  and (_31164_, _15089_, _08539_);
  or (_31165_, _31164_, _31163_);
  and (_31166_, _31165_, _06483_);
  or (_31167_, _31161_, _07142_);
  and (_31168_, _15108_, _07871_);
  or (_31169_, _31168_, _31159_);
  or (_31170_, _31169_, _06252_);
  and (_31171_, _07871_, \oc8051_golden_model_1.ACC [4]);
  or (_31174_, _31171_, _31159_);
  and (_31175_, _31174_, _07123_);
  and (_31176_, _07124_, \oc8051_golden_model_1.P3 [4]);
  or (_31177_, _31176_, _06251_);
  or (_31178_, _31177_, _31175_);
  and (_31179_, _31178_, _06476_);
  and (_31180_, _31179_, _31170_);
  and (_31181_, _15091_, _08539_);
  or (_31182_, _31181_, _31163_);
  and (_31183_, _31182_, _06475_);
  or (_31184_, _31183_, _06468_);
  or (_31185_, _31184_, _31180_);
  and (_31186_, _31185_, _31167_);
  or (_31187_, _31186_, _06466_);
  or (_31188_, _31174_, _06801_);
  and (_31189_, _31188_, _06484_);
  and (_31190_, _31189_, _31187_);
  or (_31191_, _31190_, _31166_);
  and (_31192_, _31191_, _07164_);
  and (_31193_, _15126_, _08539_);
  or (_31196_, _31193_, _31163_);
  and (_31197_, _31196_, _06461_);
  or (_31198_, _31197_, _31192_);
  and (_31199_, _31198_, _06242_);
  or (_31200_, _31163_, _15141_);
  and (_31201_, _31200_, _06241_);
  and (_31202_, _31201_, _31182_);
  or (_31203_, _31202_, _07187_);
  or (_31204_, _31203_, _31199_);
  and (_31205_, _31204_, _31162_);
  or (_31206_, _31205_, _07182_);
  and (_31207_, _09159_, _07871_);
  or (_31208_, _31159_, _07183_);
  or (_31209_, _31208_, _31207_);
  and (_31210_, _31209_, _06336_);
  and (_31211_, _31210_, _31206_);
  and (_31212_, _15198_, _07871_);
  or (_31213_, _31212_, _31159_);
  and (_31214_, _31213_, _05968_);
  or (_31215_, _31214_, _06371_);
  or (_31218_, _31215_, _31211_);
  and (_31219_, _08892_, _07871_);
  or (_31220_, _31219_, _31159_);
  or (_31221_, _31220_, _07198_);
  and (_31222_, _31221_, _31218_);
  or (_31223_, _31222_, _06367_);
  and (_31224_, _15214_, _07871_);
  or (_31225_, _31224_, _31159_);
  or (_31226_, _31225_, _07218_);
  and (_31227_, _31226_, _07216_);
  and (_31228_, _31227_, _31223_);
  and (_31229_, _11209_, _07871_);
  or (_31230_, _31229_, _31159_);
  and (_31231_, _31230_, _06533_);
  or (_31232_, _31231_, _31228_);
  and (_31233_, _31232_, _07213_);
  or (_31234_, _31159_, _08497_);
  and (_31235_, _31220_, _06366_);
  and (_31236_, _31235_, _31234_);
  or (_31237_, _31236_, _31233_);
  and (_31240_, _31237_, _07210_);
  and (_31241_, _31174_, _06541_);
  and (_31242_, _31241_, _31234_);
  or (_31243_, _31242_, _06383_);
  or (_31244_, _31243_, _31240_);
  and (_31245_, _15211_, _07871_);
  or (_31246_, _31159_, _07231_);
  or (_31247_, _31246_, _31245_);
  and (_31248_, _31247_, _07229_);
  and (_31249_, _31248_, _31244_);
  nor (_31250_, _11208_, _13138_);
  or (_31251_, _31250_, _31159_);
  and (_31252_, _31251_, _06528_);
  or (_31253_, _31252_, _06563_);
  or (_31254_, _31253_, _31249_);
  or (_31255_, _31169_, _07241_);
  and (_31256_, _31255_, _06571_);
  and (_31257_, _31256_, _31254_);
  and (_31258_, _31165_, _06199_);
  or (_31259_, _31258_, _06188_);
  or (_31262_, _31259_, _31257_);
  and (_31263_, _15280_, _07871_);
  or (_31264_, _31159_, _06189_);
  or (_31265_, _31264_, _31263_);
  and (_31266_, _31265_, _01452_);
  and (_31267_, _31266_, _31262_);
  nor (_31268_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_31269_, _31268_, _00000_);
  or (_43884_, _31269_, _31267_);
  nor (_31270_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_31271_, _31270_, _00000_);
  and (_31272_, _13138_, \oc8051_golden_model_1.P3 [5]);
  nor (_31273_, _08209_, _13138_);
  or (_31274_, _31273_, _31272_);
  or (_31275_, _31274_, _07142_);
  and (_31276_, _15311_, _07871_);
  or (_31277_, _31276_, _31272_);
  or (_31278_, _31277_, _06252_);
  and (_31279_, _07871_, \oc8051_golden_model_1.ACC [5]);
  or (_31280_, _31279_, _31272_);
  and (_31283_, _31280_, _07123_);
  and (_31284_, _07124_, \oc8051_golden_model_1.P3 [5]);
  or (_31285_, _31284_, _06251_);
  or (_31286_, _31285_, _31283_);
  and (_31287_, _31286_, _06476_);
  and (_31288_, _31287_, _31278_);
  and (_31289_, _13146_, \oc8051_golden_model_1.P3 [5]);
  and (_31290_, _15296_, _08539_);
  or (_31291_, _31290_, _31289_);
  and (_31292_, _31291_, _06475_);
  or (_31293_, _31292_, _06468_);
  or (_31294_, _31293_, _31288_);
  and (_31295_, _31294_, _31275_);
  or (_31296_, _31295_, _06466_);
  or (_31297_, _31280_, _06801_);
  and (_31298_, _31297_, _06484_);
  and (_31299_, _31298_, _31296_);
  and (_31300_, _15294_, _08539_);
  or (_31301_, _31300_, _31289_);
  and (_31302_, _31301_, _06483_);
  or (_31305_, _31302_, _06461_);
  or (_31306_, _31305_, _31299_);
  or (_31307_, _31289_, _15328_);
  and (_31308_, _31307_, _31291_);
  or (_31309_, _31308_, _07164_);
  and (_31310_, _31309_, _06242_);
  and (_31311_, _31310_, _31306_);
  or (_31312_, _31289_, _15344_);
  and (_31313_, _31312_, _06241_);
  and (_31314_, _31313_, _31291_);
  or (_31315_, _31314_, _07187_);
  or (_31316_, _31315_, _31311_);
  or (_31317_, _31274_, _07188_);
  and (_31318_, _31317_, _31316_);
  or (_31319_, _31318_, _07182_);
  and (_31320_, _09113_, _07871_);
  or (_31321_, _31272_, _07183_);
  or (_31322_, _31321_, _31320_);
  and (_31323_, _31322_, _06336_);
  and (_31324_, _31323_, _31319_);
  and (_31327_, _15400_, _07871_);
  or (_31328_, _31327_, _31272_);
  and (_31329_, _31328_, _05968_);
  or (_31330_, _31329_, _06371_);
  or (_31331_, _31330_, _31324_);
  and (_31332_, _08888_, _07871_);
  or (_31333_, _31332_, _31272_);
  or (_31334_, _31333_, _07198_);
  and (_31335_, _31334_, _31331_);
  or (_31336_, _31335_, _06367_);
  and (_31337_, _15416_, _07871_);
  or (_31338_, _31337_, _31272_);
  or (_31339_, _31338_, _07218_);
  and (_31340_, _31339_, _07216_);
  and (_31341_, _31340_, _31336_);
  and (_31342_, _11205_, _07871_);
  or (_31343_, _31342_, _31272_);
  and (_31344_, _31343_, _06533_);
  or (_31345_, _31344_, _31341_);
  and (_31346_, _31345_, _07213_);
  or (_31349_, _31272_, _08212_);
  and (_31350_, _31333_, _06366_);
  and (_31351_, _31350_, _31349_);
  or (_31352_, _31351_, _31346_);
  and (_31353_, _31352_, _07210_);
  and (_31354_, _31280_, _06541_);
  and (_31355_, _31354_, _31349_);
  or (_31356_, _31355_, _06383_);
  or (_31357_, _31356_, _31353_);
  and (_31358_, _15413_, _07871_);
  or (_31359_, _31272_, _07231_);
  or (_31360_, _31359_, _31358_);
  and (_31361_, _31360_, _07229_);
  and (_31362_, _31361_, _31357_);
  nor (_31363_, _11204_, _13138_);
  or (_31364_, _31363_, _31272_);
  and (_31365_, _31364_, _06528_);
  or (_31366_, _31365_, _06563_);
  or (_31367_, _31366_, _31362_);
  or (_31368_, _31277_, _07241_);
  and (_31371_, _31368_, _06571_);
  and (_31372_, _31371_, _31367_);
  and (_31373_, _31301_, _06199_);
  or (_31374_, _31373_, _06188_);
  or (_31375_, _31374_, _31372_);
  and (_31376_, _15477_, _07871_);
  or (_31377_, _31272_, _06189_);
  or (_31378_, _31377_, _31376_);
  and (_31379_, _31378_, _01452_);
  and (_31380_, _31379_, _31375_);
  or (_43885_, _31380_, _31271_);
  and (_31381_, _13138_, \oc8051_golden_model_1.P3 [6]);
  nor (_31382_, _08106_, _13138_);
  or (_31383_, _31382_, _31381_);
  or (_31384_, _31383_, _07142_);
  and (_31385_, _15512_, _07871_);
  or (_31386_, _31385_, _31381_);
  or (_31387_, _31386_, _06252_);
  and (_31388_, _07871_, \oc8051_golden_model_1.ACC [6]);
  or (_31389_, _31388_, _31381_);
  and (_31392_, _31389_, _07123_);
  and (_31393_, _07124_, \oc8051_golden_model_1.P3 [6]);
  or (_31394_, _31393_, _06251_);
  or (_31395_, _31394_, _31392_);
  and (_31396_, _31395_, _06476_);
  and (_31397_, _31396_, _31387_);
  and (_31398_, _13146_, \oc8051_golden_model_1.P3 [6]);
  and (_31399_, _15499_, _08539_);
  or (_31400_, _31399_, _31398_);
  and (_31401_, _31400_, _06475_);
  or (_31402_, _31401_, _06468_);
  or (_31403_, _31402_, _31397_);
  and (_31404_, _31403_, _31384_);
  or (_31405_, _31404_, _06466_);
  or (_31406_, _31389_, _06801_);
  and (_31407_, _31406_, _06484_);
  and (_31408_, _31407_, _31405_);
  and (_31409_, _15497_, _08539_);
  or (_31410_, _31409_, _31398_);
  and (_31411_, _31410_, _06483_);
  or (_31414_, _31411_, _06461_);
  or (_31415_, _31414_, _31408_);
  or (_31416_, _31398_, _15529_);
  and (_31417_, _31416_, _31400_);
  or (_31418_, _31417_, _07164_);
  and (_31419_, _31418_, _06242_);
  and (_31420_, _31419_, _31415_);
  or (_31421_, _31398_, _15545_);
  and (_31422_, _31421_, _06241_);
  and (_31423_, _31422_, _31400_);
  or (_31424_, _31423_, _07187_);
  or (_31425_, _31424_, _31420_);
  or (_31426_, _31383_, _07188_);
  and (_31427_, _31426_, _31425_);
  or (_31428_, _31427_, _07182_);
  and (_31429_, _09067_, _07871_);
  or (_31430_, _31381_, _07183_);
  or (_31431_, _31430_, _31429_);
  and (_31432_, _31431_, _06336_);
  and (_31433_, _31432_, _31428_);
  and (_31436_, _15601_, _07871_);
  or (_31437_, _31436_, _31381_);
  and (_31438_, _31437_, _05968_);
  or (_31439_, _31438_, _06371_);
  or (_31440_, _31439_, _31433_);
  and (_31441_, _15608_, _07871_);
  or (_31442_, _31441_, _31381_);
  or (_31443_, _31442_, _07198_);
  and (_31444_, _31443_, _31440_);
  or (_31445_, _31444_, _06367_);
  and (_31446_, _15618_, _07871_);
  or (_31447_, _31446_, _31381_);
  or (_31448_, _31447_, _07218_);
  and (_31449_, _31448_, _07216_);
  and (_31450_, _31449_, _31445_);
  and (_31451_, _11202_, _07871_);
  or (_31452_, _31451_, _31381_);
  and (_31453_, _31452_, _06533_);
  or (_31454_, _31453_, _31450_);
  and (_31455_, _31454_, _07213_);
  or (_31458_, _31381_, _08109_);
  and (_31459_, _31442_, _06366_);
  and (_31460_, _31459_, _31458_);
  or (_31461_, _31460_, _31455_);
  and (_31462_, _31461_, _07210_);
  and (_31463_, _31389_, _06541_);
  and (_31464_, _31463_, _31458_);
  or (_31465_, _31464_, _06383_);
  or (_31466_, _31465_, _31462_);
  and (_31467_, _15615_, _07871_);
  or (_31468_, _31381_, _07231_);
  or (_31469_, _31468_, _31467_);
  and (_31470_, _31469_, _07229_);
  and (_31471_, _31470_, _31466_);
  nor (_31472_, _11201_, _13138_);
  or (_31473_, _31472_, _31381_);
  and (_31474_, _31473_, _06528_);
  or (_31475_, _31474_, _06563_);
  or (_31476_, _31475_, _31471_);
  or (_31477_, _31386_, _07241_);
  and (_31480_, _31477_, _06571_);
  and (_31481_, _31480_, _31476_);
  and (_31482_, _31410_, _06199_);
  or (_31483_, _31482_, _06188_);
  or (_31484_, _31483_, _31481_);
  and (_31485_, _15676_, _07871_);
  or (_31486_, _31381_, _06189_);
  or (_31487_, _31486_, _31485_);
  and (_31488_, _31487_, _01452_);
  and (_31489_, _31488_, _31484_);
  nor (_31490_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_31491_, _31490_, _00000_);
  or (_43886_, _31491_, _31489_);
  nand (_31492_, _11218_, _07899_);
  not (_31493_, \oc8051_golden_model_1.P0 [0]);
  nor (_31494_, _07899_, _31493_);
  nor (_31495_, _31494_, _07210_);
  nand (_31496_, _31495_, _31492_);
  and (_31497_, _07899_, _07325_);
  or (_31498_, _31497_, _31494_);
  or (_31501_, _31498_, _07188_);
  nor (_31502_, _07920_, _31493_);
  and (_31503_, _14341_, _07920_);
  or (_31504_, _31503_, _31502_);
  and (_31505_, _31504_, _06475_);
  nor (_31506_, _08351_, _13241_);
  or (_31507_, _31506_, _31494_);
  or (_31508_, _31507_, _06252_);
  and (_31509_, _07899_, \oc8051_golden_model_1.ACC [0]);
  or (_31510_, _31509_, _31494_);
  and (_31511_, _31510_, _07123_);
  nor (_31512_, _07123_, _31493_);
  or (_31513_, _31512_, _06251_);
  or (_31514_, _31513_, _31511_);
  and (_31515_, _31514_, _06476_);
  and (_31516_, _31515_, _31508_);
  or (_31517_, _31516_, _31505_);
  and (_31518_, _31517_, _07142_);
  and (_31519_, _31498_, _06468_);
  or (_31520_, _31519_, _06466_);
  or (_31523_, _31520_, _31518_);
  or (_31524_, _31510_, _06801_);
  and (_31525_, _31524_, _06484_);
  and (_31526_, _31525_, _31523_);
  and (_31527_, _31494_, _06483_);
  or (_31528_, _31527_, _06461_);
  or (_31529_, _31528_, _31526_);
  or (_31530_, _31507_, _07164_);
  and (_31531_, _31530_, _06242_);
  and (_31532_, _31531_, _31529_);
  or (_31533_, _31502_, _14371_);
  and (_31534_, _31533_, _06241_);
  and (_31535_, _31534_, _31504_);
  or (_31536_, _31535_, _07187_);
  or (_31537_, _31536_, _31532_);
  and (_31538_, _31537_, _31501_);
  or (_31539_, _31538_, _07182_);
  and (_31540_, _09342_, _07899_);
  or (_31541_, _31494_, _07183_);
  or (_31542_, _31541_, _31540_);
  and (_31545_, _31542_, _31539_);
  or (_31546_, _31545_, _05968_);
  and (_31547_, _14427_, _07899_);
  or (_31548_, _31494_, _06336_);
  or (_31549_, _31548_, _31547_);
  and (_31550_, _31549_, _07198_);
  and (_31551_, _31550_, _31546_);
  and (_31552_, _07899_, _08908_);
  or (_31553_, _31552_, _31494_);
  and (_31554_, _31553_, _06371_);
  or (_31555_, _31554_, _06367_);
  or (_31556_, _31555_, _31551_);
  and (_31557_, _14442_, _07899_);
  or (_31558_, _31557_, _31494_);
  or (_31559_, _31558_, _07218_);
  and (_31560_, _31559_, _07216_);
  and (_31561_, _31560_, _31556_);
  nor (_31562_, _12526_, _13241_);
  or (_31563_, _31562_, _31494_);
  and (_31564_, _31492_, _06533_);
  and (_31567_, _31564_, _31563_);
  or (_31568_, _31567_, _31561_);
  and (_31569_, _31568_, _07213_);
  nand (_31570_, _31553_, _06366_);
  nor (_31571_, _31570_, _31506_);
  or (_31572_, _31571_, _06541_);
  or (_31573_, _31572_, _31569_);
  and (_31574_, _31573_, _31496_);
  or (_31575_, _31574_, _06383_);
  and (_31576_, _14325_, _07899_);
  or (_31577_, _31576_, _31494_);
  or (_31578_, _31577_, _07231_);
  and (_31579_, _31578_, _07229_);
  and (_31580_, _31579_, _31575_);
  and (_31581_, _31563_, _06528_);
  or (_31582_, _31581_, _06563_);
  or (_31583_, _31582_, _31580_);
  or (_31584_, _31507_, _07241_);
  and (_31585_, _31584_, _31583_);
  or (_31586_, _31585_, _06199_);
  or (_31589_, _31494_, _06571_);
  and (_31590_, _31589_, _31586_);
  or (_31591_, _31590_, _06188_);
  or (_31592_, _31507_, _06189_);
  and (_31593_, _31592_, _01452_);
  and (_31594_, _31593_, _31591_);
  nor (_31595_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_31596_, _31595_, _00000_);
  or (_43888_, _31596_, _31594_);
  nor (_31597_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_31598_, _31597_, _00000_);
  not (_31599_, \oc8051_golden_model_1.P0 [1]);
  nor (_31600_, _07899_, _31599_);
  nor (_31601_, _11216_, _13241_);
  or (_31602_, _31601_, _31600_);
  or (_31603_, _31602_, _07229_);
  nor (_31604_, _13241_, _07120_);
  or (_31605_, _31604_, _31600_);
  or (_31606_, _31605_, _07142_);
  or (_31607_, _07899_, \oc8051_golden_model_1.P0 [1]);
  and (_31610_, _14503_, _07899_);
  not (_31611_, _31610_);
  and (_31612_, _31611_, _31607_);
  or (_31613_, _31612_, _06252_);
  and (_31614_, _07899_, \oc8051_golden_model_1.ACC [1]);
  or (_31615_, _31614_, _31600_);
  and (_31616_, _31615_, _07123_);
  nor (_31617_, _07123_, _31599_);
  or (_31618_, _31617_, _06251_);
  or (_31619_, _31618_, _31616_);
  and (_31620_, _31619_, _06476_);
  and (_31621_, _31620_, _31613_);
  nor (_31622_, _07920_, _31599_);
  and (_31623_, _14510_, _07920_);
  or (_31624_, _31623_, _31622_);
  and (_31625_, _31624_, _06475_);
  or (_31626_, _31625_, _06468_);
  or (_31627_, _31626_, _31621_);
  and (_31628_, _31627_, _31606_);
  or (_31629_, _31628_, _06466_);
  or (_31632_, _31615_, _06801_);
  and (_31633_, _31632_, _06484_);
  and (_31634_, _31633_, _31629_);
  and (_31635_, _14513_, _07920_);
  or (_31636_, _31635_, _31622_);
  and (_31637_, _31636_, _06483_);
  or (_31638_, _31637_, _06461_);
  or (_31639_, _31638_, _31634_);
  or (_31640_, _31622_, _14509_);
  and (_31641_, _31640_, _31624_);
  or (_31642_, _31641_, _07164_);
  and (_31643_, _31642_, _06242_);
  and (_31644_, _31643_, _31639_);
  or (_31645_, _31622_, _14553_);
  and (_31646_, _31645_, _06241_);
  and (_31647_, _31646_, _31624_);
  or (_31648_, _31647_, _07187_);
  or (_31649_, _31648_, _31644_);
  or (_31650_, _31605_, _07188_);
  and (_31651_, _31650_, _31649_);
  or (_31654_, _31651_, _07182_);
  and (_31655_, _09297_, _07899_);
  or (_31656_, _31600_, _07183_);
  or (_31657_, _31656_, _31655_);
  and (_31658_, _31657_, _06336_);
  and (_31659_, _31658_, _31654_);
  and (_31660_, _14609_, _07899_);
  or (_31661_, _31660_, _31600_);
  and (_31662_, _31661_, _05968_);
  or (_31663_, _31662_, _31659_);
  and (_31664_, _31663_, _07198_);
  nand (_31665_, _07899_, _07018_);
  and (_31666_, _31607_, _06371_);
  and (_31667_, _31666_, _31665_);
  or (_31668_, _31667_, _31664_);
  and (_31669_, _31668_, _07218_);
  or (_31670_, _14625_, _13241_);
  and (_31671_, _31607_, _06367_);
  and (_31672_, _31671_, _31670_);
  or (_31673_, _31672_, _06533_);
  or (_31676_, _31673_, _31669_);
  nand (_31677_, _11215_, _07899_);
  and (_31678_, _31677_, _31602_);
  or (_31679_, _31678_, _07216_);
  and (_31680_, _31679_, _07213_);
  and (_31681_, _31680_, _31676_);
  or (_31682_, _14623_, _13241_);
  and (_31683_, _31607_, _06366_);
  and (_31684_, _31683_, _31682_);
  or (_31685_, _31684_, _06541_);
  or (_31686_, _31685_, _31681_);
  nor (_31687_, _31600_, _07210_);
  nand (_31688_, _31687_, _31677_);
  and (_31689_, _31688_, _07231_);
  and (_31690_, _31689_, _31686_);
  or (_31691_, _31665_, _08302_);
  and (_31692_, _31607_, _06383_);
  and (_31693_, _31692_, _31691_);
  or (_31694_, _31693_, _06528_);
  or (_31695_, _31694_, _31690_);
  and (_31698_, _31695_, _31603_);
  or (_31699_, _31698_, _06563_);
  or (_31700_, _31612_, _07241_);
  and (_31701_, _31700_, _06571_);
  and (_31702_, _31701_, _31699_);
  and (_31703_, _31636_, _06199_);
  or (_31704_, _31703_, _06188_);
  or (_31705_, _31704_, _31702_);
  or (_31706_, _31600_, _06189_);
  or (_31707_, _31706_, _31610_);
  and (_31708_, _31707_, _01452_);
  and (_31709_, _31708_, _31705_);
  or (_43889_, _31709_, _31598_);
  and (_31710_, _13241_, \oc8051_golden_model_1.P0 [2]);
  nor (_31711_, _13241_, _07578_);
  or (_31712_, _31711_, _31710_);
  or (_31713_, _31712_, _07188_);
  and (_31714_, _14712_, _07899_);
  or (_31715_, _31714_, _31710_);
  and (_31716_, _31715_, _06251_);
  and (_31719_, _07124_, \oc8051_golden_model_1.P0 [2]);
  and (_31720_, _07899_, \oc8051_golden_model_1.ACC [2]);
  or (_31721_, _31720_, _31710_);
  and (_31722_, _31721_, _07123_);
  or (_31723_, _31722_, _31719_);
  and (_31724_, _31723_, _06252_);
  or (_31725_, _31724_, _06475_);
  or (_31726_, _31725_, _31716_);
  and (_31727_, _13261_, \oc8051_golden_model_1.P0 [2]);
  and (_31728_, _14702_, _07920_);
  or (_31729_, _31728_, _31727_);
  or (_31730_, _31729_, _06476_);
  and (_31731_, _31730_, _31726_);
  or (_31732_, _31731_, _06468_);
  or (_31733_, _31712_, _07142_);
  and (_31734_, _31733_, _31732_);
  or (_31735_, _31734_, _06466_);
  or (_31736_, _31721_, _06801_);
  and (_31737_, _31736_, _06484_);
  and (_31738_, _31737_, _31735_);
  and (_31741_, _14706_, _07920_);
  or (_31742_, _31741_, _31727_);
  and (_31743_, _31742_, _06483_);
  or (_31744_, _31743_, _06461_);
  or (_31745_, _31744_, _31738_);
  or (_31746_, _31727_, _14739_);
  and (_31747_, _31746_, _31729_);
  or (_31748_, _31747_, _07164_);
  and (_31749_, _31748_, _06242_);
  and (_31750_, _31749_, _31745_);
  or (_31752_, _31727_, _14703_);
  and (_31753_, _31752_, _06241_);
  and (_31754_, _31753_, _31729_);
  or (_31755_, _31754_, _07187_);
  or (_31756_, _31755_, _31750_);
  and (_31757_, _31756_, _31713_);
  or (_31758_, _31757_, _07182_);
  and (_31759_, _09251_, _07899_);
  or (_31760_, _31710_, _07183_);
  or (_31761_, _31760_, _31759_);
  and (_31763_, _31761_, _06336_);
  and (_31764_, _31763_, _31758_);
  and (_31765_, _14808_, _07899_);
  or (_31766_, _31765_, _31710_);
  and (_31767_, _31766_, _05968_);
  or (_31768_, _31767_, _06371_);
  or (_31769_, _31768_, _31764_);
  and (_31770_, _07899_, _08945_);
  or (_31771_, _31770_, _31710_);
  or (_31772_, _31771_, _07198_);
  and (_31774_, _31772_, _31769_);
  or (_31775_, _31774_, _06367_);
  and (_31776_, _14824_, _07899_);
  or (_31777_, _31776_, _31710_);
  or (_31778_, _31777_, _07218_);
  and (_31779_, _31778_, _07216_);
  and (_31780_, _31779_, _31775_);
  and (_31781_, _11214_, _07899_);
  or (_31782_, _31781_, _31710_);
  and (_31783_, _31782_, _06533_);
  or (_31785_, _31783_, _31780_);
  and (_31786_, _31785_, _07213_);
  or (_31787_, _31710_, _08397_);
  and (_31788_, _31771_, _06366_);
  and (_31789_, _31788_, _31787_);
  or (_31790_, _31789_, _31786_);
  and (_31791_, _31790_, _07210_);
  and (_31792_, _31721_, _06541_);
  and (_31793_, _31792_, _31787_);
  or (_31794_, _31793_, _06383_);
  or (_31796_, _31794_, _31791_);
  and (_31797_, _14821_, _07899_);
  or (_31798_, _31710_, _07231_);
  or (_31799_, _31798_, _31797_);
  and (_31800_, _31799_, _07229_);
  and (_31801_, _31800_, _31796_);
  nor (_31802_, _11213_, _13241_);
  or (_31803_, _31802_, _31710_);
  and (_31804_, _31803_, _06528_);
  or (_31805_, _31804_, _06563_);
  or (_31807_, _31805_, _31801_);
  or (_31808_, _31715_, _07241_);
  and (_31809_, _31808_, _06571_);
  and (_31810_, _31809_, _31807_);
  and (_31811_, _31742_, _06199_);
  or (_31812_, _31811_, _06188_);
  or (_31813_, _31812_, _31810_);
  and (_31814_, _14884_, _07899_);
  or (_31815_, _31710_, _06189_);
  or (_31816_, _31815_, _31814_);
  and (_31818_, _31816_, _01452_);
  and (_31819_, _31818_, _31813_);
  nor (_31820_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_31821_, _31820_, _00000_);
  or (_43890_, _31821_, _31819_);
  and (_31822_, _13241_, \oc8051_golden_model_1.P0 [3]);
  nor (_31823_, _13241_, _07713_);
  or (_31824_, _31823_, _31822_);
  or (_31825_, _31824_, _07188_);
  or (_31826_, _31824_, _07142_);
  and (_31828_, _14898_, _07899_);
  or (_31829_, _31828_, _31822_);
  or (_31830_, _31829_, _06252_);
  and (_31831_, _07899_, \oc8051_golden_model_1.ACC [3]);
  or (_31832_, _31831_, _31822_);
  and (_31833_, _31832_, _07123_);
  and (_31834_, _07124_, \oc8051_golden_model_1.P0 [3]);
  or (_31835_, _31834_, _06251_);
  or (_31836_, _31835_, _31833_);
  and (_31837_, _31836_, _06476_);
  and (_31839_, _31837_, _31830_);
  and (_31840_, _13261_, \oc8051_golden_model_1.P0 [3]);
  and (_31841_, _14906_, _07920_);
  or (_31842_, _31841_, _31840_);
  and (_31843_, _31842_, _06475_);
  or (_31844_, _31843_, _06468_);
  or (_31845_, _31844_, _31839_);
  and (_31846_, _31845_, _31826_);
  or (_31847_, _31846_, _06466_);
  or (_31848_, _31832_, _06801_);
  and (_31850_, _31848_, _06484_);
  and (_31851_, _31850_, _31847_);
  and (_31852_, _14904_, _07920_);
  or (_31853_, _31852_, _31840_);
  and (_31854_, _31853_, _06483_);
  or (_31855_, _31854_, _06461_);
  or (_31856_, _31855_, _31851_);
  or (_31857_, _31840_, _14931_);
  and (_31858_, _31857_, _31842_);
  or (_31859_, _31858_, _07164_);
  and (_31861_, _31859_, _06242_);
  and (_31862_, _31861_, _31856_);
  or (_31863_, _31840_, _14947_);
  and (_31864_, _31863_, _06241_);
  and (_31865_, _31864_, _31842_);
  or (_31866_, _31865_, _07187_);
  or (_31867_, _31866_, _31862_);
  and (_31868_, _31867_, _31825_);
  or (_31869_, _31868_, _07182_);
  and (_31870_, _09205_, _07899_);
  or (_31872_, _31822_, _07183_);
  or (_31873_, _31872_, _31870_);
  and (_31874_, _31873_, _06336_);
  and (_31875_, _31874_, _31869_);
  and (_31876_, _15003_, _07899_);
  or (_31877_, _31876_, _31822_);
  and (_31878_, _31877_, _05968_);
  or (_31879_, _31878_, _06371_);
  or (_31880_, _31879_, _31875_);
  and (_31881_, _07899_, _08872_);
  or (_31883_, _31881_, _31822_);
  or (_31884_, _31883_, _07198_);
  and (_31885_, _31884_, _31880_);
  or (_31886_, _31885_, _06367_);
  and (_31887_, _15018_, _07899_);
  or (_31888_, _31887_, _31822_);
  or (_31889_, _31888_, _07218_);
  and (_31890_, _31889_, _07216_);
  and (_31891_, _31890_, _31886_);
  and (_31892_, _12523_, _07899_);
  or (_31894_, _31892_, _31822_);
  and (_31895_, _31894_, _06533_);
  or (_31896_, _31895_, _31891_);
  and (_31897_, _31896_, _07213_);
  or (_31898_, _31822_, _08257_);
  and (_31899_, _31883_, _06366_);
  and (_31900_, _31899_, _31898_);
  or (_31901_, _31900_, _31897_);
  and (_31902_, _31901_, _07210_);
  and (_31903_, _31832_, _06541_);
  and (_31905_, _31903_, _31898_);
  or (_31906_, _31905_, _06383_);
  or (_31907_, _31906_, _31902_);
  and (_31908_, _15015_, _07899_);
  or (_31909_, _31822_, _07231_);
  or (_31910_, _31909_, _31908_);
  and (_31911_, _31910_, _07229_);
  and (_31912_, _31911_, _31907_);
  nor (_31913_, _11211_, _13241_);
  or (_31914_, _31913_, _31822_);
  and (_31916_, _31914_, _06528_);
  or (_31917_, _31916_, _06563_);
  or (_31918_, _31917_, _31912_);
  or (_31919_, _31829_, _07241_);
  and (_31920_, _31919_, _06571_);
  and (_31921_, _31920_, _31918_);
  and (_31922_, _31853_, _06199_);
  or (_31923_, _31922_, _06188_);
  or (_31924_, _31923_, _31921_);
  and (_31925_, _15075_, _07899_);
  or (_31927_, _31822_, _06189_);
  or (_31928_, _31927_, _31925_);
  and (_31929_, _31928_, _01452_);
  and (_31930_, _31929_, _31924_);
  nor (_31931_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_31932_, _31931_, _00000_);
  or (_43892_, _31932_, _31930_);
  nor (_31933_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_31934_, _31933_, _00000_);
  and (_31935_, _13241_, \oc8051_golden_model_1.P0 [4]);
  nor (_31937_, _08494_, _13241_);
  or (_31938_, _31937_, _31935_);
  or (_31939_, _31938_, _07188_);
  and (_31940_, _13261_, \oc8051_golden_model_1.P0 [4]);
  and (_31941_, _15089_, _07920_);
  or (_31942_, _31941_, _31940_);
  and (_31943_, _31942_, _06483_);
  or (_31944_, _31938_, _07142_);
  and (_31945_, _15108_, _07899_);
  or (_31946_, _31945_, _31935_);
  or (_31948_, _31946_, _06252_);
  and (_31949_, _07899_, \oc8051_golden_model_1.ACC [4]);
  or (_31950_, _31949_, _31935_);
  and (_31951_, _31950_, _07123_);
  and (_31952_, _07124_, \oc8051_golden_model_1.P0 [4]);
  or (_31953_, _31952_, _06251_);
  or (_31954_, _31953_, _31951_);
  and (_31955_, _31954_, _06476_);
  and (_31956_, _31955_, _31948_);
  and (_31957_, _15091_, _07920_);
  or (_31959_, _31957_, _31940_);
  and (_31960_, _31959_, _06475_);
  or (_31961_, _31960_, _06468_);
  or (_31962_, _31961_, _31956_);
  and (_31963_, _31962_, _31944_);
  or (_31964_, _31963_, _06466_);
  or (_31965_, _31950_, _06801_);
  and (_31966_, _31965_, _06484_);
  and (_31967_, _31966_, _31964_);
  or (_31968_, _31967_, _31943_);
  and (_31970_, _31968_, _07164_);
  and (_31971_, _15126_, _07920_);
  or (_31972_, _31971_, _31940_);
  and (_31973_, _31972_, _06461_);
  or (_31974_, _31973_, _31970_);
  and (_31975_, _31974_, _06242_);
  or (_31976_, _31940_, _15141_);
  and (_31977_, _31976_, _06241_);
  and (_31978_, _31977_, _31959_);
  or (_31979_, _31978_, _07187_);
  or (_31980_, _31979_, _31975_);
  and (_31981_, _31980_, _31939_);
  or (_31982_, _31981_, _07182_);
  and (_31983_, _09159_, _07899_);
  or (_31984_, _31935_, _07183_);
  or (_31985_, _31984_, _31983_);
  and (_31986_, _31985_, _06336_);
  and (_31987_, _31986_, _31982_);
  and (_31988_, _15198_, _07899_);
  or (_31989_, _31988_, _31935_);
  and (_31991_, _31989_, _05968_);
  or (_31992_, _31991_, _06371_);
  or (_31993_, _31992_, _31987_);
  and (_31994_, _08892_, _07899_);
  or (_31995_, _31994_, _31935_);
  or (_31996_, _31995_, _07198_);
  and (_31997_, _31996_, _31993_);
  or (_31998_, _31997_, _06367_);
  and (_31999_, _15214_, _07899_);
  or (_32000_, _31999_, _31935_);
  or (_32002_, _32000_, _07218_);
  and (_32003_, _32002_, _07216_);
  and (_32004_, _32003_, _31998_);
  and (_32005_, _11209_, _07899_);
  or (_32006_, _32005_, _31935_);
  and (_32007_, _32006_, _06533_);
  or (_32008_, _32007_, _32004_);
  and (_32009_, _32008_, _07213_);
  or (_32010_, _31935_, _08497_);
  and (_32011_, _31995_, _06366_);
  and (_32013_, _32011_, _32010_);
  or (_32014_, _32013_, _32009_);
  and (_32015_, _32014_, _07210_);
  and (_32016_, _31950_, _06541_);
  and (_32017_, _32016_, _32010_);
  or (_32018_, _32017_, _06383_);
  or (_32019_, _32018_, _32015_);
  and (_32020_, _15211_, _07899_);
  or (_32021_, _31935_, _07231_);
  or (_32022_, _32021_, _32020_);
  and (_32024_, _32022_, _07229_);
  and (_32025_, _32024_, _32019_);
  nor (_32026_, _11208_, _13241_);
  or (_32027_, _32026_, _31935_);
  and (_32028_, _32027_, _06528_);
  or (_32029_, _32028_, _06563_);
  or (_32030_, _32029_, _32025_);
  or (_32031_, _31946_, _07241_);
  and (_32032_, _32031_, _06571_);
  and (_32033_, _32032_, _32030_);
  and (_32035_, _31942_, _06199_);
  or (_32036_, _32035_, _06188_);
  or (_32037_, _32036_, _32033_);
  and (_32038_, _15280_, _07899_);
  or (_32039_, _31935_, _06189_);
  or (_32040_, _32039_, _32038_);
  and (_32041_, _32040_, _01452_);
  and (_32042_, _32041_, _32037_);
  or (_43893_, _32042_, _31934_);
  and (_32043_, _13241_, \oc8051_golden_model_1.P0 [5]);
  nor (_32045_, _08209_, _13241_);
  or (_32046_, _32045_, _32043_);
  or (_32047_, _32046_, _07142_);
  and (_32048_, _15311_, _07899_);
  or (_32049_, _32048_, _32043_);
  or (_32050_, _32049_, _06252_);
  and (_32051_, _07899_, \oc8051_golden_model_1.ACC [5]);
  or (_32052_, _32051_, _32043_);
  and (_32053_, _32052_, _07123_);
  and (_32054_, _07124_, \oc8051_golden_model_1.P0 [5]);
  or (_32056_, _32054_, _06251_);
  or (_32057_, _32056_, _32053_);
  and (_32058_, _32057_, _06476_);
  and (_32059_, _32058_, _32050_);
  and (_32060_, _13261_, \oc8051_golden_model_1.P0 [5]);
  and (_32061_, _15296_, _07920_);
  or (_32062_, _32061_, _32060_);
  and (_32063_, _32062_, _06475_);
  or (_32064_, _32063_, _06468_);
  or (_32065_, _32064_, _32059_);
  and (_32067_, _32065_, _32047_);
  or (_32068_, _32067_, _06466_);
  or (_32069_, _32052_, _06801_);
  and (_32070_, _32069_, _06484_);
  and (_32071_, _32070_, _32068_);
  and (_32072_, _15294_, _07920_);
  or (_32073_, _32072_, _32060_);
  and (_32074_, _32073_, _06483_);
  or (_32075_, _32074_, _06461_);
  or (_32076_, _32075_, _32071_);
  or (_32078_, _32060_, _15328_);
  and (_32079_, _32078_, _32062_);
  or (_32080_, _32079_, _07164_);
  and (_32081_, _32080_, _06242_);
  and (_32082_, _32081_, _32076_);
  or (_32083_, _32060_, _15344_);
  and (_32084_, _32083_, _06241_);
  and (_32085_, _32084_, _32062_);
  or (_32086_, _32085_, _07187_);
  or (_32087_, _32086_, _32082_);
  or (_32089_, _32046_, _07188_);
  and (_32090_, _32089_, _32087_);
  or (_32091_, _32090_, _07182_);
  and (_32092_, _09113_, _07899_);
  or (_32093_, _32043_, _07183_);
  or (_32094_, _32093_, _32092_);
  and (_32095_, _32094_, _06336_);
  and (_32096_, _32095_, _32091_);
  and (_32097_, _15400_, _07899_);
  or (_32098_, _32097_, _32043_);
  and (_32100_, _32098_, _05968_);
  or (_32101_, _32100_, _06371_);
  or (_32102_, _32101_, _32096_);
  and (_32103_, _08888_, _07899_);
  or (_32104_, _32103_, _32043_);
  or (_32105_, _32104_, _07198_);
  and (_32106_, _32105_, _32102_);
  or (_32107_, _32106_, _06367_);
  and (_32108_, _15416_, _07899_);
  or (_32109_, _32108_, _32043_);
  or (_32111_, _32109_, _07218_);
  and (_32112_, _32111_, _07216_);
  and (_32113_, _32112_, _32107_);
  and (_32114_, _11205_, _07899_);
  or (_32115_, _32114_, _32043_);
  and (_32116_, _32115_, _06533_);
  or (_32117_, _32116_, _32113_);
  and (_32118_, _32117_, _07213_);
  or (_32119_, _32043_, _08212_);
  and (_32120_, _32104_, _06366_);
  and (_32122_, _32120_, _32119_);
  or (_32123_, _32122_, _32118_);
  and (_32124_, _32123_, _07210_);
  and (_32125_, _32052_, _06541_);
  and (_32126_, _32125_, _32119_);
  or (_32127_, _32126_, _06383_);
  or (_32128_, _32127_, _32124_);
  and (_32129_, _15413_, _07899_);
  or (_32130_, _32043_, _07231_);
  or (_32131_, _32130_, _32129_);
  and (_32133_, _32131_, _07229_);
  and (_32134_, _32133_, _32128_);
  nor (_32135_, _11204_, _13241_);
  or (_32136_, _32135_, _32043_);
  and (_32137_, _32136_, _06528_);
  or (_32138_, _32137_, _06563_);
  or (_32139_, _32138_, _32134_);
  or (_32140_, _32049_, _07241_);
  and (_32141_, _32140_, _06571_);
  and (_32142_, _32141_, _32139_);
  and (_32144_, _32073_, _06199_);
  or (_32145_, _32144_, _06188_);
  or (_32146_, _32145_, _32142_);
  and (_32147_, _15477_, _07899_);
  or (_32148_, _32043_, _06189_);
  or (_32149_, _32148_, _32147_);
  and (_32150_, _32149_, _01452_);
  and (_32151_, _32150_, _32146_);
  nor (_32152_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_32153_, _32152_, _00000_);
  or (_43894_, _32153_, _32151_);
  and (_32155_, _13241_, \oc8051_golden_model_1.P0 [6]);
  nor (_32156_, _08106_, _13241_);
  or (_32157_, _32156_, _32155_);
  or (_32158_, _32157_, _07142_);
  and (_32159_, _15512_, _07899_);
  or (_32160_, _32159_, _32155_);
  or (_32161_, _32160_, _06252_);
  and (_32162_, _07899_, \oc8051_golden_model_1.ACC [6]);
  or (_32163_, _32162_, _32155_);
  and (_32165_, _32163_, _07123_);
  and (_32166_, _07124_, \oc8051_golden_model_1.P0 [6]);
  or (_32167_, _32166_, _06251_);
  or (_32168_, _32167_, _32165_);
  and (_32169_, _32168_, _06476_);
  and (_32170_, _32169_, _32161_);
  and (_32171_, _13261_, \oc8051_golden_model_1.P0 [6]);
  and (_32172_, _15499_, _07920_);
  or (_32173_, _32172_, _32171_);
  and (_32174_, _32173_, _06475_);
  or (_32176_, _32174_, _06468_);
  or (_32177_, _32176_, _32170_);
  and (_32178_, _32177_, _32158_);
  or (_32179_, _32178_, _06466_);
  or (_32180_, _32163_, _06801_);
  and (_32181_, _32180_, _06484_);
  and (_32182_, _32181_, _32179_);
  and (_32183_, _15497_, _07920_);
  or (_32184_, _32183_, _32171_);
  and (_32185_, _32184_, _06483_);
  or (_32187_, _32185_, _06461_);
  or (_32188_, _32187_, _32182_);
  or (_32189_, _32171_, _15529_);
  and (_32190_, _32189_, _32173_);
  or (_32191_, _32190_, _07164_);
  and (_32192_, _32191_, _06242_);
  and (_32193_, _32192_, _32188_);
  or (_32194_, _32171_, _15545_);
  and (_32195_, _32194_, _06241_);
  and (_32196_, _32195_, _32173_);
  or (_32198_, _32196_, _07187_);
  or (_32199_, _32198_, _32193_);
  or (_32200_, _32157_, _07188_);
  and (_32201_, _32200_, _32199_);
  or (_32202_, _32201_, _07182_);
  and (_32203_, _09067_, _07899_);
  or (_32204_, _32155_, _07183_);
  or (_32205_, _32204_, _32203_);
  and (_32206_, _32205_, _06336_);
  and (_32207_, _32206_, _32202_);
  and (_32209_, _15601_, _07899_);
  or (_32210_, _32209_, _32155_);
  and (_32211_, _32210_, _05968_);
  or (_32212_, _32211_, _06371_);
  or (_32213_, _32212_, _32207_);
  and (_32214_, _15608_, _07899_);
  or (_32215_, _32214_, _32155_);
  or (_32216_, _32215_, _07198_);
  and (_32217_, _32216_, _32213_);
  or (_32218_, _32217_, _06367_);
  and (_32220_, _15618_, _07899_);
  or (_32221_, _32220_, _32155_);
  or (_32222_, _32221_, _07218_);
  and (_32223_, _32222_, _07216_);
  and (_32224_, _32223_, _32218_);
  and (_32225_, _11202_, _07899_);
  or (_32226_, _32225_, _32155_);
  and (_32227_, _32226_, _06533_);
  or (_32228_, _32227_, _32224_);
  and (_32229_, _32228_, _07213_);
  or (_32231_, _32155_, _08109_);
  and (_32232_, _32215_, _06366_);
  and (_32233_, _32232_, _32231_);
  or (_32234_, _32233_, _32229_);
  and (_32235_, _32234_, _07210_);
  and (_32236_, _32163_, _06541_);
  and (_32237_, _32236_, _32231_);
  or (_32238_, _32237_, _06383_);
  or (_32239_, _32238_, _32235_);
  and (_32240_, _15615_, _07899_);
  or (_32242_, _32155_, _07231_);
  or (_32243_, _32242_, _32240_);
  and (_32244_, _32243_, _07229_);
  and (_32245_, _32244_, _32239_);
  nor (_32246_, _11201_, _13241_);
  or (_32247_, _32246_, _32155_);
  and (_32248_, _32247_, _06528_);
  or (_32249_, _32248_, _06563_);
  or (_32250_, _32249_, _32245_);
  or (_32251_, _32160_, _07241_);
  and (_32253_, _32251_, _06571_);
  and (_32254_, _32253_, _32250_);
  and (_32255_, _32184_, _06199_);
  or (_32256_, _32255_, _06188_);
  or (_32257_, _32256_, _32254_);
  and (_32258_, _15676_, _07899_);
  or (_32259_, _32155_, _06189_);
  or (_32260_, _32259_, _32258_);
  and (_32261_, _32260_, _01452_);
  and (_32262_, _32261_, _32257_);
  nor (_32264_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_32265_, _32264_, _00000_);
  or (_43895_, _32265_, _32262_);
  nor (_32266_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_32267_, _32266_, _00000_);
  nand (_32268_, _11218_, _07945_);
  and (_32269_, _13346_, \oc8051_golden_model_1.P1 [0]);
  nor (_32270_, _32269_, _07210_);
  nand (_32271_, _32270_, _32268_);
  and (_32272_, _07945_, _07325_);
  or (_32274_, _32272_, _32269_);
  or (_32275_, _32274_, _07188_);
  and (_32276_, _13366_, \oc8051_golden_model_1.P1 [0]);
  and (_32277_, _14341_, _08531_);
  or (_32278_, _32277_, _32276_);
  and (_32279_, _32278_, _06475_);
  nor (_32280_, _08351_, _13346_);
  or (_32281_, _32280_, _32269_);
  or (_32282_, _32281_, _06252_);
  and (_32283_, _07945_, \oc8051_golden_model_1.ACC [0]);
  or (_32285_, _32283_, _32269_);
  and (_32286_, _32285_, _07123_);
  and (_32287_, _07124_, \oc8051_golden_model_1.P1 [0]);
  or (_32288_, _32287_, _06251_);
  or (_32289_, _32288_, _32286_);
  and (_32290_, _32289_, _06476_);
  and (_32291_, _32290_, _32282_);
  or (_32292_, _32291_, _32279_);
  and (_32293_, _32292_, _07142_);
  and (_32294_, _32274_, _06468_);
  or (_32296_, _32294_, _06466_);
  or (_32297_, _32296_, _32293_);
  or (_32298_, _32285_, _06801_);
  and (_32299_, _32298_, _06484_);
  and (_32300_, _32299_, _32297_);
  and (_32301_, _32269_, _06483_);
  or (_32302_, _32301_, _06461_);
  or (_32303_, _32302_, _32300_);
  or (_32304_, _32281_, _07164_);
  and (_32305_, _32304_, _06242_);
  and (_32307_, _32305_, _32303_);
  or (_32308_, _32276_, _14371_);
  and (_32309_, _32308_, _06241_);
  and (_32310_, _32309_, _32278_);
  or (_32311_, _32310_, _07187_);
  or (_32312_, _32311_, _32307_);
  and (_32313_, _32312_, _32275_);
  or (_32314_, _32313_, _07182_);
  and (_32315_, _09342_, _07945_);
  or (_32316_, _32269_, _07183_);
  or (_32318_, _32316_, _32315_);
  and (_32319_, _32318_, _32314_);
  or (_32320_, _32319_, _05968_);
  and (_32321_, _14427_, _07945_);
  or (_32322_, _32269_, _06336_);
  or (_32323_, _32322_, _32321_);
  and (_32324_, _32323_, _07198_);
  and (_32325_, _32324_, _32320_);
  and (_32326_, _07945_, _08908_);
  or (_32327_, _32326_, _32269_);
  and (_32329_, _32327_, _06371_);
  or (_32330_, _32329_, _06367_);
  or (_32331_, _32330_, _32325_);
  and (_32332_, _14442_, _07945_);
  or (_32333_, _32332_, _32269_);
  or (_32334_, _32333_, _07218_);
  and (_32335_, _32334_, _07216_);
  and (_32336_, _32335_, _32331_);
  nor (_32337_, _12526_, _13346_);
  or (_32338_, _32337_, _32269_);
  and (_32340_, _32268_, _06533_);
  and (_32341_, _32340_, _32338_);
  or (_32342_, _32341_, _32336_);
  and (_32343_, _32342_, _07213_);
  nand (_32344_, _32327_, _06366_);
  nor (_32345_, _32344_, _32280_);
  or (_32346_, _32345_, _06541_);
  or (_32347_, _32346_, _32343_);
  and (_32348_, _32347_, _32271_);
  or (_32349_, _32348_, _06383_);
  and (_32351_, _14325_, _07945_);
  or (_32352_, _32269_, _07231_);
  or (_32353_, _32352_, _32351_);
  and (_32354_, _32353_, _07229_);
  and (_32355_, _32354_, _32349_);
  and (_32356_, _32338_, _06528_);
  or (_32357_, _32356_, _06563_);
  or (_32358_, _32357_, _32355_);
  or (_32359_, _32281_, _07241_);
  and (_32360_, _32359_, _32358_);
  or (_32362_, _32360_, _06199_);
  or (_32363_, _32269_, _06571_);
  and (_32364_, _32363_, _32362_);
  or (_32365_, _32364_, _06188_);
  or (_32366_, _32281_, _06189_);
  and (_32367_, _32366_, _01452_);
  and (_32368_, _32367_, _32365_);
  or (_43897_, _32368_, _32267_);
  nor (_32369_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_32370_, _32369_, _00000_);
  and (_32372_, _13346_, \oc8051_golden_model_1.P1 [1]);
  nor (_32373_, _11216_, _13346_);
  or (_32374_, _32373_, _32372_);
  or (_32375_, _32374_, _07229_);
  nand (_32376_, _07945_, _07018_);
  or (_32377_, _07945_, \oc8051_golden_model_1.P1 [1]);
  and (_32378_, _32377_, _06371_);
  and (_32379_, _32378_, _32376_);
  nor (_32380_, _13346_, _07120_);
  or (_32381_, _32380_, _32372_);
  or (_32383_, _32381_, _07142_);
  and (_32384_, _14503_, _07945_);
  not (_32385_, _32384_);
  and (_32386_, _32385_, _32377_);
  or (_32387_, _32386_, _06252_);
  and (_32388_, _07945_, \oc8051_golden_model_1.ACC [1]);
  or (_32389_, _32388_, _32372_);
  and (_32390_, _32389_, _07123_);
  and (_32391_, _07124_, \oc8051_golden_model_1.P1 [1]);
  or (_32392_, _32391_, _06251_);
  or (_32394_, _32392_, _32390_);
  and (_32395_, _32394_, _06476_);
  and (_32396_, _32395_, _32387_);
  and (_32397_, _13366_, \oc8051_golden_model_1.P1 [1]);
  and (_32398_, _14510_, _08531_);
  or (_32399_, _32398_, _32397_);
  and (_32400_, _32399_, _06475_);
  or (_32401_, _32400_, _06468_);
  or (_32402_, _32401_, _32396_);
  and (_32403_, _32402_, _32383_);
  or (_32405_, _32403_, _06466_);
  or (_32406_, _32389_, _06801_);
  and (_32407_, _32406_, _06484_);
  and (_32408_, _32407_, _32405_);
  and (_32409_, _14513_, _08531_);
  or (_32410_, _32409_, _32397_);
  and (_32411_, _32410_, _06483_);
  or (_32412_, _32411_, _06461_);
  or (_32413_, _32412_, _32408_);
  or (_32414_, _32397_, _14509_);
  and (_32416_, _32414_, _32399_);
  or (_32417_, _32416_, _07164_);
  and (_32418_, _32417_, _06242_);
  and (_32419_, _32418_, _32413_);
  or (_32420_, _32397_, _14553_);
  and (_32421_, _32420_, _06241_);
  and (_32422_, _32421_, _32399_);
  or (_32423_, _32422_, _07187_);
  or (_32424_, _32423_, _32419_);
  or (_32425_, _32381_, _07188_);
  and (_32427_, _32425_, _32424_);
  or (_32428_, _32427_, _07182_);
  and (_32429_, _09297_, _07945_);
  or (_32430_, _32372_, _07183_);
  or (_32431_, _32430_, _32429_);
  and (_32432_, _32431_, _06336_);
  and (_32433_, _32432_, _32428_);
  and (_32434_, _14609_, _07945_);
  or (_32435_, _32434_, _32372_);
  and (_32436_, _32435_, _05968_);
  or (_32438_, _32436_, _32433_);
  and (_32439_, _32438_, _07198_);
  or (_32440_, _32439_, _32379_);
  and (_32441_, _32440_, _07218_);
  or (_32442_, _14625_, _13346_);
  and (_32443_, _32377_, _06367_);
  and (_32444_, _32443_, _32442_);
  or (_32445_, _32444_, _06533_);
  or (_32446_, _32445_, _32441_);
  and (_32447_, _11217_, _07945_);
  or (_32449_, _32447_, _32372_);
  or (_32450_, _32449_, _07216_);
  and (_32451_, _32450_, _07213_);
  and (_32452_, _32451_, _32446_);
  or (_32453_, _14623_, _13346_);
  and (_32454_, _32377_, _06366_);
  and (_32455_, _32454_, _32453_);
  or (_32456_, _32455_, _06541_);
  or (_32457_, _32456_, _32452_);
  and (_32458_, _32388_, _08302_);
  or (_32460_, _32372_, _07210_);
  or (_32461_, _32460_, _32458_);
  and (_32462_, _32461_, _07231_);
  and (_32463_, _32462_, _32457_);
  or (_32464_, _32376_, _08302_);
  and (_32465_, _32377_, _06383_);
  and (_32466_, _32465_, _32464_);
  or (_32467_, _32466_, _06528_);
  or (_32468_, _32467_, _32463_);
  and (_32469_, _32468_, _32375_);
  or (_32471_, _32469_, _06563_);
  or (_32472_, _32386_, _07241_);
  and (_32473_, _32472_, _06571_);
  and (_32474_, _32473_, _32471_);
  and (_32475_, _32410_, _06199_);
  or (_32476_, _32475_, _06188_);
  or (_32477_, _32476_, _32474_);
  or (_32478_, _32372_, _06189_);
  or (_32479_, _32478_, _32384_);
  and (_32480_, _32479_, _01452_);
  and (_32482_, _32480_, _32477_);
  or (_43898_, _32482_, _32370_);
  nor (_32483_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_32484_, _32483_, _00000_);
  and (_32485_, _13346_, \oc8051_golden_model_1.P1 [2]);
  nor (_32486_, _13346_, _07578_);
  or (_32487_, _32486_, _32485_);
  or (_32488_, _32487_, _07188_);
  and (_32489_, _14712_, _07945_);
  or (_32490_, _32489_, _32485_);
  or (_32492_, _32490_, _06252_);
  and (_32493_, _07945_, \oc8051_golden_model_1.ACC [2]);
  or (_32494_, _32493_, _32485_);
  and (_32495_, _32494_, _07123_);
  and (_32496_, _07124_, \oc8051_golden_model_1.P1 [2]);
  or (_32497_, _32496_, _06251_);
  or (_32498_, _32497_, _32495_);
  and (_32499_, _32498_, _06476_);
  and (_32500_, _32499_, _32492_);
  and (_32501_, _13366_, \oc8051_golden_model_1.P1 [2]);
  and (_32503_, _14702_, _08531_);
  or (_32504_, _32503_, _32501_);
  and (_32505_, _32504_, _06475_);
  or (_32506_, _32505_, _06468_);
  or (_32507_, _32506_, _32500_);
  or (_32508_, _32487_, _07142_);
  and (_32509_, _32508_, _32507_);
  or (_32510_, _32509_, _06466_);
  or (_32511_, _32494_, _06801_);
  and (_32512_, _32511_, _06484_);
  and (_32514_, _32512_, _32510_);
  and (_32515_, _14706_, _08531_);
  or (_32516_, _32515_, _32501_);
  and (_32517_, _32516_, _06483_);
  or (_32518_, _32517_, _06461_);
  or (_32519_, _32518_, _32514_);
  or (_32520_, _32501_, _14739_);
  and (_32521_, _32520_, _32504_);
  or (_32522_, _32521_, _07164_);
  and (_32523_, _32522_, _06242_);
  and (_32525_, _32523_, _32519_);
  or (_32526_, _32501_, _14703_);
  and (_32527_, _32526_, _06241_);
  and (_32528_, _32527_, _32504_);
  or (_32529_, _32528_, _07187_);
  or (_32530_, _32529_, _32525_);
  and (_32531_, _32530_, _32488_);
  or (_32532_, _32531_, _07182_);
  and (_32533_, _09251_, _07945_);
  or (_32534_, _32485_, _07183_);
  or (_32536_, _32534_, _32533_);
  and (_32537_, _32536_, _06336_);
  and (_32538_, _32537_, _32532_);
  and (_32539_, _14808_, _07945_);
  or (_32540_, _32539_, _32485_);
  and (_32541_, _32540_, _05968_);
  or (_32542_, _32541_, _06371_);
  or (_32543_, _32542_, _32538_);
  and (_32544_, _07945_, _08945_);
  or (_32545_, _32544_, _32485_);
  or (_32546_, _32545_, _07198_);
  and (_32547_, _32546_, _32543_);
  or (_32548_, _32547_, _06367_);
  and (_32549_, _14824_, _07945_);
  or (_32550_, _32549_, _32485_);
  or (_32551_, _32550_, _07218_);
  and (_32552_, _32551_, _07216_);
  and (_32553_, _32552_, _32548_);
  and (_32554_, _11214_, _07945_);
  or (_32555_, _32554_, _32485_);
  and (_32557_, _32555_, _06533_);
  or (_32558_, _32557_, _32553_);
  and (_32559_, _32558_, _07213_);
  or (_32560_, _32485_, _08397_);
  and (_32561_, _32545_, _06366_);
  and (_32562_, _32561_, _32560_);
  or (_32563_, _32562_, _32559_);
  and (_32564_, _32563_, _07210_);
  and (_32565_, _32494_, _06541_);
  and (_32566_, _32565_, _32560_);
  or (_32568_, _32566_, _06383_);
  or (_32569_, _32568_, _32564_);
  and (_32570_, _14821_, _07945_);
  or (_32571_, _32485_, _07231_);
  or (_32572_, _32571_, _32570_);
  and (_32573_, _32572_, _07229_);
  and (_32574_, _32573_, _32569_);
  nor (_32575_, _11213_, _13346_);
  or (_32576_, _32575_, _32485_);
  and (_32577_, _32576_, _06528_);
  or (_32579_, _32577_, _06563_);
  or (_32580_, _32579_, _32574_);
  or (_32581_, _32490_, _07241_);
  and (_32582_, _32581_, _06571_);
  and (_32583_, _32582_, _32580_);
  and (_32584_, _32516_, _06199_);
  or (_32585_, _32584_, _06188_);
  or (_32586_, _32585_, _32583_);
  and (_32587_, _14884_, _07945_);
  or (_32588_, _32485_, _06189_);
  or (_32590_, _32588_, _32587_);
  and (_32591_, _32590_, _01452_);
  and (_32592_, _32591_, _32586_);
  or (_43899_, _32592_, _32484_);
  and (_32593_, _13346_, \oc8051_golden_model_1.P1 [3]);
  nor (_32594_, _13346_, _07713_);
  or (_32595_, _32594_, _32593_);
  or (_32596_, _32595_, _07188_);
  or (_32597_, _32595_, _07142_);
  and (_32598_, _14898_, _07945_);
  or (_32600_, _32598_, _32593_);
  or (_32601_, _32600_, _06252_);
  and (_32602_, _07945_, \oc8051_golden_model_1.ACC [3]);
  or (_32603_, _32602_, _32593_);
  and (_32604_, _32603_, _07123_);
  and (_32605_, _07124_, \oc8051_golden_model_1.P1 [3]);
  or (_32606_, _32605_, _06251_);
  or (_32607_, _32606_, _32604_);
  and (_32608_, _32607_, _06476_);
  and (_32609_, _32608_, _32601_);
  and (_32611_, _13366_, \oc8051_golden_model_1.P1 [3]);
  and (_32612_, _14906_, _08531_);
  or (_32613_, _32612_, _32611_);
  and (_32614_, _32613_, _06475_);
  or (_32615_, _32614_, _06468_);
  or (_32616_, _32615_, _32609_);
  and (_32617_, _32616_, _32597_);
  or (_32618_, _32617_, _06466_);
  or (_32619_, _32603_, _06801_);
  and (_32620_, _32619_, _06484_);
  and (_32622_, _32620_, _32618_);
  and (_32623_, _14904_, _08531_);
  or (_32624_, _32623_, _32611_);
  and (_32625_, _32624_, _06483_);
  or (_32626_, _32625_, _06461_);
  or (_32627_, _32626_, _32622_);
  or (_32628_, _32611_, _14931_);
  and (_32629_, _32628_, _32613_);
  or (_32630_, _32629_, _07164_);
  and (_32631_, _32630_, _06242_);
  and (_32633_, _32631_, _32627_);
  or (_32634_, _32611_, _14947_);
  and (_32635_, _32634_, _06241_);
  and (_32636_, _32635_, _32613_);
  or (_32637_, _32636_, _07187_);
  or (_32638_, _32637_, _32633_);
  and (_32639_, _32638_, _32596_);
  or (_32640_, _32639_, _07182_);
  and (_32641_, _09205_, _07945_);
  or (_32642_, _32593_, _07183_);
  or (_32644_, _32642_, _32641_);
  and (_32645_, _32644_, _06336_);
  and (_32646_, _32645_, _32640_);
  and (_32647_, _15003_, _07945_);
  or (_32648_, _32647_, _32593_);
  and (_32649_, _32648_, _05968_);
  or (_32650_, _32649_, _06371_);
  or (_32651_, _32650_, _32646_);
  and (_32652_, _07945_, _08872_);
  or (_32653_, _32652_, _32593_);
  or (_32655_, _32653_, _07198_);
  and (_32656_, _32655_, _32651_);
  or (_32657_, _32656_, _06367_);
  and (_32658_, _15018_, _07945_);
  or (_32659_, _32658_, _32593_);
  or (_32660_, _32659_, _07218_);
  and (_32661_, _32660_, _07216_);
  and (_32662_, _32661_, _32657_);
  and (_32663_, _12523_, _07945_);
  or (_32664_, _32663_, _32593_);
  and (_32666_, _32664_, _06533_);
  or (_32667_, _32666_, _32662_);
  and (_32668_, _32667_, _07213_);
  or (_32669_, _32593_, _08257_);
  and (_32670_, _32653_, _06366_);
  and (_32671_, _32670_, _32669_);
  or (_32672_, _32671_, _32668_);
  and (_32673_, _32672_, _07210_);
  and (_32674_, _32603_, _06541_);
  and (_32675_, _32674_, _32669_);
  or (_32677_, _32675_, _06383_);
  or (_32678_, _32677_, _32673_);
  and (_32679_, _15015_, _07945_);
  or (_32680_, _32593_, _07231_);
  or (_32681_, _32680_, _32679_);
  and (_32682_, _32681_, _07229_);
  and (_32683_, _32682_, _32678_);
  nor (_32684_, _11211_, _13346_);
  or (_32685_, _32684_, _32593_);
  and (_32686_, _32685_, _06528_);
  or (_32688_, _32686_, _06563_);
  or (_32689_, _32688_, _32683_);
  or (_32690_, _32600_, _07241_);
  and (_32691_, _32690_, _06571_);
  and (_32692_, _32691_, _32689_);
  and (_32693_, _32624_, _06199_);
  or (_32694_, _32693_, _06188_);
  or (_32695_, _32694_, _32692_);
  and (_32696_, _15075_, _07945_);
  or (_32697_, _32593_, _06189_);
  or (_32699_, _32697_, _32696_);
  and (_32700_, _32699_, _01452_);
  and (_32701_, _32700_, _32695_);
  nor (_32702_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_32703_, _32702_, _00000_);
  or (_43900_, _32703_, _32701_);
  nor (_32704_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_32705_, _32704_, _00000_);
  and (_32706_, _13346_, \oc8051_golden_model_1.P1 [4]);
  nor (_32707_, _08494_, _13346_);
  or (_32709_, _32707_, _32706_);
  or (_32710_, _32709_, _07188_);
  and (_32711_, _13366_, \oc8051_golden_model_1.P1 [4]);
  and (_32712_, _15089_, _08531_);
  or (_32713_, _32712_, _32711_);
  and (_32714_, _32713_, _06483_);
  or (_32715_, _32709_, _07142_);
  and (_32716_, _15108_, _07945_);
  or (_32717_, _32716_, _32706_);
  or (_32718_, _32717_, _06252_);
  and (_32720_, _07945_, \oc8051_golden_model_1.ACC [4]);
  or (_32721_, _32720_, _32706_);
  and (_32722_, _32721_, _07123_);
  and (_32723_, _07124_, \oc8051_golden_model_1.P1 [4]);
  or (_32724_, _32723_, _06251_);
  or (_32725_, _32724_, _32722_);
  and (_32726_, _32725_, _06476_);
  and (_32727_, _32726_, _32718_);
  and (_32728_, _15091_, _08531_);
  or (_32729_, _32728_, _32711_);
  and (_32731_, _32729_, _06475_);
  or (_32732_, _32731_, _06468_);
  or (_32733_, _32732_, _32727_);
  and (_32734_, _32733_, _32715_);
  or (_32735_, _32734_, _06466_);
  or (_32736_, _32721_, _06801_);
  and (_32737_, _32736_, _06484_);
  and (_32738_, _32737_, _32735_);
  or (_32739_, _32738_, _32714_);
  and (_32740_, _32739_, _07164_);
  and (_32742_, _15126_, _08531_);
  or (_32743_, _32742_, _32711_);
  and (_32744_, _32743_, _06461_);
  or (_32745_, _32744_, _32740_);
  and (_32746_, _32745_, _06242_);
  or (_32747_, _32711_, _15141_);
  and (_32748_, _32747_, _06241_);
  and (_32749_, _32748_, _32729_);
  or (_32750_, _32749_, _07187_);
  or (_32751_, _32750_, _32746_);
  and (_32753_, _32751_, _32710_);
  or (_32754_, _32753_, _07182_);
  and (_32755_, _09159_, _07945_);
  or (_32756_, _32706_, _07183_);
  or (_32757_, _32756_, _32755_);
  and (_32758_, _32757_, _06336_);
  and (_32759_, _32758_, _32754_);
  and (_32760_, _15198_, _07945_);
  or (_32761_, _32760_, _32706_);
  and (_32762_, _32761_, _05968_);
  or (_32764_, _32762_, _06371_);
  or (_32765_, _32764_, _32759_);
  and (_32766_, _08892_, _07945_);
  or (_32767_, _32766_, _32706_);
  or (_32768_, _32767_, _07198_);
  and (_32769_, _32768_, _32765_);
  or (_32770_, _32769_, _06367_);
  and (_32771_, _15214_, _07945_);
  or (_32772_, _32771_, _32706_);
  or (_32773_, _32772_, _07218_);
  and (_32775_, _32773_, _07216_);
  and (_32776_, _32775_, _32770_);
  and (_32777_, _11209_, _07945_);
  or (_32778_, _32777_, _32706_);
  and (_32779_, _32778_, _06533_);
  or (_32780_, _32779_, _32776_);
  and (_32781_, _32780_, _07213_);
  or (_32782_, _32706_, _08497_);
  and (_32783_, _32767_, _06366_);
  and (_32784_, _32783_, _32782_);
  or (_32786_, _32784_, _32781_);
  and (_32787_, _32786_, _07210_);
  and (_32788_, _32721_, _06541_);
  and (_32789_, _32788_, _32782_);
  or (_32790_, _32789_, _06383_);
  or (_32791_, _32790_, _32787_);
  and (_32792_, _15211_, _07945_);
  or (_32793_, _32706_, _07231_);
  or (_32794_, _32793_, _32792_);
  and (_32795_, _32794_, _07229_);
  and (_32797_, _32795_, _32791_);
  nor (_32798_, _11208_, _13346_);
  or (_32799_, _32798_, _32706_);
  and (_32800_, _32799_, _06528_);
  or (_32801_, _32800_, _06563_);
  or (_32802_, _32801_, _32797_);
  or (_32803_, _32717_, _07241_);
  and (_32804_, _32803_, _06571_);
  and (_32805_, _32804_, _32802_);
  and (_32806_, _32713_, _06199_);
  or (_32808_, _32806_, _06188_);
  or (_32809_, _32808_, _32805_);
  and (_32810_, _15280_, _07945_);
  or (_32811_, _32706_, _06189_);
  or (_32812_, _32811_, _32810_);
  and (_32813_, _32812_, _01452_);
  and (_32814_, _32813_, _32809_);
  or (_43901_, _32814_, _32705_);
  and (_32815_, _13346_, \oc8051_golden_model_1.P1 [5]);
  nor (_32816_, _08209_, _13346_);
  or (_32818_, _32816_, _32815_);
  or (_32819_, _32818_, _07142_);
  and (_32820_, _15311_, _07945_);
  or (_32821_, _32820_, _32815_);
  or (_32822_, _32821_, _06252_);
  and (_32823_, _07945_, \oc8051_golden_model_1.ACC [5]);
  or (_32824_, _32823_, _32815_);
  and (_32825_, _32824_, _07123_);
  and (_32826_, _07124_, \oc8051_golden_model_1.P1 [5]);
  or (_32827_, _32826_, _06251_);
  or (_32829_, _32827_, _32825_);
  and (_32830_, _32829_, _06476_);
  and (_32831_, _32830_, _32822_);
  and (_32832_, _13366_, \oc8051_golden_model_1.P1 [5]);
  and (_32833_, _15296_, _08531_);
  or (_32834_, _32833_, _32832_);
  and (_32835_, _32834_, _06475_);
  or (_32836_, _32835_, _06468_);
  or (_32837_, _32836_, _32831_);
  and (_32838_, _32837_, _32819_);
  or (_32840_, _32838_, _06466_);
  or (_32841_, _32824_, _06801_);
  and (_32842_, _32841_, _06484_);
  and (_32843_, _32842_, _32840_);
  and (_32844_, _15294_, _08531_);
  or (_32845_, _32844_, _32832_);
  and (_32846_, _32845_, _06483_);
  or (_32847_, _32846_, _06461_);
  or (_32848_, _32847_, _32843_);
  or (_32849_, _32832_, _15328_);
  and (_32851_, _32849_, _32834_);
  or (_32852_, _32851_, _07164_);
  and (_32853_, _32852_, _06242_);
  and (_32854_, _32853_, _32848_);
  or (_32855_, _32832_, _15344_);
  and (_32856_, _32855_, _06241_);
  and (_32857_, _32856_, _32834_);
  or (_32858_, _32857_, _07187_);
  or (_32859_, _32858_, _32854_);
  or (_32860_, _32818_, _07188_);
  and (_32862_, _32860_, _32859_);
  or (_32863_, _32862_, _07182_);
  and (_32864_, _09113_, _07945_);
  or (_32865_, _32815_, _07183_);
  or (_32866_, _32865_, _32864_);
  and (_32867_, _32866_, _06336_);
  and (_32868_, _32867_, _32863_);
  and (_32869_, _15400_, _07945_);
  or (_32870_, _32869_, _32815_);
  and (_32871_, _32870_, _05968_);
  or (_32873_, _32871_, _06371_);
  or (_32874_, _32873_, _32868_);
  and (_32875_, _08888_, _07945_);
  or (_32876_, _32875_, _32815_);
  or (_32877_, _32876_, _07198_);
  and (_32878_, _32877_, _32874_);
  or (_32879_, _32878_, _06367_);
  and (_32880_, _15416_, _07945_);
  or (_32881_, _32880_, _32815_);
  or (_32882_, _32881_, _07218_);
  and (_32884_, _32882_, _07216_);
  and (_32885_, _32884_, _32879_);
  and (_32886_, _11205_, _07945_);
  or (_32887_, _32886_, _32815_);
  and (_32888_, _32887_, _06533_);
  or (_32889_, _32888_, _32885_);
  and (_32890_, _32889_, _07213_);
  or (_32891_, _32815_, _08212_);
  and (_32892_, _32876_, _06366_);
  and (_32893_, _32892_, _32891_);
  or (_32895_, _32893_, _32890_);
  and (_32896_, _32895_, _07210_);
  and (_32897_, _32824_, _06541_);
  and (_32898_, _32897_, _32891_);
  or (_32899_, _32898_, _06383_);
  or (_32900_, _32899_, _32896_);
  and (_32901_, _15413_, _07945_);
  or (_32902_, _32815_, _07231_);
  or (_32903_, _32902_, _32901_);
  and (_32904_, _32903_, _07229_);
  and (_32906_, _32904_, _32900_);
  nor (_32907_, _11204_, _13346_);
  or (_32908_, _32907_, _32815_);
  and (_32909_, _32908_, _06528_);
  or (_32910_, _32909_, _06563_);
  or (_32911_, _32910_, _32906_);
  or (_32912_, _32821_, _07241_);
  and (_32913_, _32912_, _06571_);
  and (_32914_, _32913_, _32911_);
  and (_32915_, _32845_, _06199_);
  or (_32917_, _32915_, _06188_);
  or (_32918_, _32917_, _32914_);
  and (_32919_, _15477_, _07945_);
  or (_32920_, _32815_, _06189_);
  or (_32921_, _32920_, _32919_);
  and (_32922_, _32921_, _01452_);
  and (_32923_, _32922_, _32918_);
  nor (_32924_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_32925_, _32924_, _00000_);
  or (_43902_, _32925_, _32923_);
  and (_32927_, _13346_, \oc8051_golden_model_1.P1 [6]);
  nor (_32928_, _08106_, _13346_);
  or (_32929_, _32928_, _32927_);
  or (_32930_, _32929_, _07142_);
  and (_32931_, _15512_, _07945_);
  or (_32932_, _32931_, _32927_);
  or (_32933_, _32932_, _06252_);
  and (_32934_, _07945_, \oc8051_golden_model_1.ACC [6]);
  or (_32935_, _32934_, _32927_);
  and (_32936_, _32935_, _07123_);
  and (_32938_, _07124_, \oc8051_golden_model_1.P1 [6]);
  or (_32939_, _32938_, _06251_);
  or (_32940_, _32939_, _32936_);
  and (_32941_, _32940_, _06476_);
  and (_32942_, _32941_, _32933_);
  and (_32943_, _13366_, \oc8051_golden_model_1.P1 [6]);
  and (_32944_, _15499_, _08531_);
  or (_32945_, _32944_, _32943_);
  and (_32946_, _32945_, _06475_);
  or (_32947_, _32946_, _06468_);
  or (_32949_, _32947_, _32942_);
  and (_32950_, _32949_, _32930_);
  or (_32951_, _32950_, _06466_);
  or (_32952_, _32935_, _06801_);
  and (_32953_, _32952_, _06484_);
  and (_32954_, _32953_, _32951_);
  and (_32955_, _15497_, _08531_);
  or (_32956_, _32955_, _32943_);
  and (_32957_, _32956_, _06483_);
  or (_32958_, _32957_, _06461_);
  or (_32960_, _32958_, _32954_);
  or (_32961_, _32943_, _15529_);
  and (_32962_, _32961_, _32945_);
  or (_32963_, _32962_, _07164_);
  and (_32964_, _32963_, _06242_);
  and (_32965_, _32964_, _32960_);
  or (_32966_, _32943_, _15545_);
  and (_32967_, _32966_, _06241_);
  and (_32968_, _32967_, _32945_);
  or (_32969_, _32968_, _07187_);
  or (_32971_, _32969_, _32965_);
  or (_32972_, _32929_, _07188_);
  and (_32973_, _32972_, _32971_);
  or (_32974_, _32973_, _07182_);
  and (_32975_, _09067_, _07945_);
  or (_32976_, _32927_, _07183_);
  or (_32977_, _32976_, _32975_);
  and (_32978_, _32977_, _06336_);
  and (_32979_, _32978_, _32974_);
  and (_32980_, _15601_, _07945_);
  or (_32982_, _32980_, _32927_);
  and (_32983_, _32982_, _05968_);
  or (_32984_, _32983_, _06371_);
  or (_32985_, _32984_, _32979_);
  and (_32986_, _15608_, _07945_);
  or (_32987_, _32986_, _32927_);
  or (_32988_, _32987_, _07198_);
  and (_32989_, _32988_, _32985_);
  or (_32990_, _32989_, _06367_);
  and (_32991_, _15618_, _07945_);
  or (_32993_, _32991_, _32927_);
  or (_32994_, _32993_, _07218_);
  and (_32995_, _32994_, _07216_);
  and (_32996_, _32995_, _32990_);
  and (_32997_, _11202_, _07945_);
  or (_32998_, _32997_, _32927_);
  and (_32999_, _32998_, _06533_);
  or (_33000_, _32999_, _32996_);
  and (_33001_, _33000_, _07213_);
  or (_33002_, _32927_, _08109_);
  and (_33004_, _32987_, _06366_);
  and (_33005_, _33004_, _33002_);
  or (_33006_, _33005_, _33001_);
  and (_33007_, _33006_, _07210_);
  and (_33008_, _32935_, _06541_);
  and (_33009_, _33008_, _33002_);
  or (_33010_, _33009_, _06383_);
  or (_33011_, _33010_, _33007_);
  and (_33012_, _15615_, _07945_);
  or (_33013_, _32927_, _07231_);
  or (_33015_, _33013_, _33012_);
  and (_33016_, _33015_, _07229_);
  and (_33017_, _33016_, _33011_);
  nor (_33018_, _11201_, _13346_);
  or (_33019_, _33018_, _32927_);
  and (_33020_, _33019_, _06528_);
  or (_33021_, _33020_, _06563_);
  or (_33022_, _33021_, _33017_);
  or (_33023_, _32932_, _07241_);
  and (_33024_, _33023_, _06571_);
  and (_33026_, _33024_, _33022_);
  and (_33027_, _32956_, _06199_);
  or (_33028_, _33027_, _06188_);
  or (_33029_, _33028_, _33026_);
  and (_33030_, _15676_, _07945_);
  or (_33031_, _32927_, _06189_);
  or (_33032_, _33031_, _33030_);
  and (_33033_, _33032_, _01452_);
  and (_33034_, _33033_, _33029_);
  nor (_33035_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_33037_, _33035_, _00000_);
  or (_43903_, _33037_, _33034_);
  and (_33038_, _01456_, \oc8051_golden_model_1.IP [0]);
  and (_33039_, _07918_, \oc8051_golden_model_1.ACC [0]);
  and (_33040_, _33039_, _08351_);
  and (_33041_, _13448_, \oc8051_golden_model_1.IP [0]);
  or (_33042_, _33041_, _07210_);
  or (_33043_, _33042_, _33040_);
  and (_33044_, _07918_, _07325_);
  or (_33045_, _33044_, _33041_);
  or (_33047_, _33045_, _07188_);
  and (_33048_, _13468_, \oc8051_golden_model_1.IP [0]);
  and (_33049_, _14341_, _08541_);
  or (_33050_, _33049_, _33048_);
  and (_33051_, _33050_, _06475_);
  nor (_33052_, _08351_, _13448_);
  or (_33053_, _33052_, _33041_);
  or (_33054_, _33053_, _06252_);
  or (_33055_, _33039_, _33041_);
  and (_33056_, _33055_, _07123_);
  and (_33058_, _07124_, \oc8051_golden_model_1.IP [0]);
  or (_33059_, _33058_, _06251_);
  or (_33060_, _33059_, _33056_);
  and (_33061_, _33060_, _06476_);
  and (_33062_, _33061_, _33054_);
  or (_33063_, _33062_, _33051_);
  and (_33064_, _33063_, _07142_);
  and (_33065_, _33045_, _06468_);
  or (_33066_, _33065_, _06466_);
  or (_33067_, _33066_, _33064_);
  or (_33069_, _33055_, _06801_);
  and (_33070_, _33069_, _06484_);
  and (_33071_, _33070_, _33067_);
  and (_33072_, _33041_, _06483_);
  or (_33073_, _33072_, _06461_);
  or (_33074_, _33073_, _33071_);
  or (_33075_, _33053_, _07164_);
  and (_33076_, _33075_, _06242_);
  and (_33077_, _33076_, _33074_);
  or (_33078_, _33048_, _14371_);
  and (_33080_, _33078_, _06241_);
  and (_33081_, _33080_, _33050_);
  or (_33082_, _33081_, _07187_);
  or (_33083_, _33082_, _33077_);
  and (_33084_, _33083_, _33047_);
  or (_33085_, _33084_, _07182_);
  and (_33086_, _09342_, _07918_);
  or (_33087_, _33041_, _07183_);
  or (_33088_, _33087_, _33086_);
  and (_33089_, _33088_, _33085_);
  or (_33091_, _33089_, _05968_);
  and (_33092_, _14427_, _07918_);
  or (_33093_, _33041_, _06336_);
  or (_33094_, _33093_, _33092_);
  and (_33095_, _33094_, _07198_);
  and (_33096_, _33095_, _33091_);
  and (_33097_, _07918_, _08908_);
  or (_33098_, _33097_, _33041_);
  and (_33099_, _33098_, _06371_);
  or (_33100_, _33099_, _06367_);
  or (_33102_, _33100_, _33096_);
  and (_33103_, _14442_, _07918_);
  or (_33104_, _33103_, _33041_);
  or (_33105_, _33104_, _07218_);
  and (_33106_, _33105_, _07216_);
  and (_33107_, _33106_, _33102_);
  nor (_33108_, _12526_, _13448_);
  or (_33109_, _33108_, _33041_);
  nor (_33110_, _33040_, _07216_);
  and (_33111_, _33110_, _33109_);
  or (_33113_, _33111_, _33107_);
  and (_33114_, _33113_, _07213_);
  nand (_33115_, _33098_, _06366_);
  nor (_33116_, _33115_, _33052_);
  or (_33117_, _33116_, _06541_);
  or (_33118_, _33117_, _33114_);
  and (_33119_, _33118_, _33043_);
  or (_33120_, _33119_, _06383_);
  and (_33121_, _14325_, _07918_);
  or (_33122_, _33121_, _33041_);
  or (_33124_, _33122_, _07231_);
  and (_33125_, _33124_, _07229_);
  and (_33126_, _33125_, _33120_);
  and (_33127_, _33109_, _06528_);
  or (_33128_, _33127_, _06563_);
  or (_33129_, _33128_, _33126_);
  or (_33130_, _33053_, _07241_);
  and (_33131_, _33130_, _33129_);
  or (_33132_, _33131_, _06199_);
  or (_33133_, _33041_, _06571_);
  and (_33135_, _33133_, _33132_);
  or (_33136_, _33135_, _06188_);
  or (_33137_, _33053_, _06189_);
  and (_33138_, _33137_, _01452_);
  and (_33139_, _33138_, _33136_);
  or (_33140_, _33139_, _33038_);
  and (_43904_, _33140_, _43223_);
  not (_33141_, \oc8051_golden_model_1.IP [1]);
  nor (_33142_, _01452_, _33141_);
  nor (_33143_, _07918_, _33141_);
  nor (_33145_, _11216_, _13448_);
  or (_33146_, _33145_, _33143_);
  or (_33147_, _33146_, _07229_);
  nand (_33148_, _07918_, _07018_);
  or (_33149_, _07918_, \oc8051_golden_model_1.IP [1]);
  and (_33150_, _33149_, _06371_);
  and (_33151_, _33150_, _33148_);
  nor (_33152_, _13448_, _07120_);
  or (_33153_, _33152_, _33143_);
  or (_33154_, _33153_, _07142_);
  and (_33156_, _14503_, _07918_);
  not (_33157_, _33156_);
  and (_33158_, _33157_, _33149_);
  or (_33159_, _33158_, _06252_);
  and (_33160_, _07918_, \oc8051_golden_model_1.ACC [1]);
  or (_33161_, _33160_, _33143_);
  and (_33162_, _33161_, _07123_);
  nor (_33163_, _07123_, _33141_);
  or (_33164_, _33163_, _06251_);
  or (_33165_, _33164_, _33162_);
  and (_33167_, _33165_, _06476_);
  and (_33168_, _33167_, _33159_);
  nor (_33169_, _08541_, _33141_);
  and (_33170_, _14510_, _08541_);
  or (_33171_, _33170_, _33169_);
  and (_33172_, _33171_, _06475_);
  or (_33173_, _33172_, _06468_);
  or (_33174_, _33173_, _33168_);
  and (_33175_, _33174_, _33154_);
  or (_33176_, _33175_, _06466_);
  or (_33178_, _33161_, _06801_);
  and (_33179_, _33178_, _06484_);
  and (_33180_, _33179_, _33176_);
  and (_33181_, _14513_, _08541_);
  or (_33182_, _33181_, _33169_);
  and (_33183_, _33182_, _06483_);
  or (_33184_, _33183_, _06461_);
  or (_33185_, _33184_, _33180_);
  or (_33186_, _33169_, _14509_);
  and (_33187_, _33186_, _33171_);
  or (_33189_, _33187_, _07164_);
  and (_33190_, _33189_, _06242_);
  and (_33191_, _33190_, _33185_);
  or (_33192_, _33169_, _14553_);
  and (_33193_, _33192_, _06241_);
  and (_33194_, _33193_, _33171_);
  or (_33195_, _33194_, _07187_);
  or (_33196_, _33195_, _33191_);
  or (_33197_, _33153_, _07188_);
  and (_33198_, _33197_, _33196_);
  or (_33200_, _33198_, _07182_);
  and (_33201_, _09297_, _07918_);
  or (_33202_, _33143_, _07183_);
  or (_33203_, _33202_, _33201_);
  and (_33204_, _33203_, _06336_);
  and (_33205_, _33204_, _33200_);
  and (_33206_, _14609_, _07918_);
  or (_33207_, _33206_, _33143_);
  and (_33208_, _33207_, _05968_);
  or (_33209_, _33208_, _33205_);
  and (_33211_, _33209_, _07198_);
  or (_33212_, _33211_, _33151_);
  and (_33213_, _33212_, _07218_);
  or (_33214_, _14625_, _13448_);
  and (_33215_, _33149_, _06367_);
  and (_33216_, _33215_, _33214_);
  or (_33217_, _33216_, _06533_);
  or (_33218_, _33217_, _33213_);
  nand (_33219_, _11215_, _07918_);
  and (_33220_, _33219_, _33146_);
  or (_33222_, _33220_, _07216_);
  and (_33223_, _33222_, _07213_);
  and (_33224_, _33223_, _33218_);
  or (_33225_, _14623_, _13448_);
  and (_33226_, _33149_, _06366_);
  and (_33227_, _33226_, _33225_);
  or (_33228_, _33227_, _06541_);
  or (_33229_, _33228_, _33224_);
  nor (_33230_, _33143_, _07210_);
  nand (_33231_, _33230_, _33219_);
  and (_33233_, _33231_, _07231_);
  and (_33234_, _33233_, _33229_);
  or (_33235_, _33148_, _08302_);
  and (_33236_, _33149_, _06383_);
  and (_33237_, _33236_, _33235_);
  or (_33238_, _33237_, _06528_);
  or (_33239_, _33238_, _33234_);
  and (_33240_, _33239_, _33147_);
  or (_33241_, _33240_, _06563_);
  or (_33242_, _33158_, _07241_);
  and (_33244_, _33242_, _06571_);
  and (_33245_, _33244_, _33241_);
  and (_33246_, _33182_, _06199_);
  or (_33247_, _33246_, _06188_);
  or (_33248_, _33247_, _33245_);
  or (_33249_, _33143_, _06189_);
  or (_33250_, _33249_, _33156_);
  and (_33251_, _33250_, _01452_);
  and (_33252_, _33251_, _33248_);
  or (_33253_, _33252_, _33142_);
  and (_43905_, _33253_, _43223_);
  and (_33255_, _01456_, \oc8051_golden_model_1.IP [2]);
  and (_33256_, _13448_, \oc8051_golden_model_1.IP [2]);
  nor (_33257_, _13448_, _07578_);
  or (_33258_, _33257_, _33256_);
  or (_33259_, _33258_, _07188_);
  and (_33260_, _14712_, _07918_);
  or (_33261_, _33260_, _33256_);
  or (_33262_, _33261_, _06252_);
  and (_33263_, _07918_, \oc8051_golden_model_1.ACC [2]);
  or (_33265_, _33263_, _33256_);
  and (_33266_, _33265_, _07123_);
  and (_33267_, _07124_, \oc8051_golden_model_1.IP [2]);
  or (_33268_, _33267_, _06251_);
  or (_33269_, _33268_, _33266_);
  and (_33270_, _33269_, _06476_);
  and (_33271_, _33270_, _33262_);
  and (_33272_, _13468_, \oc8051_golden_model_1.IP [2]);
  and (_33273_, _14702_, _08541_);
  or (_33274_, _33273_, _33272_);
  and (_33276_, _33274_, _06475_);
  or (_33277_, _33276_, _06468_);
  or (_33278_, _33277_, _33271_);
  or (_33279_, _33258_, _07142_);
  and (_33280_, _33279_, _33278_);
  or (_33281_, _33280_, _06466_);
  or (_33282_, _33265_, _06801_);
  and (_33283_, _33282_, _06484_);
  and (_33284_, _33283_, _33281_);
  and (_33285_, _14706_, _08541_);
  or (_33286_, _33285_, _33272_);
  and (_33287_, _33286_, _06483_);
  or (_33288_, _33287_, _06461_);
  or (_33289_, _33288_, _33284_);
  or (_33290_, _33272_, _14739_);
  and (_33291_, _33290_, _33274_);
  or (_33292_, _33291_, _07164_);
  and (_33293_, _33292_, _06242_);
  and (_33294_, _33293_, _33289_);
  or (_33295_, _33272_, _14703_);
  and (_33297_, _33295_, _06241_);
  and (_33298_, _33297_, _33274_);
  or (_33299_, _33298_, _07187_);
  or (_33300_, _33299_, _33294_);
  and (_33301_, _33300_, _33259_);
  or (_33302_, _33301_, _07182_);
  and (_33303_, _09251_, _07918_);
  or (_33304_, _33256_, _07183_);
  or (_33305_, _33304_, _33303_);
  and (_33306_, _33305_, _06336_);
  and (_33308_, _33306_, _33302_);
  and (_33309_, _14808_, _07918_);
  or (_33310_, _33309_, _33256_);
  and (_33311_, _33310_, _05968_);
  or (_33312_, _33311_, _06371_);
  or (_33313_, _33312_, _33308_);
  and (_33314_, _07918_, _08945_);
  or (_33315_, _33314_, _33256_);
  or (_33316_, _33315_, _07198_);
  and (_33317_, _33316_, _33313_);
  or (_33319_, _33317_, _06367_);
  and (_33320_, _14824_, _07918_);
  or (_33321_, _33320_, _33256_);
  or (_33322_, _33321_, _07218_);
  and (_33323_, _33322_, _07216_);
  and (_33324_, _33323_, _33319_);
  and (_33325_, _11214_, _07918_);
  or (_33326_, _33325_, _33256_);
  and (_33327_, _33326_, _06533_);
  or (_33328_, _33327_, _33324_);
  and (_33330_, _33328_, _07213_);
  or (_33331_, _33256_, _08397_);
  and (_33332_, _33315_, _06366_);
  and (_33333_, _33332_, _33331_);
  or (_33334_, _33333_, _33330_);
  and (_33335_, _33334_, _07210_);
  and (_33336_, _33265_, _06541_);
  and (_33337_, _33336_, _33331_);
  or (_33338_, _33337_, _06383_);
  or (_33339_, _33338_, _33335_);
  and (_33341_, _14821_, _07918_);
  or (_33342_, _33256_, _07231_);
  or (_33343_, _33342_, _33341_);
  and (_33344_, _33343_, _07229_);
  and (_33345_, _33344_, _33339_);
  nor (_33346_, _11213_, _13448_);
  or (_33347_, _33346_, _33256_);
  and (_33348_, _33347_, _06528_);
  or (_33349_, _33348_, _06563_);
  or (_33350_, _33349_, _33345_);
  or (_33352_, _33261_, _07241_);
  and (_33353_, _33352_, _06571_);
  and (_33354_, _33353_, _33350_);
  and (_33355_, _33286_, _06199_);
  or (_33356_, _33355_, _06188_);
  or (_33357_, _33356_, _33354_);
  and (_33358_, _14884_, _07918_);
  or (_33359_, _33256_, _06189_);
  or (_33360_, _33359_, _33358_);
  and (_33361_, _33360_, _01452_);
  and (_33363_, _33361_, _33357_);
  or (_33364_, _33363_, _33255_);
  and (_43906_, _33364_, _43223_);
  and (_33365_, _01456_, \oc8051_golden_model_1.IP [3]);
  and (_33366_, _13448_, \oc8051_golden_model_1.IP [3]);
  nor (_33367_, _13448_, _07713_);
  or (_33368_, _33367_, _33366_);
  or (_33369_, _33368_, _07188_);
  or (_33370_, _33368_, _07142_);
  and (_33371_, _14898_, _07918_);
  or (_33373_, _33371_, _33366_);
  or (_33374_, _33373_, _06252_);
  and (_33375_, _07918_, \oc8051_golden_model_1.ACC [3]);
  or (_33376_, _33375_, _33366_);
  and (_33377_, _33376_, _07123_);
  and (_33378_, _07124_, \oc8051_golden_model_1.IP [3]);
  or (_33379_, _33378_, _06251_);
  or (_33380_, _33379_, _33377_);
  and (_33381_, _33380_, _06476_);
  and (_33382_, _33381_, _33374_);
  and (_33384_, _13468_, \oc8051_golden_model_1.IP [3]);
  and (_33385_, _14906_, _08541_);
  or (_33386_, _33385_, _33384_);
  and (_33387_, _33386_, _06475_);
  or (_33388_, _33387_, _06468_);
  or (_33389_, _33388_, _33382_);
  and (_33390_, _33389_, _33370_);
  or (_33391_, _33390_, _06466_);
  or (_33392_, _33376_, _06801_);
  and (_33393_, _33392_, _06484_);
  and (_33395_, _33393_, _33391_);
  and (_33396_, _14904_, _08541_);
  or (_33397_, _33396_, _33384_);
  and (_33398_, _33397_, _06483_);
  or (_33399_, _33398_, _06461_);
  or (_33400_, _33399_, _33395_);
  or (_33401_, _33384_, _14931_);
  and (_33402_, _33401_, _33386_);
  or (_33403_, _33402_, _07164_);
  and (_33404_, _33403_, _06242_);
  and (_33406_, _33404_, _33400_);
  or (_33407_, _33384_, _14947_);
  and (_33408_, _33407_, _06241_);
  and (_33409_, _33408_, _33386_);
  or (_33410_, _33409_, _07187_);
  or (_33411_, _33410_, _33406_);
  and (_33412_, _33411_, _33369_);
  or (_33413_, _33412_, _07182_);
  and (_33414_, _09205_, _07918_);
  or (_33415_, _33366_, _07183_);
  or (_33417_, _33415_, _33414_);
  and (_33418_, _33417_, _06336_);
  and (_33419_, _33418_, _33413_);
  and (_33420_, _15003_, _07918_);
  or (_33421_, _33420_, _33366_);
  and (_33422_, _33421_, _05968_);
  or (_33423_, _33422_, _06371_);
  or (_33424_, _33423_, _33419_);
  and (_33425_, _07918_, _08872_);
  or (_33426_, _33425_, _33366_);
  or (_33428_, _33426_, _07198_);
  and (_33429_, _33428_, _33424_);
  or (_33430_, _33429_, _06367_);
  and (_33431_, _15018_, _07918_);
  or (_33432_, _33431_, _33366_);
  or (_33433_, _33432_, _07218_);
  and (_33434_, _33433_, _07216_);
  and (_33435_, _33434_, _33430_);
  and (_33436_, _12523_, _07918_);
  or (_33437_, _33436_, _33366_);
  and (_33439_, _33437_, _06533_);
  or (_33440_, _33439_, _33435_);
  and (_33441_, _33440_, _07213_);
  or (_33442_, _33366_, _08257_);
  and (_33443_, _33426_, _06366_);
  and (_33444_, _33443_, _33442_);
  or (_33445_, _33444_, _33441_);
  and (_33446_, _33445_, _07210_);
  and (_33447_, _33376_, _06541_);
  and (_33448_, _33447_, _33442_);
  or (_33450_, _33448_, _06383_);
  or (_33451_, _33450_, _33446_);
  and (_33452_, _15015_, _07918_);
  or (_33453_, _33366_, _07231_);
  or (_33454_, _33453_, _33452_);
  and (_33455_, _33454_, _07229_);
  and (_33456_, _33455_, _33451_);
  nor (_33457_, _11211_, _13448_);
  or (_33458_, _33457_, _33366_);
  and (_33459_, _33458_, _06528_);
  or (_33461_, _33459_, _06563_);
  or (_33462_, _33461_, _33456_);
  or (_33463_, _33373_, _07241_);
  and (_33464_, _33463_, _06571_);
  and (_33465_, _33464_, _33462_);
  and (_33466_, _33397_, _06199_);
  or (_33467_, _33466_, _06188_);
  or (_33468_, _33467_, _33465_);
  and (_33469_, _15075_, _07918_);
  or (_33470_, _33366_, _06189_);
  or (_33472_, _33470_, _33469_);
  and (_33473_, _33472_, _01452_);
  and (_33474_, _33473_, _33468_);
  or (_33475_, _33474_, _33365_);
  and (_43907_, _33475_, _43223_);
  and (_33476_, _01456_, \oc8051_golden_model_1.IP [4]);
  and (_33477_, _13448_, \oc8051_golden_model_1.IP [4]);
  nor (_33478_, _08494_, _13448_);
  or (_33479_, _33478_, _33477_);
  or (_33480_, _33479_, _07188_);
  and (_33482_, _13468_, \oc8051_golden_model_1.IP [4]);
  and (_33483_, _15089_, _08541_);
  or (_33484_, _33483_, _33482_);
  and (_33485_, _33484_, _06483_);
  or (_33486_, _33479_, _07142_);
  and (_33487_, _15108_, _07918_);
  or (_33488_, _33487_, _33477_);
  or (_33489_, _33488_, _06252_);
  and (_33490_, _07918_, \oc8051_golden_model_1.ACC [4]);
  or (_33491_, _33490_, _33477_);
  and (_33493_, _33491_, _07123_);
  and (_33494_, _07124_, \oc8051_golden_model_1.IP [4]);
  or (_33495_, _33494_, _06251_);
  or (_33496_, _33495_, _33493_);
  and (_33497_, _33496_, _06476_);
  and (_33498_, _33497_, _33489_);
  and (_33499_, _15091_, _08541_);
  or (_33500_, _33499_, _33482_);
  and (_33501_, _33500_, _06475_);
  or (_33502_, _33501_, _06468_);
  or (_33504_, _33502_, _33498_);
  and (_33505_, _33504_, _33486_);
  or (_33506_, _33505_, _06466_);
  or (_33507_, _33491_, _06801_);
  and (_33508_, _33507_, _06484_);
  and (_33509_, _33508_, _33506_);
  or (_33510_, _33509_, _33485_);
  and (_33511_, _33510_, _07164_);
  or (_33512_, _33482_, _15125_);
  and (_33513_, _33512_, _06461_);
  and (_33515_, _33513_, _33500_);
  or (_33516_, _33515_, _33511_);
  and (_33517_, _33516_, _06242_);
  or (_33518_, _33482_, _15141_);
  and (_33519_, _33518_, _06241_);
  and (_33520_, _33519_, _33500_);
  or (_33521_, _33520_, _07187_);
  or (_33522_, _33521_, _33517_);
  and (_33523_, _33522_, _33480_);
  or (_33524_, _33523_, _07182_);
  and (_33526_, _09159_, _07918_);
  or (_33527_, _33477_, _07183_);
  or (_33528_, _33527_, _33526_);
  and (_33529_, _33528_, _06336_);
  and (_33530_, _33529_, _33524_);
  and (_33531_, _15198_, _07918_);
  or (_33532_, _33531_, _33477_);
  and (_33533_, _33532_, _05968_);
  or (_33534_, _33533_, _06371_);
  or (_33535_, _33534_, _33530_);
  and (_33537_, _08892_, _07918_);
  or (_33538_, _33537_, _33477_);
  or (_33539_, _33538_, _07198_);
  and (_33540_, _33539_, _33535_);
  or (_33541_, _33540_, _06367_);
  and (_33542_, _15214_, _07918_);
  or (_33543_, _33542_, _33477_);
  or (_33544_, _33543_, _07218_);
  and (_33545_, _33544_, _07216_);
  and (_33546_, _33545_, _33541_);
  and (_33548_, _11209_, _07918_);
  or (_33549_, _33548_, _33477_);
  and (_33550_, _33549_, _06533_);
  or (_33551_, _33550_, _33546_);
  and (_33552_, _33551_, _07213_);
  or (_33553_, _33477_, _08497_);
  and (_33554_, _33538_, _06366_);
  and (_33555_, _33554_, _33553_);
  or (_33556_, _33555_, _33552_);
  and (_33557_, _33556_, _07210_);
  and (_33559_, _33491_, _06541_);
  and (_33560_, _33559_, _33553_);
  or (_33561_, _33560_, _06383_);
  or (_33562_, _33561_, _33557_);
  and (_33563_, _15211_, _07918_);
  or (_33564_, _33477_, _07231_);
  or (_33565_, _33564_, _33563_);
  and (_33566_, _33565_, _07229_);
  and (_33567_, _33566_, _33562_);
  nor (_33568_, _11208_, _13448_);
  or (_33570_, _33568_, _33477_);
  and (_33571_, _33570_, _06528_);
  or (_33572_, _33571_, _06563_);
  or (_33573_, _33572_, _33567_);
  or (_33574_, _33488_, _07241_);
  and (_33575_, _33574_, _06571_);
  and (_33576_, _33575_, _33573_);
  and (_33577_, _33484_, _06199_);
  or (_33578_, _33577_, _06188_);
  or (_33579_, _33578_, _33576_);
  and (_33581_, _15280_, _07918_);
  or (_33582_, _33477_, _06189_);
  or (_33583_, _33582_, _33581_);
  and (_33584_, _33583_, _01452_);
  and (_33585_, _33584_, _33579_);
  or (_33586_, _33585_, _33476_);
  and (_43908_, _33586_, _43223_);
  and (_33587_, _01456_, \oc8051_golden_model_1.IP [5]);
  and (_33588_, _13448_, \oc8051_golden_model_1.IP [5]);
  nor (_33589_, _08209_, _13448_);
  or (_33591_, _33589_, _33588_);
  or (_33592_, _33591_, _07142_);
  and (_33593_, _15311_, _07918_);
  or (_33594_, _33593_, _33588_);
  or (_33595_, _33594_, _06252_);
  and (_33596_, _07918_, \oc8051_golden_model_1.ACC [5]);
  or (_33597_, _33596_, _33588_);
  and (_33598_, _33597_, _07123_);
  and (_33599_, _07124_, \oc8051_golden_model_1.IP [5]);
  or (_33600_, _33599_, _06251_);
  or (_33602_, _33600_, _33598_);
  and (_33603_, _33602_, _06476_);
  and (_33604_, _33603_, _33595_);
  and (_33605_, _13468_, \oc8051_golden_model_1.IP [5]);
  and (_33606_, _15296_, _08541_);
  or (_33607_, _33606_, _33605_);
  and (_33608_, _33607_, _06475_);
  or (_33609_, _33608_, _06468_);
  or (_33610_, _33609_, _33604_);
  and (_33611_, _33610_, _33592_);
  or (_33613_, _33611_, _06466_);
  or (_33614_, _33597_, _06801_);
  and (_33615_, _33614_, _06484_);
  and (_33616_, _33615_, _33613_);
  and (_33617_, _15294_, _08541_);
  or (_33618_, _33617_, _33605_);
  and (_33619_, _33618_, _06483_);
  or (_33620_, _33619_, _06461_);
  or (_33621_, _33620_, _33616_);
  or (_33622_, _33605_, _15328_);
  and (_33624_, _33622_, _33607_);
  or (_33625_, _33624_, _07164_);
  and (_33626_, _33625_, _06242_);
  and (_33627_, _33626_, _33621_);
  or (_33628_, _33605_, _15344_);
  and (_33629_, _33628_, _06241_);
  and (_33630_, _33629_, _33607_);
  or (_33631_, _33630_, _07187_);
  or (_33632_, _33631_, _33627_);
  or (_33633_, _33591_, _07188_);
  and (_33635_, _33633_, _33632_);
  or (_33636_, _33635_, _07182_);
  and (_33637_, _09113_, _07918_);
  or (_33638_, _33588_, _07183_);
  or (_33639_, _33638_, _33637_);
  and (_33640_, _33639_, _06336_);
  and (_33641_, _33640_, _33636_);
  and (_33642_, _15400_, _07918_);
  or (_33643_, _33642_, _33588_);
  and (_33644_, _33643_, _05968_);
  or (_33646_, _33644_, _06371_);
  or (_33647_, _33646_, _33641_);
  and (_33648_, _08888_, _07918_);
  or (_33649_, _33648_, _33588_);
  or (_33650_, _33649_, _07198_);
  and (_33651_, _33650_, _33647_);
  or (_33652_, _33651_, _06367_);
  and (_33653_, _15416_, _07918_);
  or (_33654_, _33653_, _33588_);
  or (_33655_, _33654_, _07218_);
  and (_33657_, _33655_, _07216_);
  and (_33658_, _33657_, _33652_);
  and (_33659_, _11205_, _07918_);
  or (_33660_, _33659_, _33588_);
  and (_33661_, _33660_, _06533_);
  or (_33662_, _33661_, _33658_);
  and (_33663_, _33662_, _07213_);
  or (_33664_, _33588_, _08212_);
  and (_33665_, _33649_, _06366_);
  and (_33666_, _33665_, _33664_);
  or (_33668_, _33666_, _33663_);
  and (_33669_, _33668_, _07210_);
  and (_33670_, _33597_, _06541_);
  and (_33671_, _33670_, _33664_);
  or (_33672_, _33671_, _06383_);
  or (_33673_, _33672_, _33669_);
  and (_33674_, _15413_, _07918_);
  or (_33675_, _33588_, _07231_);
  or (_33676_, _33675_, _33674_);
  and (_33677_, _33676_, _07229_);
  and (_33679_, _33677_, _33673_);
  nor (_33680_, _11204_, _13448_);
  or (_33681_, _33680_, _33588_);
  and (_33682_, _33681_, _06528_);
  or (_33683_, _33682_, _06563_);
  or (_33684_, _33683_, _33679_);
  or (_33685_, _33594_, _07241_);
  and (_33686_, _33685_, _06571_);
  and (_33687_, _33686_, _33684_);
  and (_33688_, _33618_, _06199_);
  or (_33690_, _33688_, _06188_);
  or (_33691_, _33690_, _33687_);
  and (_33692_, _15477_, _07918_);
  or (_33693_, _33588_, _06189_);
  or (_33694_, _33693_, _33692_);
  and (_33695_, _33694_, _01452_);
  and (_33696_, _33695_, _33691_);
  or (_33697_, _33696_, _33587_);
  and (_43910_, _33697_, _43223_);
  and (_33698_, _01456_, \oc8051_golden_model_1.IP [6]);
  and (_33700_, _13448_, \oc8051_golden_model_1.IP [6]);
  nor (_33701_, _08106_, _13448_);
  or (_33702_, _33701_, _33700_);
  or (_33703_, _33702_, _07142_);
  and (_33704_, _15512_, _07918_);
  or (_33705_, _33704_, _33700_);
  or (_33706_, _33705_, _06252_);
  and (_33707_, _07918_, \oc8051_golden_model_1.ACC [6]);
  or (_33708_, _33707_, _33700_);
  and (_33709_, _33708_, _07123_);
  and (_33711_, _07124_, \oc8051_golden_model_1.IP [6]);
  or (_33712_, _33711_, _06251_);
  or (_33713_, _33712_, _33709_);
  and (_33714_, _33713_, _06476_);
  and (_33715_, _33714_, _33706_);
  and (_33716_, _13468_, \oc8051_golden_model_1.IP [6]);
  and (_33717_, _15499_, _08541_);
  or (_33718_, _33717_, _33716_);
  and (_33719_, _33718_, _06475_);
  or (_33720_, _33719_, _06468_);
  or (_33722_, _33720_, _33715_);
  and (_33723_, _33722_, _33703_);
  or (_33724_, _33723_, _06466_);
  or (_33725_, _33708_, _06801_);
  and (_33726_, _33725_, _06484_);
  and (_33727_, _33726_, _33724_);
  and (_33728_, _15497_, _08541_);
  or (_33729_, _33728_, _33716_);
  and (_33730_, _33729_, _06483_);
  or (_33731_, _33730_, _06461_);
  or (_33733_, _33731_, _33727_);
  or (_33734_, _33716_, _15529_);
  and (_33735_, _33734_, _33718_);
  or (_33736_, _33735_, _07164_);
  and (_33737_, _33736_, _06242_);
  and (_33738_, _33737_, _33733_);
  or (_33739_, _33716_, _15545_);
  and (_33740_, _33739_, _06241_);
  and (_33741_, _33740_, _33718_);
  or (_33742_, _33741_, _07187_);
  or (_33744_, _33742_, _33738_);
  or (_33745_, _33702_, _07188_);
  and (_33746_, _33745_, _33744_);
  or (_33747_, _33746_, _07182_);
  and (_33748_, _09067_, _07918_);
  or (_33749_, _33700_, _07183_);
  or (_33750_, _33749_, _33748_);
  and (_33751_, _33750_, _06336_);
  and (_33752_, _33751_, _33747_);
  and (_33753_, _15601_, _07918_);
  or (_33755_, _33753_, _33700_);
  and (_33756_, _33755_, _05968_);
  or (_33757_, _33756_, _06371_);
  or (_33758_, _33757_, _33752_);
  and (_33759_, _15608_, _07918_);
  or (_33760_, _33759_, _33700_);
  or (_33761_, _33760_, _07198_);
  and (_33762_, _33761_, _33758_);
  or (_33763_, _33762_, _06367_);
  and (_33764_, _15618_, _07918_);
  or (_33766_, _33764_, _33700_);
  or (_33767_, _33766_, _07218_);
  and (_33768_, _33767_, _07216_);
  and (_33769_, _33768_, _33763_);
  and (_33770_, _11202_, _07918_);
  or (_33771_, _33770_, _33700_);
  and (_33772_, _33771_, _06533_);
  or (_33773_, _33772_, _33769_);
  and (_33774_, _33773_, _07213_);
  or (_33775_, _33700_, _08109_);
  and (_33777_, _33760_, _06366_);
  and (_33778_, _33777_, _33775_);
  or (_33779_, _33778_, _33774_);
  and (_33780_, _33779_, _07210_);
  and (_33781_, _33708_, _06541_);
  and (_33782_, _33781_, _33775_);
  or (_33783_, _33782_, _06383_);
  or (_33784_, _33783_, _33780_);
  and (_33785_, _15615_, _07918_);
  or (_33786_, _33700_, _07231_);
  or (_33788_, _33786_, _33785_);
  and (_33789_, _33788_, _07229_);
  and (_33790_, _33789_, _33784_);
  nor (_33791_, _11201_, _13448_);
  or (_33792_, _33791_, _33700_);
  and (_33793_, _33792_, _06528_);
  or (_33794_, _33793_, _06563_);
  or (_33795_, _33794_, _33790_);
  or (_33796_, _33705_, _07241_);
  and (_33797_, _33796_, _06571_);
  and (_33799_, _33797_, _33795_);
  and (_33800_, _33729_, _06199_);
  or (_33801_, _33800_, _06188_);
  or (_33802_, _33801_, _33799_);
  and (_33803_, _15676_, _07918_);
  or (_33804_, _33700_, _06189_);
  or (_33805_, _33804_, _33803_);
  and (_33806_, _33805_, _01452_);
  and (_33807_, _33806_, _33802_);
  or (_33808_, _33807_, _33698_);
  and (_43911_, _33808_, _43223_);
  and (_33810_, _01456_, \oc8051_golden_model_1.IE [0]);
  and (_33811_, _07865_, \oc8051_golden_model_1.ACC [0]);
  and (_33812_, _33811_, _08351_);
  and (_33813_, _13551_, \oc8051_golden_model_1.IE [0]);
  or (_33814_, _33813_, _07210_);
  or (_33815_, _33814_, _33812_);
  and (_33816_, _07865_, _07325_);
  or (_33817_, _33816_, _33813_);
  or (_33818_, _33817_, _07188_);
  and (_33820_, _13571_, \oc8051_golden_model_1.IE [0]);
  and (_33821_, _14341_, _08537_);
  or (_33822_, _33821_, _33820_);
  and (_33823_, _33822_, _06475_);
  nor (_33824_, _08351_, _13551_);
  or (_33825_, _33824_, _33813_);
  or (_33826_, _33825_, _06252_);
  or (_33827_, _33811_, _33813_);
  and (_33828_, _33827_, _07123_);
  and (_33829_, _07124_, \oc8051_golden_model_1.IE [0]);
  or (_33831_, _33829_, _06251_);
  or (_33832_, _33831_, _33828_);
  and (_33833_, _33832_, _06476_);
  and (_33834_, _33833_, _33826_);
  or (_33835_, _33834_, _33823_);
  and (_33836_, _33835_, _07142_);
  and (_33837_, _33817_, _06468_);
  or (_33838_, _33837_, _06466_);
  or (_33839_, _33838_, _33836_);
  or (_33840_, _33827_, _06801_);
  and (_33842_, _33840_, _06484_);
  and (_33843_, _33842_, _33839_);
  and (_33844_, _33813_, _06483_);
  or (_33845_, _33844_, _06461_);
  or (_33846_, _33845_, _33843_);
  or (_33847_, _33825_, _07164_);
  and (_33848_, _33847_, _06242_);
  and (_33849_, _33848_, _33846_);
  or (_33850_, _33820_, _14371_);
  and (_33851_, _33850_, _06241_);
  and (_33853_, _33851_, _33822_);
  or (_33854_, _33853_, _07187_);
  or (_33855_, _33854_, _33849_);
  and (_33856_, _33855_, _33818_);
  or (_33857_, _33856_, _07182_);
  and (_33858_, _09342_, _07865_);
  or (_33859_, _33813_, _07183_);
  or (_33860_, _33859_, _33858_);
  and (_33861_, _33860_, _33857_);
  or (_33862_, _33861_, _05968_);
  and (_33864_, _14427_, _07865_);
  or (_33865_, _33813_, _06336_);
  or (_33866_, _33865_, _33864_);
  and (_33867_, _33866_, _07198_);
  and (_33868_, _33867_, _33862_);
  and (_33869_, _07865_, _08908_);
  or (_33870_, _33869_, _33813_);
  and (_33871_, _33870_, _06371_);
  or (_33872_, _33871_, _06367_);
  or (_33873_, _33872_, _33868_);
  and (_33875_, _14442_, _07865_);
  or (_33876_, _33875_, _33813_);
  or (_33877_, _33876_, _07218_);
  and (_33878_, _33877_, _07216_);
  and (_33879_, _33878_, _33873_);
  nor (_33880_, _12526_, _13551_);
  or (_33881_, _33880_, _33813_);
  nor (_33882_, _33812_, _07216_);
  and (_33883_, _33882_, _33881_);
  or (_33884_, _33883_, _33879_);
  and (_33886_, _33884_, _07213_);
  nand (_33887_, _33870_, _06366_);
  nor (_33888_, _33887_, _33824_);
  or (_33889_, _33888_, _06541_);
  or (_33890_, _33889_, _33886_);
  and (_33891_, _33890_, _33815_);
  or (_33892_, _33891_, _06383_);
  and (_33893_, _14325_, _07865_);
  or (_33894_, _33813_, _07231_);
  or (_33895_, _33894_, _33893_);
  and (_33897_, _33895_, _07229_);
  and (_33898_, _33897_, _33892_);
  and (_33899_, _33881_, _06528_);
  or (_33900_, _33899_, _06563_);
  or (_33901_, _33900_, _33898_);
  or (_33902_, _33825_, _07241_);
  and (_33903_, _33902_, _33901_);
  or (_33904_, _33903_, _06199_);
  or (_33905_, _33813_, _06571_);
  and (_33906_, _33905_, _33904_);
  or (_33908_, _33906_, _06188_);
  or (_33909_, _33825_, _06189_);
  and (_33910_, _33909_, _01452_);
  and (_33911_, _33910_, _33908_);
  or (_33912_, _33911_, _33810_);
  and (_43912_, _33912_, _43223_);
  not (_33913_, \oc8051_golden_model_1.IE [1]);
  nor (_33914_, _01452_, _33913_);
  nor (_33915_, _07865_, _33913_);
  nor (_33916_, _11216_, _13551_);
  or (_33918_, _33916_, _33915_);
  or (_33919_, _33918_, _07229_);
  nand (_33920_, _07865_, _07018_);
  or (_33921_, _07865_, \oc8051_golden_model_1.IE [1]);
  and (_33922_, _33921_, _06371_);
  and (_33923_, _33922_, _33920_);
  nor (_33924_, _13551_, _07120_);
  or (_33925_, _33924_, _33915_);
  or (_33926_, _33925_, _07142_);
  and (_33927_, _14503_, _07865_);
  not (_33929_, _33927_);
  and (_33930_, _33929_, _33921_);
  or (_33931_, _33930_, _06252_);
  and (_33932_, _07865_, \oc8051_golden_model_1.ACC [1]);
  or (_33933_, _33932_, _33915_);
  and (_33934_, _33933_, _07123_);
  nor (_33935_, _07123_, _33913_);
  or (_33936_, _33935_, _06251_);
  or (_33937_, _33936_, _33934_);
  and (_33938_, _33937_, _06476_);
  and (_33940_, _33938_, _33931_);
  nor (_33941_, _08537_, _33913_);
  and (_33942_, _14510_, _08537_);
  or (_33943_, _33942_, _33941_);
  and (_33944_, _33943_, _06475_);
  or (_33945_, _33944_, _06468_);
  or (_33946_, _33945_, _33940_);
  and (_33947_, _33946_, _33926_);
  or (_33948_, _33947_, _06466_);
  or (_33949_, _33933_, _06801_);
  and (_33951_, _33949_, _06484_);
  and (_33952_, _33951_, _33948_);
  and (_33953_, _14513_, _08537_);
  or (_33954_, _33953_, _33941_);
  and (_33955_, _33954_, _06483_);
  or (_33956_, _33955_, _06461_);
  or (_33957_, _33956_, _33952_);
  or (_33958_, _33941_, _14509_);
  and (_33959_, _33958_, _33943_);
  or (_33960_, _33959_, _07164_);
  and (_33962_, _33960_, _06242_);
  and (_33963_, _33962_, _33957_);
  or (_33964_, _33941_, _14553_);
  and (_33965_, _33964_, _06241_);
  and (_33966_, _33965_, _33943_);
  or (_33967_, _33966_, _07187_);
  or (_33968_, _33967_, _33963_);
  or (_33969_, _33925_, _07188_);
  and (_33970_, _33969_, _33968_);
  or (_33971_, _33970_, _07182_);
  and (_33973_, _09297_, _07865_);
  or (_33974_, _33915_, _07183_);
  or (_33975_, _33974_, _33973_);
  and (_33976_, _33975_, _06336_);
  and (_33977_, _33976_, _33971_);
  and (_33978_, _14609_, _07865_);
  or (_33979_, _33978_, _33915_);
  and (_33980_, _33979_, _05968_);
  or (_33981_, _33980_, _33977_);
  and (_33982_, _33981_, _07198_);
  or (_33984_, _33982_, _33923_);
  and (_33985_, _33984_, _07218_);
  or (_33986_, _14625_, _13551_);
  and (_33987_, _33921_, _06367_);
  and (_33988_, _33987_, _33986_);
  or (_33989_, _33988_, _06533_);
  or (_33990_, _33989_, _33985_);
  nand (_33991_, _11215_, _07865_);
  and (_33992_, _33991_, _33918_);
  or (_33993_, _33992_, _07216_);
  and (_33995_, _33993_, _07213_);
  and (_33996_, _33995_, _33990_);
  or (_33997_, _14623_, _13551_);
  and (_33998_, _33921_, _06366_);
  and (_33999_, _33998_, _33997_);
  or (_34000_, _33999_, _06541_);
  or (_34001_, _34000_, _33996_);
  nor (_34002_, _33915_, _07210_);
  nand (_34003_, _34002_, _33991_);
  and (_34004_, _34003_, _07231_);
  and (_34006_, _34004_, _34001_);
  or (_34007_, _33920_, _08302_);
  and (_34008_, _33921_, _06383_);
  and (_34009_, _34008_, _34007_);
  or (_34010_, _34009_, _06528_);
  or (_34011_, _34010_, _34006_);
  and (_34012_, _34011_, _33919_);
  or (_34013_, _34012_, _06563_);
  or (_34014_, _33930_, _07241_);
  and (_34015_, _34014_, _06571_);
  and (_34017_, _34015_, _34013_);
  and (_34018_, _33954_, _06199_);
  or (_34019_, _34018_, _06188_);
  or (_34020_, _34019_, _34017_);
  or (_34021_, _33915_, _06189_);
  or (_34022_, _34021_, _33927_);
  and (_34023_, _34022_, _01452_);
  and (_34024_, _34023_, _34020_);
  or (_34025_, _34024_, _33914_);
  and (_43913_, _34025_, _43223_);
  and (_34027_, _01456_, \oc8051_golden_model_1.IE [2]);
  and (_34028_, _13551_, \oc8051_golden_model_1.IE [2]);
  nor (_34029_, _13551_, _07578_);
  or (_34030_, _34029_, _34028_);
  or (_34031_, _34030_, _07188_);
  and (_34032_, _14712_, _07865_);
  or (_34033_, _34032_, _34028_);
  or (_34034_, _34033_, _06252_);
  and (_34035_, _07865_, \oc8051_golden_model_1.ACC [2]);
  or (_34036_, _34035_, _34028_);
  and (_34038_, _34036_, _07123_);
  and (_34039_, _07124_, \oc8051_golden_model_1.IE [2]);
  or (_34040_, _34039_, _06251_);
  or (_34041_, _34040_, _34038_);
  and (_34042_, _34041_, _06476_);
  and (_34043_, _34042_, _34034_);
  and (_34044_, _13571_, \oc8051_golden_model_1.IE [2]);
  and (_34045_, _14702_, _08537_);
  or (_34046_, _34045_, _34044_);
  and (_34047_, _34046_, _06475_);
  or (_34049_, _34047_, _06468_);
  or (_34050_, _34049_, _34043_);
  or (_34051_, _34030_, _07142_);
  and (_34052_, _34051_, _34050_);
  or (_34053_, _34052_, _06466_);
  or (_34054_, _34036_, _06801_);
  and (_34055_, _34054_, _06484_);
  and (_34056_, _34055_, _34053_);
  and (_34057_, _14706_, _08537_);
  or (_34058_, _34057_, _34044_);
  and (_34060_, _34058_, _06483_);
  or (_34061_, _34060_, _06461_);
  or (_34062_, _34061_, _34056_);
  or (_34063_, _34044_, _14739_);
  and (_34064_, _34063_, _34046_);
  or (_34065_, _34064_, _07164_);
  and (_34066_, _34065_, _06242_);
  and (_34067_, _34066_, _34062_);
  or (_34068_, _34044_, _14703_);
  and (_34069_, _34068_, _06241_);
  and (_34070_, _34069_, _34046_);
  or (_34071_, _34070_, _07187_);
  or (_34072_, _34071_, _34067_);
  and (_34073_, _34072_, _34031_);
  or (_34074_, _34073_, _07182_);
  and (_34075_, _09251_, _07865_);
  or (_34076_, _34028_, _07183_);
  or (_34077_, _34076_, _34075_);
  and (_34078_, _34077_, _06336_);
  and (_34079_, _34078_, _34074_);
  and (_34081_, _14808_, _07865_);
  or (_34082_, _34081_, _34028_);
  and (_34083_, _34082_, _05968_);
  or (_34084_, _34083_, _06371_);
  or (_34085_, _34084_, _34079_);
  and (_34086_, _07865_, _08945_);
  or (_34087_, _34086_, _34028_);
  or (_34088_, _34087_, _07198_);
  and (_34089_, _34088_, _34085_);
  or (_34090_, _34089_, _06367_);
  and (_34092_, _14824_, _07865_);
  or (_34093_, _34092_, _34028_);
  or (_34094_, _34093_, _07218_);
  and (_34095_, _34094_, _07216_);
  and (_34096_, _34095_, _34090_);
  and (_34097_, _11214_, _07865_);
  or (_34098_, _34097_, _34028_);
  and (_34099_, _34098_, _06533_);
  or (_34100_, _34099_, _34096_);
  and (_34101_, _34100_, _07213_);
  or (_34103_, _34028_, _08397_);
  and (_34104_, _34087_, _06366_);
  and (_34105_, _34104_, _34103_);
  or (_34106_, _34105_, _34101_);
  and (_34107_, _34106_, _07210_);
  and (_34108_, _34036_, _06541_);
  and (_34109_, _34108_, _34103_);
  or (_34110_, _34109_, _06383_);
  or (_34111_, _34110_, _34107_);
  and (_34112_, _14821_, _07865_);
  or (_34114_, _34028_, _07231_);
  or (_34115_, _34114_, _34112_);
  and (_34116_, _34115_, _07229_);
  and (_34117_, _34116_, _34111_);
  nor (_34118_, _11213_, _13551_);
  or (_34119_, _34118_, _34028_);
  and (_34120_, _34119_, _06528_);
  or (_34121_, _34120_, _06563_);
  or (_34122_, _34121_, _34117_);
  or (_34123_, _34033_, _07241_);
  and (_34125_, _34123_, _06571_);
  and (_34126_, _34125_, _34122_);
  and (_34127_, _34058_, _06199_);
  or (_34128_, _34127_, _06188_);
  or (_34129_, _34128_, _34126_);
  and (_34130_, _14884_, _07865_);
  or (_34131_, _34028_, _06189_);
  or (_34132_, _34131_, _34130_);
  and (_34133_, _34132_, _01452_);
  and (_34134_, _34133_, _34129_);
  or (_34136_, _34134_, _34027_);
  and (_43914_, _34136_, _43223_);
  and (_34137_, _01456_, \oc8051_golden_model_1.IE [3]);
  and (_34138_, _13551_, \oc8051_golden_model_1.IE [3]);
  nor (_34139_, _13551_, _07713_);
  or (_34140_, _34139_, _34138_);
  or (_34141_, _34140_, _07188_);
  or (_34142_, _34140_, _07142_);
  and (_34143_, _14898_, _07865_);
  or (_34144_, _34143_, _34138_);
  or (_34146_, _34144_, _06252_);
  and (_34147_, _07865_, \oc8051_golden_model_1.ACC [3]);
  or (_34148_, _34147_, _34138_);
  and (_34149_, _34148_, _07123_);
  and (_34150_, _07124_, \oc8051_golden_model_1.IE [3]);
  or (_34151_, _34150_, _06251_);
  or (_34152_, _34151_, _34149_);
  and (_34153_, _34152_, _06476_);
  and (_34154_, _34153_, _34146_);
  and (_34155_, _13571_, \oc8051_golden_model_1.IE [3]);
  and (_34157_, _14906_, _08537_);
  or (_34158_, _34157_, _34155_);
  and (_34159_, _34158_, _06475_);
  or (_34160_, _34159_, _06468_);
  or (_34161_, _34160_, _34154_);
  and (_34162_, _34161_, _34142_);
  or (_34163_, _34162_, _06466_);
  or (_34164_, _34148_, _06801_);
  and (_34166_, _34164_, _06484_);
  and (_34168_, _34166_, _34163_);
  and (_34171_, _14904_, _08537_);
  or (_34173_, _34171_, _34155_);
  and (_34175_, _34173_, _06483_);
  or (_34177_, _34175_, _06461_);
  or (_34179_, _34177_, _34168_);
  or (_34181_, _34155_, _14931_);
  and (_34183_, _34181_, _34158_);
  or (_34185_, _34183_, _07164_);
  and (_34186_, _34185_, _06242_);
  and (_34187_, _34186_, _34179_);
  or (_34189_, _34155_, _14947_);
  and (_34190_, _34189_, _06241_);
  and (_34191_, _34190_, _34158_);
  or (_34192_, _34191_, _07187_);
  or (_34193_, _34192_, _34187_);
  and (_34194_, _34193_, _34141_);
  or (_34195_, _34194_, _07182_);
  and (_34196_, _09205_, _07865_);
  or (_34197_, _34138_, _07183_);
  or (_34198_, _34197_, _34196_);
  and (_34200_, _34198_, _06336_);
  and (_34201_, _34200_, _34195_);
  and (_34202_, _15003_, _07865_);
  or (_34203_, _34202_, _34138_);
  and (_34204_, _34203_, _05968_);
  or (_34205_, _34204_, _06371_);
  or (_34206_, _34205_, _34201_);
  and (_34207_, _07865_, _08872_);
  or (_34208_, _34207_, _34138_);
  or (_34209_, _34208_, _07198_);
  and (_34211_, _34209_, _34206_);
  or (_34212_, _34211_, _06367_);
  and (_34213_, _15018_, _07865_);
  or (_34214_, _34213_, _34138_);
  or (_34215_, _34214_, _07218_);
  and (_34216_, _34215_, _07216_);
  and (_34217_, _34216_, _34212_);
  and (_34218_, _12523_, _07865_);
  or (_34219_, _34218_, _34138_);
  and (_34220_, _34219_, _06533_);
  or (_34222_, _34220_, _34217_);
  and (_34223_, _34222_, _07213_);
  or (_34224_, _34138_, _08257_);
  and (_34225_, _34208_, _06366_);
  and (_34226_, _34225_, _34224_);
  or (_34227_, _34226_, _34223_);
  and (_34228_, _34227_, _07210_);
  and (_34229_, _34148_, _06541_);
  and (_34230_, _34229_, _34224_);
  or (_34231_, _34230_, _06383_);
  or (_34233_, _34231_, _34228_);
  and (_34234_, _15015_, _07865_);
  or (_34235_, _34138_, _07231_);
  or (_34236_, _34235_, _34234_);
  and (_34237_, _34236_, _07229_);
  and (_34238_, _34237_, _34233_);
  nor (_34239_, _11211_, _13551_);
  or (_34240_, _34239_, _34138_);
  and (_34241_, _34240_, _06528_);
  or (_34242_, _34241_, _06563_);
  or (_34244_, _34242_, _34238_);
  or (_34245_, _34144_, _07241_);
  and (_34246_, _34245_, _06571_);
  and (_34247_, _34246_, _34244_);
  and (_34248_, _34173_, _06199_);
  or (_34249_, _34248_, _06188_);
  or (_34250_, _34249_, _34247_);
  and (_34251_, _15075_, _07865_);
  or (_34252_, _34138_, _06189_);
  or (_34253_, _34252_, _34251_);
  and (_34255_, _34253_, _01452_);
  and (_34256_, _34255_, _34250_);
  or (_34257_, _34256_, _34137_);
  and (_43915_, _34257_, _43223_);
  and (_34258_, _01456_, \oc8051_golden_model_1.IE [4]);
  and (_34259_, _13551_, \oc8051_golden_model_1.IE [4]);
  nor (_34260_, _08494_, _13551_);
  or (_34261_, _34260_, _34259_);
  or (_34262_, _34261_, _07188_);
  and (_34263_, _13571_, \oc8051_golden_model_1.IE [4]);
  and (_34265_, _15089_, _08537_);
  or (_34266_, _34265_, _34263_);
  and (_34267_, _34266_, _06483_);
  or (_34268_, _34261_, _07142_);
  and (_34269_, _15108_, _07865_);
  or (_34270_, _34269_, _34259_);
  or (_34271_, _34270_, _06252_);
  and (_34272_, _07865_, \oc8051_golden_model_1.ACC [4]);
  or (_34273_, _34272_, _34259_);
  and (_34274_, _34273_, _07123_);
  and (_34276_, _07124_, \oc8051_golden_model_1.IE [4]);
  or (_34277_, _34276_, _06251_);
  or (_34278_, _34277_, _34274_);
  and (_34279_, _34278_, _06476_);
  and (_34280_, _34279_, _34271_);
  and (_34281_, _15091_, _08537_);
  or (_34282_, _34281_, _34263_);
  and (_34283_, _34282_, _06475_);
  or (_34284_, _34283_, _06468_);
  or (_34285_, _34284_, _34280_);
  and (_34287_, _34285_, _34268_);
  or (_34288_, _34287_, _06466_);
  or (_34289_, _34273_, _06801_);
  and (_34290_, _34289_, _06484_);
  and (_34291_, _34290_, _34288_);
  or (_34292_, _34291_, _34267_);
  and (_34293_, _34292_, _07164_);
  and (_34294_, _15126_, _08537_);
  or (_34295_, _34294_, _34263_);
  and (_34296_, _34295_, _06461_);
  or (_34298_, _34296_, _34293_);
  and (_34299_, _34298_, _06242_);
  or (_34300_, _34263_, _15141_);
  and (_34301_, _34300_, _06241_);
  and (_34302_, _34301_, _34282_);
  or (_34303_, _34302_, _07187_);
  or (_34304_, _34303_, _34299_);
  and (_34305_, _34304_, _34262_);
  or (_34306_, _34305_, _07182_);
  and (_34307_, _09159_, _07865_);
  or (_34309_, _34259_, _07183_);
  or (_34310_, _34309_, _34307_);
  and (_34311_, _34310_, _06336_);
  and (_34312_, _34311_, _34306_);
  and (_34313_, _15198_, _07865_);
  or (_34314_, _34313_, _34259_);
  and (_34315_, _34314_, _05968_);
  or (_34316_, _34315_, _06371_);
  or (_34317_, _34316_, _34312_);
  and (_34318_, _08892_, _07865_);
  or (_34320_, _34318_, _34259_);
  or (_34321_, _34320_, _07198_);
  and (_34322_, _34321_, _34317_);
  or (_34323_, _34322_, _06367_);
  and (_34324_, _15214_, _07865_);
  or (_34325_, _34324_, _34259_);
  or (_34326_, _34325_, _07218_);
  and (_34327_, _34326_, _07216_);
  and (_34328_, _34327_, _34323_);
  and (_34329_, _11209_, _07865_);
  or (_34331_, _34329_, _34259_);
  and (_34332_, _34331_, _06533_);
  or (_34333_, _34332_, _34328_);
  and (_34334_, _34333_, _07213_);
  or (_34335_, _34259_, _08497_);
  and (_34336_, _34320_, _06366_);
  and (_34337_, _34336_, _34335_);
  or (_34338_, _34337_, _34334_);
  and (_34339_, _34338_, _07210_);
  and (_34340_, _34273_, _06541_);
  and (_34342_, _34340_, _34335_);
  or (_34343_, _34342_, _06383_);
  or (_34344_, _34343_, _34339_);
  and (_34345_, _15211_, _07865_);
  or (_34346_, _34259_, _07231_);
  or (_34347_, _34346_, _34345_);
  and (_34348_, _34347_, _07229_);
  and (_34349_, _34348_, _34344_);
  nor (_34350_, _11208_, _13551_);
  or (_34351_, _34350_, _34259_);
  and (_34353_, _34351_, _06528_);
  or (_34354_, _34353_, _06563_);
  or (_34355_, _34354_, _34349_);
  or (_34356_, _34270_, _07241_);
  and (_34357_, _34356_, _06571_);
  and (_34358_, _34357_, _34355_);
  and (_34359_, _34266_, _06199_);
  or (_34360_, _34359_, _06188_);
  or (_34361_, _34360_, _34358_);
  and (_34362_, _15280_, _07865_);
  or (_34364_, _34259_, _06189_);
  or (_34365_, _34364_, _34362_);
  and (_34366_, _34365_, _01452_);
  and (_34367_, _34366_, _34361_);
  or (_34368_, _34367_, _34258_);
  and (_43916_, _34368_, _43223_);
  and (_34369_, _01456_, \oc8051_golden_model_1.IE [5]);
  and (_34370_, _13551_, \oc8051_golden_model_1.IE [5]);
  nor (_34371_, _08209_, _13551_);
  or (_34372_, _34371_, _34370_);
  or (_34374_, _34372_, _07142_);
  and (_34375_, _15311_, _07865_);
  or (_34376_, _34375_, _34370_);
  or (_34377_, _34376_, _06252_);
  and (_34378_, _07865_, \oc8051_golden_model_1.ACC [5]);
  or (_34379_, _34378_, _34370_);
  and (_34380_, _34379_, _07123_);
  and (_34381_, _07124_, \oc8051_golden_model_1.IE [5]);
  or (_34382_, _34381_, _06251_);
  or (_34383_, _34382_, _34380_);
  and (_34385_, _34383_, _06476_);
  and (_34386_, _34385_, _34377_);
  and (_34387_, _13571_, \oc8051_golden_model_1.IE [5]);
  and (_34388_, _15296_, _08537_);
  or (_34389_, _34388_, _34387_);
  and (_34390_, _34389_, _06475_);
  or (_34391_, _34390_, _06468_);
  or (_34392_, _34391_, _34386_);
  and (_34393_, _34392_, _34374_);
  or (_34394_, _34393_, _06466_);
  or (_34396_, _34379_, _06801_);
  and (_34397_, _34396_, _06484_);
  and (_34398_, _34397_, _34394_);
  and (_34399_, _15294_, _08537_);
  or (_34400_, _34399_, _34387_);
  and (_34401_, _34400_, _06483_);
  or (_34402_, _34401_, _06461_);
  or (_34403_, _34402_, _34398_);
  or (_34404_, _34387_, _15328_);
  and (_34405_, _34404_, _34389_);
  or (_34407_, _34405_, _07164_);
  and (_34408_, _34407_, _06242_);
  and (_34409_, _34408_, _34403_);
  or (_34410_, _34387_, _15344_);
  and (_34411_, _34410_, _06241_);
  and (_34412_, _34411_, _34389_);
  or (_34413_, _34412_, _07187_);
  or (_34414_, _34413_, _34409_);
  or (_34415_, _34372_, _07188_);
  and (_34416_, _34415_, _34414_);
  or (_34418_, _34416_, _07182_);
  and (_34419_, _09113_, _07865_);
  or (_34420_, _34370_, _07183_);
  or (_34421_, _34420_, _34419_);
  and (_34422_, _34421_, _06336_);
  and (_34423_, _34422_, _34418_);
  and (_34424_, _15400_, _07865_);
  or (_34425_, _34424_, _34370_);
  and (_34426_, _34425_, _05968_);
  or (_34427_, _34426_, _06371_);
  or (_34429_, _34427_, _34423_);
  and (_34430_, _08888_, _07865_);
  or (_34431_, _34430_, _34370_);
  or (_34432_, _34431_, _07198_);
  and (_34433_, _34432_, _34429_);
  or (_34434_, _34433_, _06367_);
  and (_34435_, _15416_, _07865_);
  or (_34436_, _34435_, _34370_);
  or (_34437_, _34436_, _07218_);
  and (_34438_, _34437_, _07216_);
  and (_34440_, _34438_, _34434_);
  and (_34441_, _11205_, _07865_);
  or (_34442_, _34441_, _34370_);
  and (_34443_, _34442_, _06533_);
  or (_34444_, _34443_, _34440_);
  and (_34445_, _34444_, _07213_);
  or (_34446_, _34370_, _08212_);
  and (_34447_, _34431_, _06366_);
  and (_34448_, _34447_, _34446_);
  or (_34449_, _34448_, _34445_);
  and (_34451_, _34449_, _07210_);
  and (_34452_, _34379_, _06541_);
  and (_34453_, _34452_, _34446_);
  or (_34454_, _34453_, _06383_);
  or (_34455_, _34454_, _34451_);
  and (_34456_, _15413_, _07865_);
  or (_34457_, _34370_, _07231_);
  or (_34458_, _34457_, _34456_);
  and (_34459_, _34458_, _07229_);
  and (_34460_, _34459_, _34455_);
  nor (_34462_, _11204_, _13551_);
  or (_34463_, _34462_, _34370_);
  and (_34464_, _34463_, _06528_);
  or (_34465_, _34464_, _06563_);
  or (_34466_, _34465_, _34460_);
  or (_34467_, _34376_, _07241_);
  and (_34468_, _34467_, _06571_);
  and (_34469_, _34468_, _34466_);
  and (_34470_, _34400_, _06199_);
  or (_34471_, _34470_, _06188_);
  or (_34473_, _34471_, _34469_);
  and (_34474_, _15477_, _07865_);
  or (_34475_, _34370_, _06189_);
  or (_34476_, _34475_, _34474_);
  and (_34477_, _34476_, _01452_);
  and (_34478_, _34477_, _34473_);
  or (_34479_, _34478_, _34369_);
  and (_43917_, _34479_, _43223_);
  and (_34480_, _01456_, \oc8051_golden_model_1.IE [6]);
  and (_34481_, _13551_, \oc8051_golden_model_1.IE [6]);
  nor (_34483_, _08106_, _13551_);
  or (_34484_, _34483_, _34481_);
  or (_34485_, _34484_, _07142_);
  and (_34486_, _15512_, _07865_);
  or (_34487_, _34486_, _34481_);
  or (_34488_, _34487_, _06252_);
  and (_34489_, _07865_, \oc8051_golden_model_1.ACC [6]);
  or (_34490_, _34489_, _34481_);
  and (_34491_, _34490_, _07123_);
  and (_34492_, _07124_, \oc8051_golden_model_1.IE [6]);
  or (_34494_, _34492_, _06251_);
  or (_34495_, _34494_, _34491_);
  and (_34496_, _34495_, _06476_);
  and (_34497_, _34496_, _34488_);
  and (_34498_, _13571_, \oc8051_golden_model_1.IE [6]);
  and (_34499_, _15499_, _08537_);
  or (_34500_, _34499_, _34498_);
  and (_34501_, _34500_, _06475_);
  or (_34502_, _34501_, _06468_);
  or (_34503_, _34502_, _34497_);
  and (_34505_, _34503_, _34485_);
  or (_34506_, _34505_, _06466_);
  or (_34507_, _34490_, _06801_);
  and (_34508_, _34507_, _06484_);
  and (_34509_, _34508_, _34506_);
  and (_34510_, _15497_, _08537_);
  or (_34511_, _34510_, _34498_);
  and (_34512_, _34511_, _06483_);
  or (_34513_, _34512_, _06461_);
  or (_34514_, _34513_, _34509_);
  or (_34516_, _34498_, _15529_);
  and (_34517_, _34516_, _34500_);
  or (_34518_, _34517_, _07164_);
  and (_34519_, _34518_, _06242_);
  and (_34520_, _34519_, _34514_);
  or (_34521_, _34498_, _15545_);
  and (_34522_, _34521_, _06241_);
  and (_34523_, _34522_, _34500_);
  or (_34524_, _34523_, _07187_);
  or (_34525_, _34524_, _34520_);
  or (_34527_, _34484_, _07188_);
  and (_34528_, _34527_, _34525_);
  or (_34529_, _34528_, _07182_);
  and (_34530_, _09067_, _07865_);
  or (_34531_, _34481_, _07183_);
  or (_34532_, _34531_, _34530_);
  and (_34533_, _34532_, _06336_);
  and (_34534_, _34533_, _34529_);
  and (_34535_, _15601_, _07865_);
  or (_34536_, _34535_, _34481_);
  and (_34538_, _34536_, _05968_);
  or (_34539_, _34538_, _06371_);
  or (_34540_, _34539_, _34534_);
  and (_34541_, _15608_, _07865_);
  or (_34542_, _34541_, _34481_);
  or (_34543_, _34542_, _07198_);
  and (_34544_, _34543_, _34540_);
  or (_34545_, _34544_, _06367_);
  and (_34546_, _15618_, _07865_);
  or (_34547_, _34546_, _34481_);
  or (_34549_, _34547_, _07218_);
  and (_34550_, _34549_, _07216_);
  and (_34551_, _34550_, _34545_);
  and (_34552_, _11202_, _07865_);
  or (_34553_, _34552_, _34481_);
  and (_34554_, _34553_, _06533_);
  or (_34555_, _34554_, _34551_);
  and (_34556_, _34555_, _07213_);
  or (_34557_, _34481_, _08109_);
  and (_34558_, _34542_, _06366_);
  and (_34560_, _34558_, _34557_);
  or (_34561_, _34560_, _34556_);
  and (_34562_, _34561_, _07210_);
  and (_34563_, _34490_, _06541_);
  and (_34564_, _34563_, _34557_);
  or (_34565_, _34564_, _06383_);
  or (_34566_, _34565_, _34562_);
  and (_34567_, _15615_, _07865_);
  or (_34568_, _34481_, _07231_);
  or (_34569_, _34568_, _34567_);
  and (_34571_, _34569_, _07229_);
  and (_34572_, _34571_, _34566_);
  nor (_34573_, _11201_, _13551_);
  or (_34574_, _34573_, _34481_);
  and (_34575_, _34574_, _06528_);
  or (_34576_, _34575_, _06563_);
  or (_34577_, _34576_, _34572_);
  or (_34578_, _34487_, _07241_);
  and (_34579_, _34578_, _06571_);
  and (_34580_, _34579_, _34577_);
  and (_34582_, _34511_, _06199_);
  or (_34583_, _34582_, _06188_);
  or (_34584_, _34583_, _34580_);
  and (_34585_, _15676_, _07865_);
  or (_34586_, _34481_, _06189_);
  or (_34587_, _34586_, _34585_);
  and (_34588_, _34587_, _01452_);
  and (_34589_, _34588_, _34584_);
  or (_34590_, _34589_, _34480_);
  and (_43918_, _34590_, _43223_);
  not (_34592_, \oc8051_golden_model_1.SCON [0]);
  nor (_34593_, _01452_, _34592_);
  nand (_34594_, _11218_, _07943_);
  nor (_34595_, _07943_, _34592_);
  nor (_34596_, _34595_, _07210_);
  nand (_34597_, _34596_, _34594_);
  and (_34598_, _07943_, _07325_);
  or (_34599_, _34598_, _34595_);
  or (_34600_, _34599_, _07188_);
  nor (_34601_, _08533_, _34592_);
  and (_34603_, _14341_, _08533_);
  or (_34604_, _34603_, _34601_);
  and (_34605_, _34604_, _06475_);
  nor (_34606_, _08351_, _13660_);
  or (_34607_, _34606_, _34595_);
  or (_34608_, _34607_, _06252_);
  and (_34609_, _07943_, \oc8051_golden_model_1.ACC [0]);
  or (_34610_, _34609_, _34595_);
  and (_34611_, _34610_, _07123_);
  nor (_34612_, _07123_, _34592_);
  or (_34614_, _34612_, _06251_);
  or (_34615_, _34614_, _34611_);
  and (_34616_, _34615_, _06476_);
  and (_34617_, _34616_, _34608_);
  or (_34618_, _34617_, _34605_);
  and (_34619_, _34618_, _07142_);
  and (_34620_, _34599_, _06468_);
  or (_34621_, _34620_, _06466_);
  or (_34622_, _34621_, _34619_);
  or (_34623_, _34610_, _06801_);
  and (_34625_, _34623_, _06484_);
  and (_34626_, _34625_, _34622_);
  and (_34627_, _34595_, _06483_);
  or (_34628_, _34627_, _06461_);
  or (_34629_, _34628_, _34626_);
  or (_34630_, _34607_, _07164_);
  and (_34631_, _34630_, _06242_);
  and (_34632_, _34631_, _34629_);
  or (_34633_, _34601_, _14371_);
  and (_34634_, _34633_, _06241_);
  and (_34636_, _34634_, _34604_);
  or (_34637_, _34636_, _07187_);
  or (_34638_, _34637_, _34632_);
  and (_34639_, _34638_, _34600_);
  or (_34640_, _34639_, _07182_);
  and (_34641_, _09342_, _07943_);
  or (_34642_, _34595_, _07183_);
  or (_34643_, _34642_, _34641_);
  and (_34644_, _34643_, _34640_);
  or (_34645_, _34644_, _05968_);
  and (_34647_, _14427_, _07943_);
  or (_34648_, _34595_, _06336_);
  or (_34649_, _34648_, _34647_);
  and (_34650_, _34649_, _07198_);
  and (_34651_, _34650_, _34645_);
  and (_34652_, _07943_, _08908_);
  or (_34653_, _34652_, _34595_);
  and (_34654_, _34653_, _06371_);
  or (_34655_, _34654_, _06367_);
  or (_34656_, _34655_, _34651_);
  and (_34658_, _14442_, _07943_);
  or (_34659_, _34658_, _34595_);
  or (_34660_, _34659_, _07218_);
  and (_34661_, _34660_, _07216_);
  and (_34662_, _34661_, _34656_);
  nor (_34663_, _12526_, _13660_);
  or (_34664_, _34663_, _34595_);
  and (_34665_, _34594_, _06533_);
  and (_34666_, _34665_, _34664_);
  or (_34667_, _34666_, _34662_);
  and (_34669_, _34667_, _07213_);
  nand (_34670_, _34653_, _06366_);
  nor (_34671_, _34670_, _34606_);
  or (_34672_, _34671_, _06541_);
  or (_34673_, _34672_, _34669_);
  and (_34674_, _34673_, _34597_);
  or (_34675_, _34674_, _06383_);
  and (_34676_, _14325_, _07943_);
  or (_34677_, _34676_, _34595_);
  or (_34678_, _34677_, _07231_);
  and (_34680_, _34678_, _07229_);
  and (_34681_, _34680_, _34675_);
  and (_34682_, _34664_, _06528_);
  or (_34683_, _34682_, _06563_);
  or (_34684_, _34683_, _34681_);
  or (_34685_, _34607_, _07241_);
  and (_34686_, _34685_, _34684_);
  or (_34687_, _34686_, _06199_);
  or (_34688_, _34595_, _06571_);
  and (_34689_, _34688_, _34687_);
  or (_34691_, _34689_, _06188_);
  or (_34692_, _34607_, _06189_);
  and (_34693_, _34692_, _01452_);
  and (_34694_, _34693_, _34691_);
  or (_34695_, _34694_, _34593_);
  and (_43920_, _34695_, _43223_);
  not (_34696_, \oc8051_golden_model_1.SCON [1]);
  nor (_34697_, _01452_, _34696_);
  nor (_34698_, _07943_, _34696_);
  nor (_34699_, _11216_, _13660_);
  or (_34701_, _34699_, _34698_);
  or (_34702_, _34701_, _07229_);
  nand (_34703_, _07943_, _07018_);
  or (_34704_, _07943_, \oc8051_golden_model_1.SCON [1]);
  and (_34705_, _34704_, _06371_);
  and (_34706_, _34705_, _34703_);
  nor (_34707_, _13660_, _07120_);
  or (_34708_, _34707_, _34698_);
  or (_34709_, _34708_, _07142_);
  and (_34710_, _14503_, _07943_);
  not (_34712_, _34710_);
  and (_34713_, _34712_, _34704_);
  or (_34714_, _34713_, _06252_);
  and (_34715_, _07943_, \oc8051_golden_model_1.ACC [1]);
  or (_34716_, _34715_, _34698_);
  and (_34717_, _34716_, _07123_);
  nor (_34718_, _07123_, _34696_);
  or (_34719_, _34718_, _06251_);
  or (_34720_, _34719_, _34717_);
  and (_34721_, _34720_, _06476_);
  and (_34723_, _34721_, _34714_);
  nor (_34724_, _08533_, _34696_);
  and (_34725_, _14510_, _08533_);
  or (_34726_, _34725_, _34724_);
  and (_34727_, _34726_, _06475_);
  or (_34728_, _34727_, _06468_);
  or (_34729_, _34728_, _34723_);
  and (_34730_, _34729_, _34709_);
  or (_34731_, _34730_, _06466_);
  or (_34732_, _34716_, _06801_);
  and (_34734_, _34732_, _06484_);
  and (_34735_, _34734_, _34731_);
  and (_34736_, _14513_, _08533_);
  or (_34737_, _34736_, _34724_);
  and (_34738_, _34737_, _06483_);
  or (_34739_, _34738_, _06461_);
  or (_34740_, _34739_, _34735_);
  or (_34741_, _34724_, _14509_);
  and (_34742_, _34741_, _34726_);
  or (_34743_, _34742_, _07164_);
  and (_34745_, _34743_, _06242_);
  and (_34746_, _34745_, _34740_);
  or (_34747_, _34724_, _14553_);
  and (_34748_, _34747_, _06241_);
  and (_34749_, _34748_, _34726_);
  or (_34750_, _34749_, _07187_);
  or (_34751_, _34750_, _34746_);
  or (_34752_, _34708_, _07188_);
  and (_34753_, _34752_, _34751_);
  or (_34754_, _34753_, _07182_);
  and (_34756_, _09297_, _07943_);
  or (_34757_, _34698_, _07183_);
  or (_34758_, _34757_, _34756_);
  and (_34759_, _34758_, _06336_);
  and (_34760_, _34759_, _34754_);
  and (_34761_, _14609_, _07943_);
  or (_34762_, _34761_, _34698_);
  and (_34763_, _34762_, _05968_);
  or (_34764_, _34763_, _34760_);
  and (_34765_, _34764_, _07198_);
  or (_34767_, _34765_, _34706_);
  and (_34768_, _34767_, _07218_);
  or (_34769_, _14625_, _13660_);
  and (_34770_, _34704_, _06367_);
  and (_34771_, _34770_, _34769_);
  or (_34772_, _34771_, _06533_);
  or (_34773_, _34772_, _34768_);
  nand (_34774_, _11215_, _07943_);
  and (_34775_, _34774_, _34701_);
  or (_34776_, _34775_, _07216_);
  and (_34778_, _34776_, _07213_);
  and (_34779_, _34778_, _34773_);
  or (_34780_, _14623_, _13660_);
  and (_34781_, _34704_, _06366_);
  and (_34782_, _34781_, _34780_);
  or (_34783_, _34782_, _06541_);
  or (_34784_, _34783_, _34779_);
  nor (_34785_, _34698_, _07210_);
  nand (_34786_, _34785_, _34774_);
  and (_34787_, _34786_, _07231_);
  and (_34789_, _34787_, _34784_);
  or (_34790_, _34703_, _08302_);
  and (_34791_, _34704_, _06383_);
  and (_34792_, _34791_, _34790_);
  or (_34793_, _34792_, _06528_);
  or (_34794_, _34793_, _34789_);
  and (_34795_, _34794_, _34702_);
  or (_34796_, _34795_, _06563_);
  or (_34797_, _34713_, _07241_);
  and (_34798_, _34797_, _06571_);
  and (_34799_, _34798_, _34796_);
  and (_34800_, _34737_, _06199_);
  or (_34801_, _34800_, _06188_);
  or (_34802_, _34801_, _34799_);
  or (_34803_, _34698_, _06189_);
  or (_34804_, _34803_, _34710_);
  and (_34805_, _34804_, _01452_);
  and (_34806_, _34805_, _34802_);
  or (_34807_, _34806_, _34697_);
  and (_43921_, _34807_, _43223_);
  and (_34809_, _01456_, \oc8051_golden_model_1.SCON [2]);
  and (_34810_, _13660_, \oc8051_golden_model_1.SCON [2]);
  nor (_34811_, _13660_, _07578_);
  or (_34812_, _34811_, _34810_);
  or (_34813_, _34812_, _07188_);
  and (_34814_, _14712_, _07943_);
  or (_34815_, _34814_, _34810_);
  or (_34816_, _34815_, _06252_);
  and (_34817_, _07943_, \oc8051_golden_model_1.ACC [2]);
  or (_34818_, _34817_, _34810_);
  and (_34820_, _34818_, _07123_);
  and (_34821_, _07124_, \oc8051_golden_model_1.SCON [2]);
  or (_34822_, _34821_, _06251_);
  or (_34823_, _34822_, _34820_);
  and (_34824_, _34823_, _06476_);
  and (_34825_, _34824_, _34816_);
  and (_34826_, _13682_, \oc8051_golden_model_1.SCON [2]);
  and (_34827_, _14702_, _08533_);
  or (_34828_, _34827_, _34826_);
  and (_34829_, _34828_, _06475_);
  or (_34831_, _34829_, _06468_);
  or (_34832_, _34831_, _34825_);
  or (_34833_, _34812_, _07142_);
  and (_34834_, _34833_, _34832_);
  or (_34835_, _34834_, _06466_);
  or (_34836_, _34818_, _06801_);
  and (_34837_, _34836_, _06484_);
  and (_34838_, _34837_, _34835_);
  and (_34839_, _14706_, _08533_);
  or (_34840_, _34839_, _34826_);
  and (_34842_, _34840_, _06483_);
  or (_34843_, _34842_, _06461_);
  or (_34844_, _34843_, _34838_);
  or (_34845_, _34826_, _14739_);
  and (_34846_, _34845_, _34828_);
  or (_34847_, _34846_, _07164_);
  and (_34848_, _34847_, _06242_);
  and (_34849_, _34848_, _34844_);
  or (_34850_, _34826_, _14703_);
  and (_34851_, _34850_, _06241_);
  and (_34853_, _34851_, _34828_);
  or (_34854_, _34853_, _07187_);
  or (_34855_, _34854_, _34849_);
  and (_34856_, _34855_, _34813_);
  or (_34857_, _34856_, _07182_);
  and (_34858_, _09251_, _07943_);
  or (_34859_, _34810_, _07183_);
  or (_34860_, _34859_, _34858_);
  and (_34861_, _34860_, _06336_);
  and (_34862_, _34861_, _34857_);
  and (_34864_, _14808_, _07943_);
  or (_34865_, _34864_, _34810_);
  and (_34866_, _34865_, _05968_);
  or (_34867_, _34866_, _06371_);
  or (_34868_, _34867_, _34862_);
  and (_34869_, _07943_, _08945_);
  or (_34870_, _34869_, _34810_);
  or (_34871_, _34870_, _07198_);
  and (_34872_, _34871_, _34868_);
  or (_34873_, _34872_, _06367_);
  and (_34875_, _14824_, _07943_);
  or (_34876_, _34875_, _34810_);
  or (_34877_, _34876_, _07218_);
  and (_34878_, _34877_, _07216_);
  and (_34879_, _34878_, _34873_);
  and (_34880_, _11214_, _07943_);
  or (_34881_, _34880_, _34810_);
  and (_34882_, _34881_, _06533_);
  or (_34883_, _34882_, _34879_);
  and (_34884_, _34883_, _07213_);
  or (_34886_, _34810_, _08397_);
  and (_34887_, _34870_, _06366_);
  and (_34888_, _34887_, _34886_);
  or (_34889_, _34888_, _34884_);
  and (_34890_, _34889_, _07210_);
  and (_34891_, _34818_, _06541_);
  and (_34892_, _34891_, _34886_);
  or (_34893_, _34892_, _06383_);
  or (_34894_, _34893_, _34890_);
  and (_34895_, _14821_, _07943_);
  or (_34897_, _34810_, _07231_);
  or (_34898_, _34897_, _34895_);
  and (_34899_, _34898_, _07229_);
  and (_34900_, _34899_, _34894_);
  nor (_34901_, _11213_, _13660_);
  or (_34902_, _34901_, _34810_);
  and (_34903_, _34902_, _06528_);
  or (_34904_, _34903_, _06563_);
  or (_34905_, _34904_, _34900_);
  or (_34906_, _34815_, _07241_);
  and (_34908_, _34906_, _06571_);
  and (_34909_, _34908_, _34905_);
  and (_34910_, _34840_, _06199_);
  or (_34911_, _34910_, _06188_);
  or (_34912_, _34911_, _34909_);
  and (_34913_, _14884_, _07943_);
  or (_34914_, _34810_, _06189_);
  or (_34915_, _34914_, _34913_);
  and (_34916_, _34915_, _01452_);
  and (_34917_, _34916_, _34912_);
  or (_34919_, _34917_, _34809_);
  and (_43922_, _34919_, _43223_);
  and (_34920_, _01456_, \oc8051_golden_model_1.SCON [3]);
  and (_34921_, _13660_, \oc8051_golden_model_1.SCON [3]);
  nor (_34922_, _13660_, _07713_);
  or (_34923_, _34922_, _34921_);
  or (_34924_, _34923_, _07188_);
  or (_34925_, _34923_, _07142_);
  and (_34926_, _14898_, _07943_);
  or (_34927_, _34926_, _34921_);
  or (_34929_, _34927_, _06252_);
  and (_34930_, _07943_, \oc8051_golden_model_1.ACC [3]);
  or (_34931_, _34930_, _34921_);
  and (_34932_, _34931_, _07123_);
  and (_34933_, _07124_, \oc8051_golden_model_1.SCON [3]);
  or (_34934_, _34933_, _06251_);
  or (_34935_, _34934_, _34932_);
  and (_34936_, _34935_, _06476_);
  and (_34937_, _34936_, _34929_);
  and (_34938_, _13682_, \oc8051_golden_model_1.SCON [3]);
  and (_34940_, _14906_, _08533_);
  or (_34941_, _34940_, _34938_);
  and (_34942_, _34941_, _06475_);
  or (_34943_, _34942_, _06468_);
  or (_34944_, _34943_, _34937_);
  and (_34945_, _34944_, _34925_);
  or (_34946_, _34945_, _06466_);
  or (_34947_, _34931_, _06801_);
  and (_34948_, _34947_, _06484_);
  and (_34949_, _34948_, _34946_);
  and (_34951_, _14904_, _08533_);
  or (_34952_, _34951_, _34938_);
  and (_34953_, _34952_, _06483_);
  or (_34954_, _34953_, _06461_);
  or (_34955_, _34954_, _34949_);
  or (_34956_, _34938_, _14931_);
  and (_34957_, _34956_, _34941_);
  or (_34958_, _34957_, _07164_);
  and (_34959_, _34958_, _06242_);
  and (_34960_, _34959_, _34955_);
  or (_34962_, _34938_, _14947_);
  and (_34963_, _34962_, _06241_);
  and (_34964_, _34963_, _34941_);
  or (_34965_, _34964_, _07187_);
  or (_34966_, _34965_, _34960_);
  and (_34967_, _34966_, _34924_);
  or (_34968_, _34967_, _07182_);
  and (_34969_, _09205_, _07943_);
  or (_34970_, _34921_, _07183_);
  or (_34971_, _34970_, _34969_);
  and (_34973_, _34971_, _06336_);
  and (_34974_, _34973_, _34968_);
  and (_34975_, _15003_, _07943_);
  or (_34976_, _34975_, _34921_);
  and (_34977_, _34976_, _05968_);
  or (_34978_, _34977_, _06371_);
  or (_34979_, _34978_, _34974_);
  and (_34980_, _07943_, _08872_);
  or (_34981_, _34980_, _34921_);
  or (_34982_, _34981_, _07198_);
  and (_34984_, _34982_, _34979_);
  or (_34985_, _34984_, _06367_);
  and (_34986_, _15018_, _07943_);
  or (_34987_, _34986_, _34921_);
  or (_34988_, _34987_, _07218_);
  and (_34989_, _34988_, _07216_);
  and (_34990_, _34989_, _34985_);
  and (_34991_, _12523_, _07943_);
  or (_34992_, _34991_, _34921_);
  and (_34993_, _34992_, _06533_);
  or (_34995_, _34993_, _34990_);
  and (_34996_, _34995_, _07213_);
  or (_34997_, _34921_, _08257_);
  and (_34998_, _34981_, _06366_);
  and (_34999_, _34998_, _34997_);
  or (_35000_, _34999_, _34996_);
  and (_35001_, _35000_, _07210_);
  and (_35002_, _34931_, _06541_);
  and (_35003_, _35002_, _34997_);
  or (_35004_, _35003_, _06383_);
  or (_35006_, _35004_, _35001_);
  and (_35007_, _15015_, _07943_);
  or (_35008_, _34921_, _07231_);
  or (_35009_, _35008_, _35007_);
  and (_35010_, _35009_, _07229_);
  and (_35011_, _35010_, _35006_);
  nor (_35012_, _11211_, _13660_);
  or (_35013_, _35012_, _34921_);
  and (_35014_, _35013_, _06528_);
  or (_35015_, _35014_, _06563_);
  or (_35017_, _35015_, _35011_);
  or (_35018_, _34927_, _07241_);
  and (_35019_, _35018_, _06571_);
  and (_35020_, _35019_, _35017_);
  and (_35021_, _34952_, _06199_);
  or (_35022_, _35021_, _06188_);
  or (_35023_, _35022_, _35020_);
  and (_35024_, _15075_, _07943_);
  or (_35025_, _34921_, _06189_);
  or (_35026_, _35025_, _35024_);
  and (_35028_, _35026_, _01452_);
  and (_35029_, _35028_, _35023_);
  or (_35030_, _35029_, _34920_);
  and (_43923_, _35030_, _43223_);
  and (_35031_, _01456_, \oc8051_golden_model_1.SCON [4]);
  and (_35032_, _13660_, \oc8051_golden_model_1.SCON [4]);
  nor (_35033_, _08494_, _13660_);
  or (_35034_, _35033_, _35032_);
  or (_35035_, _35034_, _07188_);
  and (_35036_, _13682_, \oc8051_golden_model_1.SCON [4]);
  and (_35038_, _15089_, _08533_);
  or (_35039_, _35038_, _35036_);
  and (_35040_, _35039_, _06483_);
  or (_35041_, _35034_, _07142_);
  and (_35042_, _15108_, _07943_);
  or (_35043_, _35042_, _35032_);
  or (_35044_, _35043_, _06252_);
  and (_35045_, _07943_, \oc8051_golden_model_1.ACC [4]);
  or (_35046_, _35045_, _35032_);
  and (_35047_, _35046_, _07123_);
  and (_35049_, _07124_, \oc8051_golden_model_1.SCON [4]);
  or (_35050_, _35049_, _06251_);
  or (_35051_, _35050_, _35047_);
  and (_35052_, _35051_, _06476_);
  and (_35053_, _35052_, _35044_);
  and (_35054_, _15091_, _08533_);
  or (_35055_, _35054_, _35036_);
  and (_35056_, _35055_, _06475_);
  or (_35057_, _35056_, _06468_);
  or (_35058_, _35057_, _35053_);
  and (_35060_, _35058_, _35041_);
  or (_35061_, _35060_, _06466_);
  or (_35062_, _35046_, _06801_);
  and (_35063_, _35062_, _06484_);
  and (_35064_, _35063_, _35061_);
  or (_35065_, _35064_, _35040_);
  and (_35066_, _35065_, _07164_);
  or (_35067_, _35036_, _15125_);
  and (_35068_, _35067_, _06461_);
  and (_35069_, _35068_, _35055_);
  or (_35071_, _35069_, _35066_);
  and (_35072_, _35071_, _06242_);
  or (_35073_, _35036_, _15141_);
  and (_35074_, _35073_, _06241_);
  and (_35075_, _35074_, _35055_);
  or (_35076_, _35075_, _07187_);
  or (_35077_, _35076_, _35072_);
  and (_35078_, _35077_, _35035_);
  or (_35079_, _35078_, _07182_);
  and (_35080_, _09159_, _07943_);
  or (_35082_, _35032_, _07183_);
  or (_35083_, _35082_, _35080_);
  and (_35084_, _35083_, _06336_);
  and (_35085_, _35084_, _35079_);
  and (_35086_, _15198_, _07943_);
  or (_35087_, _35086_, _35032_);
  and (_35088_, _35087_, _05968_);
  or (_35089_, _35088_, _06371_);
  or (_35090_, _35089_, _35085_);
  and (_35091_, _08892_, _07943_);
  or (_35093_, _35091_, _35032_);
  or (_35094_, _35093_, _07198_);
  and (_35095_, _35094_, _35090_);
  or (_35096_, _35095_, _06367_);
  and (_35097_, _15214_, _07943_);
  or (_35098_, _35097_, _35032_);
  or (_35099_, _35098_, _07218_);
  and (_35100_, _35099_, _07216_);
  and (_35101_, _35100_, _35096_);
  and (_35102_, _11209_, _07943_);
  or (_35104_, _35102_, _35032_);
  and (_35105_, _35104_, _06533_);
  or (_35106_, _35105_, _35101_);
  and (_35107_, _35106_, _07213_);
  or (_35108_, _35032_, _08497_);
  and (_35109_, _35093_, _06366_);
  and (_35110_, _35109_, _35108_);
  or (_35111_, _35110_, _35107_);
  and (_35112_, _35111_, _07210_);
  and (_35113_, _35046_, _06541_);
  and (_35115_, _35113_, _35108_);
  or (_35116_, _35115_, _06383_);
  or (_35117_, _35116_, _35112_);
  and (_35118_, _15211_, _07943_);
  or (_35119_, _35032_, _07231_);
  or (_35120_, _35119_, _35118_);
  and (_35121_, _35120_, _07229_);
  and (_35122_, _35121_, _35117_);
  nor (_35123_, _11208_, _13660_);
  or (_35124_, _35123_, _35032_);
  and (_35126_, _35124_, _06528_);
  or (_35127_, _35126_, _06563_);
  or (_35128_, _35127_, _35122_);
  or (_35129_, _35043_, _07241_);
  and (_35130_, _35129_, _06571_);
  and (_35131_, _35130_, _35128_);
  and (_35132_, _35039_, _06199_);
  or (_35133_, _35132_, _06188_);
  or (_35134_, _35133_, _35131_);
  and (_35135_, _15280_, _07943_);
  or (_35137_, _35032_, _06189_);
  or (_35138_, _35137_, _35135_);
  and (_35139_, _35138_, _01452_);
  and (_35140_, _35139_, _35134_);
  or (_35141_, _35140_, _35031_);
  and (_43924_, _35141_, _43223_);
  and (_35142_, _01456_, \oc8051_golden_model_1.SCON [5]);
  and (_35143_, _13660_, \oc8051_golden_model_1.SCON [5]);
  nor (_35144_, _08209_, _13660_);
  or (_35145_, _35144_, _35143_);
  or (_35147_, _35145_, _07142_);
  and (_35148_, _15311_, _07943_);
  or (_35149_, _35148_, _35143_);
  or (_35150_, _35149_, _06252_);
  and (_35151_, _07943_, \oc8051_golden_model_1.ACC [5]);
  or (_35152_, _35151_, _35143_);
  and (_35153_, _35152_, _07123_);
  and (_35154_, _07124_, \oc8051_golden_model_1.SCON [5]);
  or (_35155_, _35154_, _06251_);
  or (_35156_, _35155_, _35153_);
  and (_35158_, _35156_, _06476_);
  and (_35159_, _35158_, _35150_);
  and (_35160_, _13682_, \oc8051_golden_model_1.SCON [5]);
  and (_35161_, _15296_, _08533_);
  or (_35162_, _35161_, _35160_);
  and (_35163_, _35162_, _06475_);
  or (_35164_, _35163_, _06468_);
  or (_35165_, _35164_, _35159_);
  and (_35166_, _35165_, _35147_);
  or (_35167_, _35166_, _06466_);
  or (_35169_, _35152_, _06801_);
  and (_35170_, _35169_, _06484_);
  and (_35171_, _35170_, _35167_);
  and (_35172_, _15294_, _08533_);
  or (_35173_, _35172_, _35160_);
  and (_35174_, _35173_, _06483_);
  or (_35175_, _35174_, _06461_);
  or (_35176_, _35175_, _35171_);
  or (_35177_, _35160_, _15328_);
  and (_35178_, _35177_, _35162_);
  or (_35180_, _35178_, _07164_);
  and (_35181_, _35180_, _06242_);
  and (_35182_, _35181_, _35176_);
  or (_35183_, _35160_, _15344_);
  and (_35184_, _35183_, _06241_);
  and (_35185_, _35184_, _35162_);
  or (_35186_, _35185_, _07187_);
  or (_35187_, _35186_, _35182_);
  or (_35188_, _35145_, _07188_);
  and (_35189_, _35188_, _35187_);
  or (_35191_, _35189_, _07182_);
  and (_35192_, _09113_, _07943_);
  or (_35193_, _35143_, _07183_);
  or (_35194_, _35193_, _35192_);
  and (_35195_, _35194_, _06336_);
  and (_35196_, _35195_, _35191_);
  and (_35197_, _15400_, _07943_);
  or (_35198_, _35197_, _35143_);
  and (_35199_, _35198_, _05968_);
  or (_35200_, _35199_, _06371_);
  or (_35202_, _35200_, _35196_);
  and (_35203_, _08888_, _07943_);
  or (_35204_, _35203_, _35143_);
  or (_35205_, _35204_, _07198_);
  and (_35206_, _35205_, _35202_);
  or (_35207_, _35206_, _06367_);
  and (_35208_, _15416_, _07943_);
  or (_35209_, _35208_, _35143_);
  or (_35210_, _35209_, _07218_);
  and (_35211_, _35210_, _07216_);
  and (_35213_, _35211_, _35207_);
  and (_35214_, _11205_, _07943_);
  or (_35215_, _35214_, _35143_);
  and (_35216_, _35215_, _06533_);
  or (_35217_, _35216_, _35213_);
  and (_35218_, _35217_, _07213_);
  or (_35219_, _35143_, _08212_);
  and (_35220_, _35204_, _06366_);
  and (_35221_, _35220_, _35219_);
  or (_35222_, _35221_, _35218_);
  and (_35224_, _35222_, _07210_);
  and (_35225_, _35152_, _06541_);
  and (_35226_, _35225_, _35219_);
  or (_35227_, _35226_, _06383_);
  or (_35228_, _35227_, _35224_);
  and (_35229_, _15413_, _07943_);
  or (_35230_, _35143_, _07231_);
  or (_35231_, _35230_, _35229_);
  and (_35232_, _35231_, _07229_);
  and (_35233_, _35232_, _35228_);
  nor (_35235_, _11204_, _13660_);
  or (_35236_, _35235_, _35143_);
  and (_35237_, _35236_, _06528_);
  or (_35238_, _35237_, _06563_);
  or (_35239_, _35238_, _35233_);
  or (_35240_, _35149_, _07241_);
  and (_35241_, _35240_, _06571_);
  and (_35242_, _35241_, _35239_);
  and (_35243_, _35173_, _06199_);
  or (_35244_, _35243_, _06188_);
  or (_35246_, _35244_, _35242_);
  and (_35247_, _15477_, _07943_);
  or (_35248_, _35143_, _06189_);
  or (_35249_, _35248_, _35247_);
  and (_35250_, _35249_, _01452_);
  and (_35251_, _35250_, _35246_);
  or (_35252_, _35251_, _35142_);
  and (_43925_, _35252_, _43223_);
  and (_35253_, _01456_, \oc8051_golden_model_1.SCON [6]);
  and (_35254_, _13660_, \oc8051_golden_model_1.SCON [6]);
  nor (_35256_, _08106_, _13660_);
  or (_35257_, _35256_, _35254_);
  or (_35258_, _35257_, _07142_);
  and (_35259_, _15512_, _07943_);
  or (_35260_, _35259_, _35254_);
  or (_35261_, _35260_, _06252_);
  and (_35262_, _07943_, \oc8051_golden_model_1.ACC [6]);
  or (_35263_, _35262_, _35254_);
  and (_35264_, _35263_, _07123_);
  and (_35265_, _07124_, \oc8051_golden_model_1.SCON [6]);
  or (_35267_, _35265_, _06251_);
  or (_35268_, _35267_, _35264_);
  and (_35269_, _35268_, _06476_);
  and (_35270_, _35269_, _35261_);
  and (_35271_, _13682_, \oc8051_golden_model_1.SCON [6]);
  and (_35272_, _15499_, _08533_);
  or (_35273_, _35272_, _35271_);
  and (_35274_, _35273_, _06475_);
  or (_35275_, _35274_, _06468_);
  or (_35276_, _35275_, _35270_);
  and (_35278_, _35276_, _35258_);
  or (_35279_, _35278_, _06466_);
  or (_35280_, _35263_, _06801_);
  and (_35281_, _35280_, _06484_);
  and (_35282_, _35281_, _35279_);
  and (_35283_, _15497_, _08533_);
  or (_35284_, _35283_, _35271_);
  and (_35285_, _35284_, _06483_);
  or (_35286_, _35285_, _06461_);
  or (_35287_, _35286_, _35282_);
  or (_35289_, _35271_, _15529_);
  and (_35290_, _35289_, _35273_);
  or (_35291_, _35290_, _07164_);
  and (_35292_, _35291_, _06242_);
  and (_35293_, _35292_, _35287_);
  or (_35294_, _35271_, _15545_);
  and (_35295_, _35294_, _06241_);
  and (_35296_, _35295_, _35273_);
  or (_35297_, _35296_, _07187_);
  or (_35298_, _35297_, _35293_);
  or (_35300_, _35257_, _07188_);
  and (_35301_, _35300_, _35298_);
  or (_35302_, _35301_, _07182_);
  and (_35303_, _09067_, _07943_);
  or (_35304_, _35254_, _07183_);
  or (_35305_, _35304_, _35303_);
  and (_35306_, _35305_, _06336_);
  and (_35307_, _35306_, _35302_);
  and (_35308_, _15601_, _07943_);
  or (_35309_, _35308_, _35254_);
  and (_35311_, _35309_, _05968_);
  or (_35312_, _35311_, _06371_);
  or (_35313_, _35312_, _35307_);
  and (_35314_, _15608_, _07943_);
  or (_35315_, _35314_, _35254_);
  or (_35316_, _35315_, _07198_);
  and (_35317_, _35316_, _35313_);
  or (_35318_, _35317_, _06367_);
  and (_35319_, _15618_, _07943_);
  or (_35320_, _35319_, _35254_);
  or (_35322_, _35320_, _07218_);
  and (_35323_, _35322_, _07216_);
  and (_35324_, _35323_, _35318_);
  and (_35325_, _11202_, _07943_);
  or (_35326_, _35325_, _35254_);
  and (_35327_, _35326_, _06533_);
  or (_35328_, _35327_, _35324_);
  and (_35329_, _35328_, _07213_);
  or (_35330_, _35254_, _08109_);
  and (_35331_, _35315_, _06366_);
  and (_35333_, _35331_, _35330_);
  or (_35334_, _35333_, _35329_);
  and (_35335_, _35334_, _07210_);
  and (_35336_, _35263_, _06541_);
  and (_35337_, _35336_, _35330_);
  or (_35338_, _35337_, _06383_);
  or (_35339_, _35338_, _35335_);
  and (_35340_, _15615_, _07943_);
  or (_35341_, _35254_, _07231_);
  or (_35342_, _35341_, _35340_);
  and (_35344_, _35342_, _07229_);
  and (_35345_, _35344_, _35339_);
  nor (_35346_, _11201_, _13660_);
  or (_35347_, _35346_, _35254_);
  and (_35348_, _35347_, _06528_);
  or (_35349_, _35348_, _06563_);
  or (_35350_, _35349_, _35345_);
  or (_35351_, _35260_, _07241_);
  and (_35352_, _35351_, _06571_);
  and (_35353_, _35352_, _35350_);
  and (_35355_, _35284_, _06199_);
  or (_35356_, _35355_, _06188_);
  or (_35357_, _35356_, _35353_);
  and (_35358_, _15676_, _07943_);
  or (_35359_, _35254_, _06189_);
  or (_35360_, _35359_, _35358_);
  and (_35361_, _35360_, _01452_);
  and (_35362_, _35361_, _35357_);
  or (_35363_, _35362_, _35253_);
  and (_43926_, _35363_, _43223_);
  nor (_35365_, _01452_, _06235_);
  nor (_35366_, _07928_, _06235_);
  and (_35367_, _07928_, \oc8051_golden_model_1.ACC [0]);
  and (_35368_, _35367_, _08351_);
  or (_35369_, _35368_, _35366_);
  or (_35370_, _35369_, _07210_);
  nor (_35371_, _08351_, _13775_);
  or (_35372_, _35371_, _35366_);
  or (_35373_, _35372_, _06252_);
  or (_35374_, _35367_, _35366_);
  and (_35376_, _35374_, _07123_);
  nor (_35377_, _07123_, _06235_);
  or (_35378_, _35377_, _06251_);
  or (_35379_, _35378_, _35376_);
  and (_35380_, _35379_, _07142_);
  nand (_35381_, _35380_, _35373_);
  nand (_35382_, _35381_, _06838_);
  or (_35383_, _35374_, _06801_);
  and (_35384_, _35383_, _07523_);
  and (_35385_, _35384_, _35382_);
  or (_35387_, _07187_, _07362_);
  or (_35388_, _35387_, _35385_);
  and (_35389_, _08135_, _07325_);
  or (_35390_, _35366_, _07188_);
  or (_35391_, _35390_, _35389_);
  and (_35392_, _35391_, _35388_);
  or (_35393_, _35392_, _07182_);
  or (_35394_, _35366_, _07183_);
  and (_35395_, _09342_, _07928_);
  or (_35396_, _35395_, _35394_);
  and (_35398_, _35396_, _35393_);
  or (_35399_, _35398_, _05968_);
  and (_35400_, _14427_, _08135_);
  or (_35401_, _35366_, _06336_);
  or (_35402_, _35401_, _35400_);
  and (_35403_, _35402_, _07198_);
  and (_35404_, _35403_, _35399_);
  and (_35405_, _07928_, _08908_);
  or (_35406_, _35405_, _35366_);
  and (_35407_, _35406_, _06371_);
  or (_35409_, _35407_, _06367_);
  or (_35410_, _35409_, _35404_);
  and (_35411_, _14442_, _07928_);
  or (_35412_, _35411_, _35366_);
  or (_35413_, _35412_, _07218_);
  and (_35414_, _35413_, _07216_);
  and (_35415_, _35414_, _35410_);
  nor (_35416_, _12526_, _13775_);
  or (_35417_, _35416_, _35366_);
  nor (_35418_, _35368_, _07216_);
  and (_35420_, _35418_, _35417_);
  or (_35421_, _35420_, _35415_);
  and (_35422_, _35421_, _07213_);
  nand (_35423_, _35406_, _06366_);
  nor (_35424_, _35423_, _35371_);
  or (_35425_, _35424_, _06541_);
  or (_35426_, _35425_, _35422_);
  and (_35427_, _35426_, _35370_);
  or (_35428_, _35427_, _06383_);
  and (_35429_, _14325_, _07928_);
  or (_35431_, _35429_, _35366_);
  or (_35432_, _35431_, _07231_);
  and (_35433_, _35432_, _07229_);
  and (_35434_, _35433_, _35428_);
  and (_35435_, _35417_, _06528_);
  or (_35436_, _35435_, _19442_);
  or (_35437_, _35436_, _35434_);
  or (_35438_, _35372_, _06756_);
  and (_35439_, _35438_, _01452_);
  and (_35440_, _35439_, _35437_);
  or (_35442_, _35440_, _35365_);
  and (_43928_, _35442_, _43223_);
  nand (_35443_, _06547_, \oc8051_golden_model_1.SP [1]);
  nand (_35444_, _08135_, _07018_);
  or (_35445_, _35444_, _08302_);
  or (_35446_, _07928_, \oc8051_golden_model_1.SP [1]);
  and (_35447_, _35446_, _06383_);
  and (_35448_, _35447_, _35445_);
  and (_35449_, _11215_, _08135_);
  nor (_35450_, _07928_, _06233_);
  or (_35452_, _35450_, _07210_);
  or (_35453_, _35452_, _35449_);
  and (_35454_, _06237_, _06468_);
  or (_35455_, _35454_, _06466_);
  and (_35456_, _14503_, _08135_);
  not (_35457_, _35456_);
  and (_35458_, _35457_, _35446_);
  or (_35459_, _35458_, _06252_);
  nand (_35460_, _06705_, \oc8051_golden_model_1.SP [1]);
  and (_35461_, _07928_, \oc8051_golden_model_1.ACC [1]);
  or (_35463_, _35461_, _35450_);
  and (_35464_, _35463_, _07123_);
  nor (_35465_, _07123_, _06233_);
  or (_35466_, _35465_, _06705_);
  or (_35467_, _35466_, _35464_);
  and (_35468_, _35467_, _35460_);
  or (_35469_, _35468_, _06251_);
  and (_35470_, _35469_, _12446_);
  and (_35471_, _35470_, _35459_);
  nor (_35472_, _05950_, \oc8051_golden_model_1.SP [1]);
  or (_35474_, _35472_, _35471_);
  or (_35475_, _35474_, _35455_);
  or (_35476_, _35463_, _06801_);
  and (_35477_, _35476_, _07523_);
  and (_35478_, _35477_, _35475_);
  or (_35479_, _07472_, _06249_);
  or (_35480_, _35479_, _35478_);
  nand (_35481_, _07472_, \oc8051_golden_model_1.SP [1]);
  and (_35482_, _35481_, _07188_);
  and (_35483_, _35482_, _35480_);
  nand (_35485_, _08135_, _07120_);
  and (_35486_, _35446_, _07187_);
  and (_35487_, _35486_, _35485_);
  or (_35488_, _35487_, _07182_);
  or (_35489_, _35488_, _35483_);
  or (_35490_, _35450_, _07183_);
  and (_35491_, _09297_, _07928_);
  or (_35492_, _35491_, _35490_);
  and (_35493_, _35492_, _06336_);
  and (_35494_, _35493_, _35489_);
  and (_35496_, _35446_, _05968_);
  or (_35497_, _14609_, _13775_);
  and (_35498_, _35497_, _35496_);
  or (_35499_, _35498_, _35494_);
  and (_35500_, _35499_, _07198_);
  and (_35501_, _35446_, _06371_);
  and (_35502_, _35501_, _35444_);
  or (_35503_, _35502_, _05895_);
  or (_35504_, _35503_, _35500_);
  nand (_35505_, _05895_, \oc8051_golden_model_1.SP [1]);
  and (_35507_, _35505_, _07218_);
  and (_35508_, _35507_, _35504_);
  or (_35509_, _14625_, _13775_);
  and (_35510_, _35446_, _06367_);
  and (_35511_, _35510_, _35509_);
  or (_35512_, _35511_, _06533_);
  or (_35513_, _35512_, _35508_);
  and (_35514_, _11217_, _07928_);
  or (_35515_, _35514_, _35450_);
  or (_35516_, _35515_, _07216_);
  and (_35517_, _35516_, _07213_);
  and (_35518_, _35517_, _35513_);
  or (_35519_, _14623_, _13775_);
  and (_35520_, _35446_, _06366_);
  and (_35521_, _35520_, _35519_);
  or (_35522_, _35521_, _06541_);
  or (_35523_, _35522_, _35518_);
  and (_35524_, _35523_, _35453_);
  or (_35525_, _35524_, _07209_);
  nor (_35526_, _05919_, _06233_);
  nor (_35528_, _35526_, _06383_);
  and (_35529_, _35528_, _35525_);
  or (_35530_, _35529_, _35448_);
  and (_35531_, _35530_, _07229_);
  nor (_35532_, _11216_, _13775_);
  or (_35533_, _35532_, _35450_);
  and (_35534_, _35533_, _06528_);
  or (_35535_, _35534_, _06547_);
  or (_35536_, _35535_, _35531_);
  nand (_35537_, _35536_, _35443_);
  nor (_35539_, _06260_, _07228_);
  nand (_35540_, _35539_, _35537_);
  or (_35541_, _35539_, _06233_);
  and (_35542_, _35541_, _07241_);
  and (_35543_, _35542_, _35540_);
  and (_35544_, _35458_, _06563_);
  or (_35545_, _35544_, _07812_);
  or (_35546_, _35545_, _35543_);
  or (_35547_, _07250_, _06233_);
  and (_35548_, _35547_, _06189_);
  and (_35550_, _35548_, _35546_);
  or (_35551_, _35456_, _35450_);
  and (_35552_, _35551_, _06188_);
  or (_35553_, _35552_, _01456_);
  or (_35554_, _35553_, _35550_);
  or (_35555_, _01452_, \oc8051_golden_model_1.SP [1]);
  and (_35556_, _35555_, _43223_);
  and (_43929_, _35556_, _35554_);
  nor (_35557_, _01452_, _06670_);
  nand (_35558_, _16022_, _05895_);
  nor (_35560_, _13775_, _07578_);
  nor (_35561_, _07928_, _06670_);
  or (_35562_, _35561_, _07188_);
  or (_35563_, _35562_, _35560_);
  and (_35564_, _14712_, _08135_);
  or (_35565_, _35564_, _35561_);
  or (_35566_, _35565_, _06252_);
  and (_35567_, _07928_, \oc8051_golden_model_1.ACC [2]);
  or (_35568_, _35567_, _35561_);
  or (_35569_, _35568_, _07124_);
  or (_35571_, _07123_, \oc8051_golden_model_1.SP [2]);
  and (_35572_, _35571_, _07272_);
  and (_35573_, _35572_, _35569_);
  and (_35574_, _07837_, _06705_);
  or (_35575_, _35574_, _06251_);
  or (_35576_, _35575_, _35573_);
  and (_35577_, _35576_, _05950_);
  and (_35578_, _35577_, _35566_);
  nor (_35579_, _16022_, _05950_);
  or (_35580_, _35579_, _06468_);
  or (_35582_, _35580_, _35578_);
  nand (_35583_, _08614_, _06468_);
  and (_35584_, _35583_, _35582_);
  or (_35585_, _35584_, _06466_);
  or (_35586_, _35568_, _06801_);
  and (_35587_, _35586_, _07523_);
  and (_35588_, _35587_, _35585_);
  or (_35589_, _07522_, _07471_);
  or (_35590_, _35589_, _35588_);
  nor (_35591_, _07837_, _05947_);
  nor (_35593_, _35591_, _05970_);
  and (_35594_, _35593_, _35590_);
  and (_35595_, _07837_, _05970_);
  or (_35596_, _35595_, _07187_);
  or (_35597_, _35596_, _35594_);
  and (_35598_, _35597_, _35563_);
  or (_35599_, _35598_, _07182_);
  or (_35600_, _35561_, _07183_);
  and (_35601_, _09251_, _07928_);
  or (_35602_, _35601_, _35600_);
  and (_35604_, _35602_, _06336_);
  and (_35605_, _35604_, _35599_);
  and (_35606_, _14808_, _07928_);
  or (_35607_, _35606_, _35561_);
  and (_35608_, _35607_, _05968_);
  or (_35609_, _35608_, _06371_);
  or (_35610_, _35609_, _35605_);
  and (_35611_, _07928_, _08945_);
  or (_35612_, _35611_, _35561_);
  or (_35613_, _35612_, _07198_);
  and (_35615_, _35613_, _35610_);
  or (_35616_, _35615_, _05895_);
  and (_35617_, _35616_, _35558_);
  or (_35618_, _35617_, _06367_);
  and (_35619_, _14824_, _07928_);
  or (_35620_, _35619_, _35561_);
  or (_35621_, _35620_, _07218_);
  and (_35622_, _35621_, _07216_);
  and (_35623_, _35622_, _35618_);
  and (_35624_, _11214_, _07928_);
  or (_35626_, _35624_, _35561_);
  and (_35627_, _35626_, _06533_);
  or (_35628_, _35627_, _35623_);
  and (_35629_, _35628_, _07213_);
  or (_35630_, _35561_, _08397_);
  and (_35631_, _35612_, _06366_);
  and (_35632_, _35631_, _35630_);
  or (_35633_, _35632_, _35629_);
  and (_35634_, _35633_, _12719_);
  and (_35635_, _35568_, _06541_);
  and (_35637_, _35635_, _35630_);
  nor (_35638_, _16022_, _05919_);
  or (_35639_, _35638_, _06383_);
  or (_35640_, _35639_, _35637_);
  or (_35641_, _35640_, _35634_);
  and (_35642_, _14821_, _07928_);
  or (_35643_, _35642_, _35561_);
  or (_35644_, _35643_, _07231_);
  and (_35645_, _35644_, _35641_);
  or (_35646_, _35645_, _06528_);
  nor (_35648_, _11213_, _13775_);
  or (_35649_, _35648_, _35561_);
  or (_35650_, _35649_, _07229_);
  and (_35651_, _35650_, _13873_);
  and (_35652_, _35651_, _35646_);
  and (_35653_, _16022_, _06547_);
  or (_35654_, _35653_, _07228_);
  or (_35655_, _35654_, _35652_);
  nor (_35656_, _07837_, _05916_);
  nor (_35657_, _35656_, _06260_);
  and (_35659_, _35657_, _35655_);
  and (_35660_, _16022_, _06260_);
  or (_35661_, _35660_, _06563_);
  or (_35662_, _35661_, _35659_);
  or (_35663_, _35565_, _07241_);
  and (_35664_, _35663_, _07250_);
  and (_35665_, _35664_, _35662_);
  nor (_35666_, _16022_, _07250_);
  or (_35667_, _35666_, _06188_);
  or (_35668_, _35667_, _35665_);
  and (_35670_, _14884_, _08135_);
  or (_35671_, _35561_, _06189_);
  or (_35672_, _35671_, _35670_);
  and (_35673_, _35672_, _01452_);
  and (_35674_, _35673_, _35668_);
  or (_35675_, _35674_, _35557_);
  and (_43930_, _35675_, _43223_);
  nor (_35676_, _01452_, _06559_);
  or (_35677_, _07840_, _07250_);
  or (_35678_, _07840_, _05916_);
  nand (_35680_, _15841_, _05895_);
  nor (_35681_, _13775_, _07713_);
  nor (_35682_, _07928_, _06559_);
  or (_35683_, _35682_, _07182_);
  or (_35684_, _35683_, _35681_);
  and (_35685_, _35684_, _12604_);
  and (_35686_, _14898_, _08135_);
  or (_35687_, _35686_, _35682_);
  or (_35688_, _35687_, _06252_);
  and (_35689_, _07928_, \oc8051_golden_model_1.ACC [3]);
  or (_35691_, _35689_, _35682_);
  and (_35692_, _35691_, _07123_);
  nor (_35693_, _07123_, _06559_);
  or (_35694_, _35693_, _06705_);
  or (_35695_, _35694_, _35692_);
  nand (_35696_, _15841_, _06705_);
  and (_35697_, _35696_, _35695_);
  or (_35698_, _35697_, _06251_);
  and (_35699_, _35698_, _05950_);
  and (_35700_, _35699_, _35688_);
  nor (_35702_, _15841_, _05950_);
  or (_35703_, _35702_, _06468_);
  or (_35704_, _35703_, _35700_);
  nand (_35705_, _08594_, _06468_);
  and (_35706_, _35705_, _35704_);
  or (_35707_, _35706_, _06466_);
  or (_35708_, _35691_, _06801_);
  and (_35709_, _35708_, _07523_);
  and (_35710_, _35709_, _35707_);
  or (_35711_, _07764_, _07472_);
  or (_35713_, _35711_, _35710_);
  nand (_35714_, _15841_, _07472_);
  and (_35715_, _35714_, _07188_);
  and (_35716_, _35715_, _35713_);
  or (_35717_, _35716_, _35685_);
  or (_35718_, _35682_, _07183_);
  and (_35719_, _09205_, _07928_);
  or (_35720_, _35719_, _35718_);
  and (_35721_, _35720_, _06336_);
  and (_35722_, _35721_, _35717_);
  and (_35724_, _15003_, _07928_);
  or (_35725_, _35724_, _35682_);
  and (_35726_, _35725_, _05968_);
  or (_35727_, _35726_, _06371_);
  or (_35728_, _35727_, _35722_);
  and (_35729_, _07928_, _08872_);
  or (_35730_, _35729_, _35682_);
  or (_35731_, _35730_, _07198_);
  and (_35732_, _35731_, _35728_);
  or (_35733_, _35732_, _05895_);
  and (_35735_, _35733_, _35680_);
  or (_35736_, _35735_, _06367_);
  and (_35737_, _15018_, _07928_);
  or (_35738_, _35737_, _35682_);
  or (_35739_, _35738_, _07218_);
  and (_35740_, _35739_, _07216_);
  and (_35741_, _35740_, _35736_);
  and (_35742_, _12523_, _07928_);
  or (_35743_, _35742_, _35682_);
  and (_35744_, _35743_, _06533_);
  or (_35746_, _35744_, _35741_);
  and (_35747_, _35746_, _07213_);
  or (_35748_, _35682_, _08257_);
  and (_35749_, _35730_, _06366_);
  and (_35750_, _35749_, _35748_);
  or (_35751_, _35750_, _35747_);
  and (_35752_, _35751_, _12719_);
  and (_35753_, _35691_, _06541_);
  and (_35754_, _35753_, _35748_);
  nor (_35755_, _15841_, _05919_);
  or (_35757_, _35755_, _06383_);
  or (_35758_, _35757_, _35754_);
  or (_35759_, _35758_, _35752_);
  and (_35760_, _15015_, _08135_);
  or (_35761_, _35682_, _07231_);
  or (_35762_, _35761_, _35760_);
  and (_35763_, _35762_, _35759_);
  or (_35764_, _35763_, _06528_);
  nor (_35765_, _11211_, _13775_);
  or (_35766_, _35765_, _35682_);
  or (_35768_, _35766_, _07229_);
  and (_35769_, _35768_, _13873_);
  and (_35770_, _35769_, _35764_);
  nor (_35771_, _08591_, _06559_);
  or (_35772_, _35771_, _08592_);
  and (_35773_, _35772_, _06547_);
  or (_35774_, _35773_, _07228_);
  or (_35775_, _35774_, _35770_);
  and (_35776_, _35775_, _35678_);
  or (_35777_, _35776_, _06260_);
  or (_35779_, _35772_, _06261_);
  and (_35780_, _35779_, _07241_);
  and (_35781_, _35780_, _35777_);
  and (_35782_, _35687_, _06563_);
  or (_35783_, _35782_, _07812_);
  or (_35784_, _35783_, _35781_);
  and (_35785_, _35784_, _35677_);
  or (_35786_, _35785_, _06188_);
  and (_35787_, _15075_, _08135_);
  or (_35788_, _35682_, _06189_);
  or (_35790_, _35788_, _35787_);
  and (_35791_, _35790_, _01452_);
  and (_35792_, _35791_, _35786_);
  or (_35793_, _35792_, _35676_);
  and (_43932_, _35793_, _43223_);
  nor (_35794_, _01452_, _13805_);
  nor (_35795_, _07719_, \oc8051_golden_model_1.SP [4]);
  nor (_35796_, _35795_, _13789_);
  or (_35797_, _35796_, _07250_);
  or (_35798_, _35796_, _05916_);
  nor (_35800_, _08494_, _13775_);
  nor (_35801_, _07928_, _13805_);
  or (_35802_, _35801_, _07182_);
  or (_35803_, _35802_, _35800_);
  and (_35804_, _35803_, _12604_);
  and (_35805_, _15108_, _08135_);
  or (_35806_, _35805_, _35801_);
  or (_35807_, _35806_, _06252_);
  and (_35808_, _07928_, \oc8051_golden_model_1.ACC [4]);
  or (_35809_, _35808_, _35801_);
  or (_35811_, _35809_, _07124_);
  or (_35812_, _07123_, \oc8051_golden_model_1.SP [4]);
  and (_35813_, _35812_, _07272_);
  and (_35814_, _35813_, _35811_);
  and (_35815_, _35796_, _06705_);
  or (_35816_, _35815_, _06251_);
  or (_35817_, _35816_, _35814_);
  and (_35818_, _35817_, _05950_);
  and (_35819_, _35818_, _35807_);
  and (_35820_, _35796_, _07474_);
  or (_35822_, _35820_, _06468_);
  or (_35823_, _35822_, _35819_);
  and (_35824_, _13806_, _06235_);
  nor (_35825_, _08593_, _13805_);
  nor (_35826_, _35825_, _35824_);
  nand (_35827_, _35826_, _06468_);
  and (_35828_, _35827_, _35823_);
  or (_35829_, _35828_, _06466_);
  or (_35830_, _35809_, _06801_);
  and (_35831_, _35830_, _07523_);
  and (_35833_, _35831_, _35829_);
  and (_35834_, _07720_, \oc8051_golden_model_1.SP [4]);
  nor (_35835_, _07720_, \oc8051_golden_model_1.SP [4]);
  nor (_35836_, _35835_, _35834_);
  and (_35837_, _35836_, _06247_);
  or (_35838_, _35837_, _07472_);
  or (_35839_, _35838_, _35833_);
  or (_35840_, _35796_, _07473_);
  and (_35841_, _35840_, _07188_);
  and (_35842_, _35841_, _35839_);
  or (_35844_, _35842_, _35804_);
  or (_35845_, _35801_, _07183_);
  and (_35846_, _09159_, _07928_);
  or (_35847_, _35846_, _35845_);
  and (_35848_, _35847_, _06336_);
  and (_35849_, _35848_, _35844_);
  and (_35850_, _15198_, _07928_);
  or (_35851_, _35850_, _35801_);
  and (_35852_, _35851_, _05968_);
  or (_35853_, _35852_, _06371_);
  or (_35855_, _35853_, _35849_);
  and (_35856_, _08892_, _07928_);
  or (_35857_, _35856_, _35801_);
  or (_35858_, _35857_, _07198_);
  and (_35859_, _35858_, _35855_);
  or (_35860_, _35859_, _05895_);
  or (_35861_, _35796_, _13846_);
  and (_35862_, _35861_, _35860_);
  or (_35863_, _35862_, _06367_);
  and (_35864_, _15214_, _07928_);
  or (_35866_, _35864_, _35801_);
  or (_35867_, _35866_, _07218_);
  and (_35868_, _35867_, _07216_);
  and (_35869_, _35868_, _35863_);
  and (_35870_, _11209_, _07928_);
  or (_35871_, _35870_, _35801_);
  and (_35872_, _35871_, _06533_);
  or (_35873_, _35872_, _35869_);
  and (_35874_, _35873_, _07213_);
  or (_35875_, _35801_, _08497_);
  and (_35877_, _35857_, _06366_);
  and (_35878_, _35877_, _35875_);
  or (_35879_, _35878_, _35874_);
  and (_35880_, _35879_, _12719_);
  and (_35881_, _35809_, _06541_);
  and (_35882_, _35881_, _35875_);
  and (_35883_, _35796_, _07209_);
  or (_35884_, _35883_, _06383_);
  or (_35885_, _35884_, _35882_);
  or (_35886_, _35885_, _35880_);
  and (_35888_, _15211_, _07928_);
  or (_35889_, _35888_, _35801_);
  or (_35890_, _35889_, _07231_);
  and (_35891_, _35890_, _35886_);
  or (_35892_, _35891_, _06528_);
  nor (_35893_, _11208_, _13775_);
  or (_35894_, _35893_, _35801_);
  or (_35895_, _35894_, _07229_);
  and (_35896_, _35895_, _13873_);
  and (_35897_, _35896_, _35892_);
  nor (_35899_, _08592_, _13805_);
  or (_35900_, _35899_, _13806_);
  and (_35901_, _35900_, _06547_);
  or (_35902_, _35901_, _07228_);
  or (_35903_, _35902_, _35897_);
  and (_35904_, _35903_, _35798_);
  or (_35905_, _35904_, _06260_);
  or (_35906_, _35900_, _06261_);
  and (_35907_, _35906_, _07241_);
  and (_35908_, _35907_, _35905_);
  and (_35910_, _35806_, _06563_);
  or (_35911_, _35910_, _07812_);
  or (_35912_, _35911_, _35908_);
  and (_35913_, _35912_, _35797_);
  or (_35914_, _35913_, _06188_);
  and (_35915_, _15280_, _08135_);
  or (_35916_, _35801_, _06189_);
  or (_35917_, _35916_, _35915_);
  and (_35918_, _35917_, _01452_);
  and (_35919_, _35918_, _35914_);
  or (_35921_, _35919_, _35794_);
  and (_43933_, _35921_, _43223_);
  nor (_35922_, _01452_, _13804_);
  nor (_35923_, _13789_, \oc8051_golden_model_1.SP [5]);
  nor (_35924_, _35923_, _13790_);
  or (_35925_, _35924_, _07250_);
  or (_35926_, _35924_, _05916_);
  nor (_35927_, _08209_, _13775_);
  nor (_35928_, _07928_, _13804_);
  or (_35929_, _35928_, _07182_);
  or (_35931_, _35929_, _35927_);
  and (_35932_, _35931_, _12604_);
  and (_35933_, _15311_, _08135_);
  or (_35934_, _35933_, _35928_);
  or (_35935_, _35934_, _06252_);
  and (_35936_, _07928_, \oc8051_golden_model_1.ACC [5]);
  or (_35937_, _35936_, _35928_);
  or (_35938_, _35937_, _07124_);
  or (_35939_, _07123_, \oc8051_golden_model_1.SP [5]);
  and (_35940_, _35939_, _07272_);
  and (_35942_, _35940_, _35938_);
  and (_35943_, _35924_, _06705_);
  or (_35944_, _35943_, _06251_);
  or (_35945_, _35944_, _35942_);
  and (_35946_, _35945_, _05950_);
  and (_35947_, _35946_, _35935_);
  and (_35948_, _35924_, _07474_);
  or (_35949_, _35948_, _06468_);
  or (_35950_, _35949_, _35947_);
  and (_35951_, _13807_, _06235_);
  nor (_35953_, _35824_, _13804_);
  nor (_35954_, _35953_, _35951_);
  nand (_35955_, _35954_, _06468_);
  and (_35956_, _35955_, _35950_);
  or (_35957_, _35956_, _06466_);
  or (_35958_, _35937_, _06801_);
  and (_35959_, _35958_, _07523_);
  and (_35960_, _35959_, _35957_);
  nor (_35961_, _35834_, \oc8051_golden_model_1.SP [5]);
  nor (_35962_, _35961_, _13819_);
  and (_35964_, _35962_, _06247_);
  or (_35965_, _35964_, _07472_);
  or (_35966_, _35965_, _35960_);
  or (_35967_, _35924_, _07473_);
  and (_35968_, _35967_, _07188_);
  and (_35969_, _35968_, _35966_);
  or (_35970_, _35969_, _35932_);
  or (_35971_, _35928_, _07183_);
  and (_35972_, _09113_, _07928_);
  or (_35973_, _35972_, _35971_);
  and (_35975_, _35973_, _06336_);
  and (_35976_, _35975_, _35970_);
  and (_35977_, _15400_, _07928_);
  or (_35978_, _35977_, _35928_);
  and (_35979_, _35978_, _05968_);
  or (_35980_, _35979_, _06371_);
  or (_35981_, _35980_, _35976_);
  and (_35982_, _08888_, _07928_);
  or (_35983_, _35982_, _35928_);
  or (_35984_, _35983_, _07198_);
  and (_35986_, _35984_, _35981_);
  or (_35987_, _35986_, _05895_);
  or (_35988_, _35924_, _13846_);
  and (_35989_, _35988_, _35987_);
  or (_35990_, _35989_, _06367_);
  and (_35991_, _15416_, _07928_);
  or (_35992_, _35991_, _35928_);
  or (_35993_, _35992_, _07218_);
  and (_35994_, _35993_, _07216_);
  and (_35995_, _35994_, _35990_);
  and (_35997_, _11205_, _07928_);
  or (_35998_, _35997_, _35928_);
  and (_35999_, _35998_, _06533_);
  or (_36000_, _35999_, _35995_);
  and (_36001_, _36000_, _07213_);
  or (_36002_, _35928_, _08212_);
  and (_36003_, _35983_, _06366_);
  and (_36004_, _36003_, _36002_);
  or (_36005_, _36004_, _36001_);
  and (_36006_, _36005_, _12719_);
  and (_36008_, _35937_, _06541_);
  and (_36009_, _36008_, _36002_);
  and (_36010_, _35924_, _07209_);
  or (_36011_, _36010_, _06383_);
  or (_36012_, _36011_, _36009_);
  or (_36013_, _36012_, _36006_);
  and (_36014_, _15413_, _07928_);
  or (_36015_, _36014_, _35928_);
  or (_36016_, _36015_, _07231_);
  and (_36017_, _36016_, _36013_);
  or (_36019_, _36017_, _06528_);
  nor (_36020_, _11204_, _13775_);
  or (_36021_, _36020_, _35928_);
  or (_36022_, _36021_, _07229_);
  and (_36023_, _36022_, _13873_);
  and (_36024_, _36023_, _36019_);
  nor (_36025_, _13806_, _13804_);
  or (_36026_, _36025_, _13807_);
  and (_36027_, _36026_, _06547_);
  or (_36028_, _36027_, _07228_);
  or (_36030_, _36028_, _36024_);
  and (_36031_, _36030_, _35926_);
  or (_36032_, _36031_, _06260_);
  or (_36033_, _36026_, _06261_);
  and (_36034_, _36033_, _07241_);
  and (_36035_, _36034_, _36032_);
  and (_36036_, _35934_, _06563_);
  or (_36037_, _36036_, _07812_);
  or (_36038_, _36037_, _36035_);
  and (_36039_, _36038_, _35925_);
  or (_36041_, _36039_, _06188_);
  and (_36042_, _15477_, _08135_);
  or (_36043_, _35928_, _06189_);
  or (_36044_, _36043_, _36042_);
  and (_36045_, _36044_, _01452_);
  and (_36046_, _36045_, _36041_);
  or (_36047_, _36046_, _35922_);
  and (_43934_, _36047_, _43223_);
  nor (_36048_, _01452_, _13803_);
  nor (_36049_, _07928_, _13803_);
  and (_36051_, _15512_, _08135_);
  or (_36052_, _36051_, _36049_);
  or (_36053_, _36052_, _06252_);
  nor (_36054_, _07123_, _13803_);
  and (_36055_, _07928_, \oc8051_golden_model_1.ACC [6]);
  or (_36056_, _36055_, _36049_);
  and (_36057_, _36056_, _07123_);
  or (_36058_, _36057_, _36054_);
  and (_36059_, _36058_, _07272_);
  nor (_36060_, _13790_, \oc8051_golden_model_1.SP [6]);
  nor (_36062_, _36060_, _13791_);
  and (_36063_, _36062_, _06705_);
  or (_36064_, _36063_, _06251_);
  or (_36065_, _36064_, _36059_);
  and (_36066_, _36065_, _05950_);
  and (_36067_, _36066_, _36053_);
  and (_36068_, _36062_, _07474_);
  or (_36069_, _36068_, _06468_);
  or (_36070_, _36069_, _36067_);
  nor (_36071_, _35951_, _13803_);
  nor (_36073_, _36071_, _13809_);
  nand (_36074_, _36073_, _06468_);
  and (_36075_, _36074_, _36070_);
  or (_36076_, _36075_, _06466_);
  or (_36077_, _36056_, _06801_);
  and (_36078_, _36077_, _07523_);
  and (_36079_, _36078_, _36076_);
  nor (_36080_, _13819_, \oc8051_golden_model_1.SP [6]);
  nor (_36081_, _36080_, _13820_);
  and (_36082_, _36081_, _06247_);
  or (_36084_, _36082_, _36079_);
  and (_36085_, _36084_, _07473_);
  and (_36086_, _36062_, _07472_);
  or (_36087_, _36086_, _07187_);
  or (_36088_, _36087_, _36085_);
  nor (_36089_, _08106_, _13775_);
  or (_36090_, _36049_, _07188_);
  or (_36091_, _36090_, _36089_);
  and (_36092_, _36091_, _36088_);
  or (_36093_, _36092_, _07182_);
  and (_36095_, _09067_, _07928_);
  or (_36096_, _36049_, _07183_);
  or (_36097_, _36096_, _36095_);
  and (_36098_, _36097_, _06336_);
  and (_36099_, _36098_, _36093_);
  and (_36100_, _15601_, _08135_);
  or (_36101_, _36100_, _36049_);
  and (_36102_, _36101_, _05968_);
  or (_36103_, _36102_, _06371_);
  or (_36104_, _36103_, _36099_);
  and (_36106_, _15608_, _07928_);
  or (_36107_, _36106_, _36049_);
  or (_36108_, _36107_, _07198_);
  and (_36109_, _36108_, _36104_);
  or (_36110_, _36109_, _05895_);
  or (_36111_, _36062_, _13846_);
  and (_36112_, _36111_, _36110_);
  or (_36113_, _36112_, _06367_);
  and (_36114_, _15618_, _07928_);
  or (_36115_, _36114_, _36049_);
  or (_36117_, _36115_, _07218_);
  and (_36118_, _36117_, _07216_);
  and (_36119_, _36118_, _36113_);
  and (_36120_, _11202_, _07928_);
  or (_36121_, _36120_, _36049_);
  and (_36122_, _36121_, _06533_);
  or (_36123_, _36122_, _36119_);
  and (_36124_, _36123_, _07213_);
  or (_36125_, _36049_, _08109_);
  and (_36126_, _36107_, _06366_);
  and (_36128_, _36126_, _36125_);
  or (_36129_, _36128_, _36124_);
  and (_36130_, _36129_, _12719_);
  and (_36131_, _36056_, _06541_);
  and (_36132_, _36131_, _36125_);
  and (_36133_, _36062_, _07209_);
  or (_36134_, _36133_, _06383_);
  or (_36135_, _36134_, _36132_);
  or (_36136_, _36135_, _36130_);
  and (_36137_, _15615_, _07928_);
  or (_36139_, _36137_, _36049_);
  or (_36140_, _36139_, _07231_);
  and (_36141_, _36140_, _36136_);
  or (_36142_, _36141_, _06528_);
  nor (_36143_, _11201_, _13775_);
  or (_36144_, _36143_, _36049_);
  or (_36145_, _36144_, _07229_);
  and (_36146_, _36145_, _13873_);
  and (_36147_, _36146_, _36142_);
  nor (_36148_, _13807_, _13803_);
  or (_36150_, _36148_, _13808_);
  and (_36151_, _36150_, _06547_);
  or (_36152_, _36151_, _07228_);
  or (_36153_, _36152_, _36147_);
  nor (_36154_, _36062_, _05916_);
  nor (_36155_, _36154_, _06260_);
  and (_36156_, _36155_, _36153_);
  and (_36157_, _36150_, _06260_);
  or (_36158_, _36157_, _06563_);
  or (_36159_, _36158_, _36156_);
  or (_36161_, _36052_, _07241_);
  and (_36162_, _36161_, _07250_);
  and (_36163_, _36162_, _36159_);
  and (_36164_, _36062_, _07812_);
  or (_36165_, _36164_, _06188_);
  or (_36166_, _36165_, _36163_);
  and (_36167_, _15676_, _08135_);
  or (_36168_, _36049_, _06189_);
  or (_36169_, _36168_, _36167_);
  and (_36170_, _36169_, _01452_);
  and (_36172_, _36170_, _36166_);
  or (_36173_, _36172_, _36048_);
  and (_43935_, _36173_, _43223_);
  not (_36174_, \oc8051_golden_model_1.SBUF [0]);
  nor (_36175_, _01452_, _36174_);
  nand (_36176_, _11218_, _07857_);
  nor (_36177_, _07857_, _36174_);
  nor (_36178_, _36177_, _07210_);
  nand (_36179_, _36178_, _36176_);
  and (_36180_, _07857_, \oc8051_golden_model_1.ACC [0]);
  or (_36182_, _36180_, _36177_);
  and (_36183_, _36182_, _06466_);
  or (_36184_, _36183_, _07187_);
  nor (_36185_, _08351_, _13904_);
  or (_36186_, _36185_, _36177_);
  and (_36187_, _36186_, _06251_);
  nor (_36188_, _07123_, _36174_);
  and (_36189_, _36182_, _07123_);
  or (_36190_, _36189_, _36188_);
  and (_36191_, _36190_, _06252_);
  or (_36193_, _36191_, _06468_);
  or (_36194_, _36193_, _36187_);
  and (_36195_, _36194_, _06801_);
  or (_36196_, _36195_, _36184_);
  and (_36197_, _07857_, _07325_);
  or (_36198_, _36177_, _19463_);
  or (_36199_, _36198_, _36197_);
  and (_36200_, _36199_, _36196_);
  or (_36201_, _36200_, _07182_);
  and (_36202_, _09342_, _07857_);
  or (_36204_, _36177_, _07183_);
  or (_36205_, _36204_, _36202_);
  and (_36206_, _36205_, _36201_);
  or (_36207_, _36206_, _05968_);
  and (_36208_, _14427_, _07857_);
  or (_36209_, _36177_, _06336_);
  or (_36210_, _36209_, _36208_);
  and (_36211_, _36210_, _07198_);
  and (_36212_, _36211_, _36207_);
  and (_36213_, _07857_, _08908_);
  or (_36215_, _36213_, _36177_);
  and (_36216_, _36215_, _06371_);
  or (_36217_, _36216_, _06367_);
  or (_36218_, _36217_, _36212_);
  and (_36219_, _14442_, _07857_);
  or (_36220_, _36219_, _36177_);
  or (_36221_, _36220_, _07218_);
  and (_36222_, _36221_, _07216_);
  and (_36223_, _36222_, _36218_);
  nor (_36224_, _12526_, _13904_);
  or (_36226_, _36224_, _36177_);
  and (_36227_, _36176_, _06533_);
  and (_36228_, _36227_, _36226_);
  or (_36229_, _36228_, _36223_);
  and (_36230_, _36229_, _07213_);
  nand (_36231_, _36215_, _06366_);
  nor (_36232_, _36231_, _36185_);
  or (_36233_, _36232_, _06541_);
  or (_36234_, _36233_, _36230_);
  and (_36235_, _36234_, _36179_);
  or (_36237_, _36235_, _06383_);
  and (_36238_, _14325_, _07857_);
  or (_36239_, _36177_, _07231_);
  or (_36240_, _36239_, _36238_);
  and (_36241_, _36240_, _07229_);
  and (_36242_, _36241_, _36237_);
  and (_36243_, _36226_, _06528_);
  or (_36244_, _36243_, _19442_);
  or (_36245_, _36244_, _36242_);
  or (_36246_, _36186_, _06756_);
  and (_36248_, _36246_, _01452_);
  and (_36249_, _36248_, _36245_);
  or (_36250_, _36249_, _36175_);
  and (_43937_, _36250_, _43223_);
  not (_36251_, \oc8051_golden_model_1.SBUF [1]);
  nor (_36252_, _01452_, _36251_);
  or (_36253_, _07857_, \oc8051_golden_model_1.SBUF [1]);
  and (_36254_, _14503_, _07857_);
  not (_36255_, _36254_);
  and (_36256_, _36255_, _36253_);
  or (_36257_, _36256_, _06252_);
  nor (_36258_, _07857_, _36251_);
  and (_36259_, _07857_, \oc8051_golden_model_1.ACC [1]);
  or (_36260_, _36259_, _36258_);
  and (_36261_, _36260_, _07123_);
  nor (_36262_, _07123_, _36251_);
  or (_36263_, _36262_, _06251_);
  or (_36264_, _36263_, _36261_);
  and (_36265_, _36264_, _07142_);
  and (_36266_, _36265_, _36257_);
  nor (_36268_, _13904_, _07120_);
  or (_36269_, _36268_, _36258_);
  and (_36270_, _36269_, _06468_);
  or (_36271_, _36270_, _36266_);
  and (_36272_, _36271_, _06801_);
  and (_36273_, _36260_, _06466_);
  or (_36274_, _36273_, _07187_);
  or (_36275_, _36274_, _36272_);
  or (_36276_, _36269_, _07188_);
  and (_36277_, _36276_, _07183_);
  and (_36279_, _36277_, _36275_);
  or (_36280_, _09297_, _13904_);
  and (_36281_, _36253_, _07182_);
  and (_36282_, _36281_, _36280_);
  or (_36283_, _36282_, _36279_);
  and (_36284_, _36283_, _06336_);
  or (_36285_, _14609_, _13904_);
  and (_36286_, _36253_, _05968_);
  and (_36287_, _36286_, _36285_);
  or (_36288_, _36287_, _36284_);
  and (_36290_, _36288_, _07198_);
  nand (_36291_, _07857_, _07018_);
  and (_36292_, _36253_, _06371_);
  and (_36293_, _36292_, _36291_);
  or (_36294_, _36293_, _36290_);
  and (_36295_, _36294_, _07218_);
  or (_36296_, _14625_, _13904_);
  and (_36297_, _36253_, _06367_);
  and (_36298_, _36297_, _36296_);
  or (_36299_, _36298_, _06533_);
  or (_36301_, _36299_, _36295_);
  nor (_36302_, _11216_, _13904_);
  or (_36303_, _36302_, _36258_);
  nand (_36304_, _11215_, _07857_);
  and (_36305_, _36304_, _36303_);
  or (_36306_, _36305_, _07216_);
  and (_36307_, _36306_, _07213_);
  and (_36308_, _36307_, _36301_);
  or (_36309_, _14623_, _13904_);
  and (_36310_, _36253_, _06366_);
  and (_36312_, _36310_, _36309_);
  or (_36313_, _36312_, _06541_);
  or (_36314_, _36313_, _36308_);
  nor (_36315_, _36258_, _07210_);
  nand (_36316_, _36315_, _36304_);
  and (_36317_, _36316_, _07231_);
  and (_36318_, _36317_, _36314_);
  or (_36319_, _36291_, _08302_);
  and (_36320_, _36253_, _06383_);
  and (_36321_, _36320_, _36319_);
  or (_36323_, _36321_, _06528_);
  or (_36324_, _36323_, _36318_);
  or (_36325_, _36303_, _07229_);
  and (_36326_, _36325_, _07241_);
  and (_36327_, _36326_, _36324_);
  and (_36328_, _36256_, _06563_);
  or (_36329_, _36328_, _06188_);
  or (_36330_, _36329_, _36327_);
  or (_36331_, _36258_, _06189_);
  or (_36332_, _36331_, _36254_);
  and (_36334_, _36332_, _01452_);
  and (_36335_, _36334_, _36330_);
  or (_36336_, _36335_, _36252_);
  and (_43938_, _36336_, _43223_);
  and (_36337_, _01456_, \oc8051_golden_model_1.SBUF [2]);
  and (_36338_, _13904_, \oc8051_golden_model_1.SBUF [2]);
  and (_36339_, _09251_, _07857_);
  or (_36340_, _36339_, _36338_);
  and (_36341_, _36340_, _07182_);
  and (_36342_, _14712_, _07857_);
  or (_36344_, _36342_, _36338_);
  or (_36345_, _36344_, _06252_);
  and (_36346_, _07857_, \oc8051_golden_model_1.ACC [2]);
  or (_36347_, _36346_, _36338_);
  and (_36348_, _36347_, _07123_);
  and (_36349_, _07124_, \oc8051_golden_model_1.SBUF [2]);
  or (_36350_, _36349_, _06251_);
  or (_36351_, _36350_, _36348_);
  and (_36352_, _36351_, _07142_);
  and (_36353_, _36352_, _36345_);
  nor (_36355_, _13904_, _07578_);
  or (_36356_, _36355_, _36338_);
  and (_36357_, _36356_, _06468_);
  or (_36358_, _36357_, _36353_);
  and (_36359_, _36358_, _06801_);
  and (_36360_, _36347_, _06466_);
  or (_36361_, _36360_, _07187_);
  or (_36362_, _36361_, _36359_);
  or (_36363_, _36356_, _07188_);
  and (_36364_, _36363_, _07183_);
  and (_36366_, _36364_, _36362_);
  or (_36367_, _36366_, _05968_);
  or (_36368_, _36367_, _36341_);
  and (_36369_, _14808_, _07857_);
  or (_36370_, _36338_, _06336_);
  or (_36371_, _36370_, _36369_);
  and (_36372_, _36371_, _07198_);
  and (_36373_, _36372_, _36368_);
  and (_36374_, _07857_, _08945_);
  or (_36375_, _36374_, _36338_);
  and (_36377_, _36375_, _06371_);
  or (_36378_, _36377_, _06367_);
  or (_36379_, _36378_, _36373_);
  and (_36380_, _14824_, _07857_);
  or (_36381_, _36380_, _36338_);
  or (_36382_, _36381_, _07218_);
  and (_36383_, _36382_, _07216_);
  and (_36384_, _36383_, _36379_);
  and (_36385_, _11214_, _07857_);
  or (_36386_, _36385_, _36338_);
  and (_36388_, _36386_, _06533_);
  or (_36389_, _36388_, _36384_);
  and (_36390_, _36389_, _07213_);
  or (_36391_, _36338_, _08397_);
  and (_36392_, _36375_, _06366_);
  and (_36393_, _36392_, _36391_);
  or (_36394_, _36393_, _36390_);
  and (_36395_, _36394_, _07210_);
  and (_36396_, _36347_, _06541_);
  and (_36397_, _36396_, _36391_);
  or (_36399_, _36397_, _06383_);
  or (_36400_, _36399_, _36395_);
  and (_36401_, _14821_, _07857_);
  or (_36402_, _36338_, _07231_);
  or (_36403_, _36402_, _36401_);
  and (_36404_, _36403_, _07229_);
  and (_36405_, _36404_, _36400_);
  nor (_36406_, _11213_, _13904_);
  or (_36407_, _36406_, _36338_);
  and (_36408_, _36407_, _06528_);
  or (_36410_, _36408_, _36405_);
  and (_36411_, _36410_, _07241_);
  and (_36412_, _36344_, _06563_);
  or (_36413_, _36412_, _06188_);
  or (_36414_, _36413_, _36411_);
  and (_36415_, _14884_, _07857_);
  or (_36416_, _36338_, _06189_);
  or (_36417_, _36416_, _36415_);
  and (_36418_, _36417_, _01452_);
  and (_36419_, _36418_, _36414_);
  or (_36421_, _36419_, _36337_);
  and (_43939_, _36421_, _43223_);
  and (_36422_, _13904_, \oc8051_golden_model_1.SBUF [3]);
  and (_36423_, _14898_, _07857_);
  or (_36424_, _36423_, _36422_);
  or (_36425_, _36424_, _06252_);
  and (_36426_, _07857_, \oc8051_golden_model_1.ACC [3]);
  or (_36427_, _36426_, _36422_);
  and (_36428_, _36427_, _07123_);
  and (_36429_, _07124_, \oc8051_golden_model_1.SBUF [3]);
  or (_36431_, _36429_, _06251_);
  or (_36432_, _36431_, _36428_);
  and (_36433_, _36432_, _07142_);
  and (_36434_, _36433_, _36425_);
  nor (_36435_, _13904_, _07713_);
  or (_36436_, _36435_, _36422_);
  and (_36437_, _36436_, _06468_);
  or (_36438_, _36437_, _36434_);
  and (_36439_, _36438_, _06801_);
  and (_36440_, _36427_, _06466_);
  or (_36442_, _36440_, _07187_);
  or (_36443_, _36442_, _36439_);
  or (_36444_, _36436_, _07188_);
  and (_36445_, _36444_, _36443_);
  or (_36446_, _36445_, _07182_);
  and (_36447_, _09205_, _07857_);
  or (_36448_, _36422_, _07183_);
  or (_36449_, _36448_, _36447_);
  and (_36450_, _36449_, _06336_);
  and (_36451_, _36450_, _36446_);
  and (_36453_, _15003_, _07857_);
  or (_36454_, _36453_, _36422_);
  and (_36455_, _36454_, _05968_);
  or (_36456_, _36455_, _06371_);
  or (_36457_, _36456_, _36451_);
  and (_36458_, _07857_, _08872_);
  or (_36459_, _36458_, _36422_);
  or (_36460_, _36459_, _07198_);
  and (_36461_, _36460_, _36457_);
  or (_36462_, _36461_, _06367_);
  and (_36464_, _15018_, _07857_);
  or (_36465_, _36464_, _36422_);
  or (_36466_, _36465_, _07218_);
  and (_36467_, _36466_, _07216_);
  and (_36468_, _36467_, _36462_);
  and (_36469_, _12523_, _07857_);
  or (_36470_, _36469_, _36422_);
  and (_36471_, _36470_, _06533_);
  or (_36472_, _36471_, _36468_);
  and (_36473_, _36472_, _07213_);
  or (_36475_, _36422_, _08257_);
  and (_36476_, _36459_, _06366_);
  and (_36477_, _36476_, _36475_);
  or (_36478_, _36477_, _36473_);
  and (_36479_, _36478_, _07210_);
  and (_36480_, _36427_, _06541_);
  and (_36481_, _36480_, _36475_);
  or (_36482_, _36481_, _06383_);
  or (_36483_, _36482_, _36479_);
  and (_36484_, _15015_, _07857_);
  or (_36486_, _36422_, _07231_);
  or (_36487_, _36486_, _36484_);
  and (_36488_, _36487_, _07229_);
  and (_36489_, _36488_, _36483_);
  nor (_36490_, _11211_, _13904_);
  or (_36491_, _36490_, _36422_);
  and (_36492_, _36491_, _06528_);
  or (_36493_, _36492_, _06563_);
  or (_36494_, _36493_, _36489_);
  or (_36495_, _36424_, _07241_);
  and (_36497_, _36495_, _06189_);
  and (_36498_, _36497_, _36494_);
  and (_36499_, _15075_, _07857_);
  or (_36500_, _36499_, _36422_);
  and (_36501_, _36500_, _06188_);
  or (_36502_, _36501_, _01456_);
  or (_36503_, _36502_, _36498_);
  or (_36504_, _01452_, \oc8051_golden_model_1.SBUF [3]);
  and (_36505_, _36504_, _43223_);
  and (_43940_, _36505_, _36503_);
  and (_36507_, _13904_, \oc8051_golden_model_1.SBUF [4]);
  and (_36508_, _15108_, _07857_);
  or (_36509_, _36508_, _36507_);
  or (_36510_, _36509_, _06252_);
  and (_36511_, _07857_, \oc8051_golden_model_1.ACC [4]);
  or (_36512_, _36511_, _36507_);
  and (_36513_, _36512_, _07123_);
  and (_36514_, _07124_, \oc8051_golden_model_1.SBUF [4]);
  or (_36515_, _36514_, _06251_);
  or (_36516_, _36515_, _36513_);
  and (_36518_, _36516_, _07142_);
  and (_36519_, _36518_, _36510_);
  nor (_36520_, _08494_, _13904_);
  or (_36521_, _36520_, _36507_);
  and (_36522_, _36521_, _06468_);
  or (_36523_, _36522_, _36519_);
  and (_36524_, _36523_, _06801_);
  and (_36525_, _36512_, _06466_);
  or (_36526_, _36525_, _07187_);
  or (_36527_, _36526_, _36524_);
  and (_36529_, _36521_, _07183_);
  or (_36530_, _36529_, _12603_);
  and (_36531_, _36530_, _36527_);
  and (_36532_, _09159_, _07857_);
  or (_36533_, _36532_, _36507_);
  and (_36534_, _36533_, _07182_);
  or (_36535_, _36534_, _05968_);
  or (_36536_, _36535_, _36531_);
  and (_36537_, _15198_, _07857_);
  or (_36538_, _36507_, _06336_);
  or (_36540_, _36538_, _36537_);
  and (_36541_, _36540_, _07198_);
  and (_36542_, _36541_, _36536_);
  and (_36543_, _08892_, _07857_);
  or (_36544_, _36543_, _36507_);
  and (_36545_, _36544_, _06371_);
  or (_36546_, _36545_, _06367_);
  or (_36547_, _36546_, _36542_);
  and (_36548_, _15214_, _07857_);
  or (_36549_, _36548_, _36507_);
  or (_36551_, _36549_, _07218_);
  and (_36552_, _36551_, _07216_);
  and (_36553_, _36552_, _36547_);
  and (_36554_, _11209_, _07857_);
  or (_36555_, _36554_, _36507_);
  and (_36556_, _36555_, _06533_);
  or (_36557_, _36556_, _36553_);
  and (_36558_, _36557_, _07213_);
  or (_36559_, _36507_, _08497_);
  and (_36560_, _36544_, _06366_);
  and (_36562_, _36560_, _36559_);
  or (_36563_, _36562_, _36558_);
  and (_36564_, _36563_, _07210_);
  and (_36565_, _36512_, _06541_);
  and (_36566_, _36565_, _36559_);
  or (_36567_, _36566_, _06383_);
  or (_36568_, _36567_, _36564_);
  and (_36569_, _15211_, _07857_);
  or (_36570_, _36507_, _07231_);
  or (_36571_, _36570_, _36569_);
  and (_36573_, _36571_, _07229_);
  and (_36574_, _36573_, _36568_);
  nor (_36575_, _11208_, _13904_);
  or (_36576_, _36575_, _36507_);
  and (_36577_, _36576_, _06528_);
  or (_36578_, _36577_, _06563_);
  or (_36579_, _36578_, _36574_);
  or (_36580_, _36509_, _07241_);
  and (_36581_, _36580_, _06189_);
  and (_36582_, _36581_, _36579_);
  and (_36584_, _15280_, _07857_);
  or (_36585_, _36584_, _36507_);
  and (_36586_, _36585_, _06188_);
  or (_36587_, _36586_, _01456_);
  or (_36588_, _36587_, _36582_);
  or (_36589_, _01452_, \oc8051_golden_model_1.SBUF [4]);
  and (_36590_, _36589_, _43223_);
  and (_43941_, _36590_, _36588_);
  and (_36591_, _13904_, \oc8051_golden_model_1.SBUF [5]);
  and (_36592_, _15311_, _07857_);
  or (_36594_, _36592_, _36591_);
  or (_36595_, _36594_, _06252_);
  and (_36596_, _07857_, \oc8051_golden_model_1.ACC [5]);
  or (_36597_, _36596_, _36591_);
  and (_36598_, _36597_, _07123_);
  and (_36599_, _07124_, \oc8051_golden_model_1.SBUF [5]);
  or (_36600_, _36599_, _06251_);
  or (_36601_, _36600_, _36598_);
  and (_36602_, _36601_, _07142_);
  and (_36603_, _36602_, _36595_);
  nor (_36605_, _08209_, _13904_);
  or (_36606_, _36605_, _36591_);
  and (_36607_, _36606_, _06468_);
  or (_36608_, _36607_, _36603_);
  and (_36609_, _36608_, _06801_);
  and (_36610_, _36597_, _06466_);
  or (_36611_, _36610_, _07187_);
  or (_36612_, _36611_, _36609_);
  or (_36613_, _36606_, _07188_);
  and (_36614_, _36613_, _36612_);
  or (_36616_, _36614_, _07182_);
  and (_36617_, _09113_, _07857_);
  or (_36618_, _36591_, _07183_);
  or (_36619_, _36618_, _36617_);
  and (_36620_, _36619_, _06336_);
  and (_36621_, _36620_, _36616_);
  and (_36622_, _15400_, _07857_);
  or (_36623_, _36622_, _36591_);
  and (_36624_, _36623_, _05968_);
  or (_36625_, _36624_, _06371_);
  or (_36627_, _36625_, _36621_);
  and (_36628_, _08888_, _07857_);
  or (_36629_, _36628_, _36591_);
  or (_36630_, _36629_, _07198_);
  and (_36631_, _36630_, _36627_);
  or (_36632_, _36631_, _06367_);
  and (_36633_, _15416_, _07857_);
  or (_36634_, _36633_, _36591_);
  or (_36635_, _36634_, _07218_);
  and (_36636_, _36635_, _07216_);
  and (_36638_, _36636_, _36632_);
  and (_36639_, _11205_, _07857_);
  or (_36640_, _36639_, _36591_);
  and (_36641_, _36640_, _06533_);
  or (_36642_, _36641_, _36638_);
  and (_36643_, _36642_, _07213_);
  or (_36644_, _36591_, _08212_);
  and (_36645_, _36629_, _06366_);
  and (_36646_, _36645_, _36644_);
  or (_36647_, _36646_, _36643_);
  and (_36649_, _36647_, _07210_);
  and (_36650_, _36597_, _06541_);
  and (_36651_, _36650_, _36644_);
  or (_36652_, _36651_, _06383_);
  or (_36653_, _36652_, _36649_);
  and (_36654_, _15413_, _07857_);
  or (_36655_, _36591_, _07231_);
  or (_36656_, _36655_, _36654_);
  and (_36657_, _36656_, _07229_);
  and (_36658_, _36657_, _36653_);
  nor (_36660_, _11204_, _13904_);
  or (_36661_, _36660_, _36591_);
  and (_36662_, _36661_, _06528_);
  or (_36663_, _36662_, _06563_);
  or (_36664_, _36663_, _36658_);
  or (_36665_, _36594_, _07241_);
  and (_36666_, _36665_, _06189_);
  and (_36667_, _36666_, _36664_);
  and (_36668_, _15477_, _07857_);
  or (_36669_, _36668_, _36591_);
  and (_36671_, _36669_, _06188_);
  or (_36672_, _36671_, _01456_);
  or (_36673_, _36672_, _36667_);
  or (_36674_, _01452_, \oc8051_golden_model_1.SBUF [5]);
  and (_36675_, _36674_, _43223_);
  and (_43942_, _36675_, _36673_);
  and (_36676_, _13904_, \oc8051_golden_model_1.SBUF [6]);
  nor (_36677_, _08106_, _13904_);
  or (_36678_, _36677_, _36676_);
  or (_36679_, _36678_, _07188_);
  and (_36681_, _15512_, _07857_);
  or (_36682_, _36681_, _36676_);
  or (_36683_, _36682_, _06252_);
  and (_36684_, _07857_, \oc8051_golden_model_1.ACC [6]);
  or (_36685_, _36684_, _36676_);
  and (_36686_, _36685_, _07123_);
  and (_36687_, _07124_, \oc8051_golden_model_1.SBUF [6]);
  or (_36688_, _36687_, _06251_);
  or (_36689_, _36688_, _36686_);
  and (_36690_, _36689_, _07142_);
  and (_36692_, _36690_, _36683_);
  and (_36693_, _36678_, _06468_);
  or (_36694_, _36693_, _36692_);
  and (_36695_, _36694_, _06801_);
  and (_36696_, _36685_, _06466_);
  or (_36697_, _36696_, _07187_);
  or (_36698_, _36697_, _36695_);
  and (_36699_, _36698_, _07183_);
  and (_36700_, _36699_, _36679_);
  and (_36701_, _09067_, _07857_);
  or (_36703_, _36701_, _36676_);
  and (_36704_, _36703_, _07182_);
  or (_36705_, _36704_, _05968_);
  or (_36706_, _36705_, _36700_);
  and (_36707_, _15601_, _07857_);
  or (_36708_, _36676_, _06336_);
  or (_36709_, _36708_, _36707_);
  and (_36710_, _36709_, _07198_);
  and (_36711_, _36710_, _36706_);
  and (_36712_, _15608_, _07857_);
  or (_36714_, _36712_, _36676_);
  and (_36715_, _36714_, _06371_);
  or (_36716_, _36715_, _06367_);
  or (_36717_, _36716_, _36711_);
  and (_36718_, _15618_, _07857_);
  or (_36719_, _36718_, _36676_);
  or (_36720_, _36719_, _07218_);
  and (_36721_, _36720_, _07216_);
  and (_36722_, _36721_, _36717_);
  and (_36723_, _11202_, _07857_);
  or (_36725_, _36723_, _36676_);
  and (_36726_, _36725_, _06533_);
  or (_36727_, _36726_, _36722_);
  and (_36728_, _36727_, _07213_);
  or (_36729_, _36676_, _08109_);
  and (_36730_, _36714_, _06366_);
  and (_36731_, _36730_, _36729_);
  or (_36732_, _36731_, _36728_);
  and (_36733_, _36732_, _07210_);
  and (_36734_, _36685_, _06541_);
  and (_36736_, _36734_, _36729_);
  or (_36737_, _36736_, _06383_);
  or (_36738_, _36737_, _36733_);
  and (_36739_, _15615_, _07857_);
  or (_36740_, _36676_, _07231_);
  or (_36741_, _36740_, _36739_);
  and (_36742_, _36741_, _07229_);
  and (_36743_, _36742_, _36738_);
  nor (_36744_, _11201_, _13904_);
  or (_36745_, _36744_, _36676_);
  and (_36747_, _36745_, _06528_);
  or (_36748_, _36747_, _06563_);
  or (_36749_, _36748_, _36743_);
  or (_36750_, _36682_, _07241_);
  and (_36751_, _36750_, _06189_);
  and (_36752_, _36751_, _36749_);
  and (_36753_, _15676_, _07857_);
  or (_36754_, _36753_, _36676_);
  and (_36755_, _36754_, _06188_);
  or (_36756_, _36755_, _01456_);
  or (_36758_, _36756_, _36752_);
  or (_36759_, _01452_, \oc8051_golden_model_1.SBUF [6]);
  and (_36760_, _36759_, _43223_);
  and (_43943_, _36760_, _36758_);
  not (_36761_, \oc8051_golden_model_1.PSW [0]);
  nor (_36762_, _01452_, _36761_);
  nand (_36763_, _11218_, _07907_);
  nor (_36764_, _07907_, _36761_);
  nor (_36765_, _36764_, _07210_);
  nand (_36766_, _36765_, _36763_);
  and (_36768_, _07907_, _07325_);
  or (_36769_, _36768_, _36764_);
  or (_36770_, _36769_, _07188_);
  nor (_36771_, _08543_, _36761_);
  and (_36772_, _14341_, _08543_);
  or (_36773_, _36772_, _36771_);
  and (_36774_, _36773_, _06475_);
  nor (_36775_, _08351_, _13994_);
  or (_36776_, _36775_, _36764_);
  or (_36777_, _36776_, _06252_);
  and (_36779_, _07907_, \oc8051_golden_model_1.ACC [0]);
  or (_36780_, _36779_, _36764_);
  and (_36781_, _36780_, _07123_);
  nor (_36782_, _07123_, _36761_);
  or (_36783_, _36782_, _06251_);
  or (_36784_, _36783_, _36781_);
  and (_36785_, _36784_, _06476_);
  and (_36786_, _36785_, _36777_);
  or (_36787_, _36786_, _36774_);
  and (_36788_, _36787_, _07142_);
  and (_36790_, _36769_, _06468_);
  or (_36791_, _36790_, _06466_);
  or (_36792_, _36791_, _36788_);
  or (_36793_, _36780_, _06801_);
  and (_36794_, _36793_, _06484_);
  and (_36795_, _36794_, _36792_);
  and (_36796_, _36764_, _06483_);
  or (_36797_, _36796_, _06461_);
  or (_36798_, _36797_, _36795_);
  or (_36799_, _36776_, _07164_);
  and (_36801_, _36799_, _06242_);
  and (_36802_, _36801_, _36798_);
  or (_36803_, _36771_, _14371_);
  and (_36804_, _36803_, _06241_);
  and (_36805_, _36804_, _36773_);
  or (_36806_, _36805_, _07187_);
  or (_36807_, _36806_, _36802_);
  and (_36808_, _36807_, _36770_);
  or (_36809_, _36808_, _07182_);
  and (_36810_, _09342_, _07907_);
  or (_36812_, _36764_, _07183_);
  or (_36813_, _36812_, _36810_);
  and (_36814_, _36813_, _36809_);
  or (_36815_, _36814_, _05968_);
  and (_36816_, _14427_, _07907_);
  or (_36817_, _36764_, _06336_);
  or (_36818_, _36817_, _36816_);
  and (_36819_, _36818_, _07198_);
  and (_36820_, _36819_, _36815_);
  and (_36821_, _07907_, _08908_);
  or (_36823_, _36821_, _36764_);
  and (_36824_, _36823_, _06371_);
  or (_36825_, _36824_, _06367_);
  or (_36826_, _36825_, _36820_);
  and (_36827_, _14442_, _07907_);
  or (_36828_, _36827_, _36764_);
  or (_36829_, _36828_, _07218_);
  and (_36830_, _36829_, _07216_);
  and (_36831_, _36830_, _36826_);
  nor (_36832_, _12526_, _13994_);
  or (_36834_, _36832_, _36764_);
  and (_36835_, _36763_, _06533_);
  and (_36836_, _36835_, _36834_);
  or (_36837_, _36836_, _36831_);
  and (_36838_, _36837_, _07213_);
  nand (_36839_, _36823_, _06366_);
  nor (_36840_, _36839_, _36775_);
  or (_36841_, _36840_, _06541_);
  or (_36842_, _36841_, _36838_);
  and (_36843_, _36842_, _36766_);
  or (_36845_, _36843_, _06383_);
  and (_36846_, _14325_, _07907_);
  or (_36847_, _36764_, _07231_);
  or (_36848_, _36847_, _36846_);
  and (_36849_, _36848_, _07229_);
  and (_36850_, _36849_, _36845_);
  and (_36851_, _36834_, _06528_);
  or (_36852_, _36851_, _06563_);
  or (_36853_, _36852_, _36850_);
  or (_36854_, _36776_, _07241_);
  and (_36856_, _36854_, _36853_);
  or (_36857_, _36856_, _06199_);
  or (_36858_, _36764_, _06571_);
  and (_36859_, _36858_, _36857_);
  or (_36860_, _36859_, _06188_);
  or (_36861_, _36776_, _06189_);
  and (_36862_, _36861_, _01452_);
  and (_36863_, _36862_, _36860_);
  or (_36864_, _36863_, _36762_);
  and (_43945_, _36864_, _43223_);
  not (_36866_, \oc8051_golden_model_1.PSW [1]);
  nor (_36867_, _01452_, _36866_);
  nor (_36868_, _07907_, _36866_);
  nor (_36869_, _11216_, _13994_);
  or (_36870_, _36869_, _36868_);
  or (_36871_, _36870_, _07229_);
  nor (_36872_, _13994_, _07120_);
  or (_36873_, _36872_, _36868_);
  or (_36874_, _36873_, _07142_);
  or (_36875_, _07907_, \oc8051_golden_model_1.PSW [1]);
  and (_36877_, _14503_, _07907_);
  not (_36878_, _36877_);
  and (_36879_, _36878_, _36875_);
  or (_36880_, _36879_, _06252_);
  and (_36881_, _07907_, \oc8051_golden_model_1.ACC [1]);
  or (_36882_, _36881_, _36868_);
  and (_36883_, _36882_, _07123_);
  nor (_36884_, _07123_, _36866_);
  or (_36885_, _36884_, _06251_);
  or (_36886_, _36885_, _36883_);
  and (_36888_, _36886_, _06476_);
  and (_36889_, _36888_, _36880_);
  nor (_36890_, _08543_, _36866_);
  and (_36891_, _14510_, _08543_);
  or (_36892_, _36891_, _36890_);
  and (_36893_, _36892_, _06475_);
  or (_36894_, _36893_, _06468_);
  or (_36895_, _36894_, _36889_);
  and (_36896_, _36895_, _36874_);
  or (_36897_, _36896_, _06466_);
  or (_36899_, _36882_, _06801_);
  and (_36900_, _36899_, _06484_);
  and (_36901_, _36900_, _36897_);
  and (_36902_, _14513_, _08543_);
  or (_36903_, _36902_, _36890_);
  and (_36904_, _36903_, _06483_);
  or (_36905_, _36904_, _06461_);
  or (_36906_, _36905_, _36901_);
  or (_36907_, _36890_, _14509_);
  and (_36908_, _36907_, _36892_);
  or (_36910_, _36908_, _07164_);
  and (_36911_, _36910_, _06242_);
  and (_36912_, _36911_, _36906_);
  or (_36913_, _36890_, _14553_);
  and (_36914_, _36913_, _06241_);
  and (_36915_, _36914_, _36892_);
  or (_36916_, _36915_, _07187_);
  or (_36917_, _36916_, _36912_);
  or (_36918_, _36873_, _07188_);
  and (_36919_, _36918_, _36917_);
  or (_36921_, _36919_, _07182_);
  and (_36922_, _09297_, _07907_);
  or (_36923_, _36922_, _36868_);
  or (_36924_, _36923_, _07183_);
  and (_36925_, _36924_, _06336_);
  and (_36926_, _36925_, _36921_);
  or (_36927_, _14609_, _13994_);
  and (_36928_, _36875_, _05968_);
  and (_36929_, _36928_, _36927_);
  or (_36930_, _36929_, _36926_);
  and (_36932_, _36930_, _07198_);
  nand (_36933_, _07907_, _07018_);
  and (_36934_, _36875_, _06371_);
  and (_36935_, _36934_, _36933_);
  or (_36936_, _36935_, _36932_);
  and (_36937_, _36936_, _07218_);
  or (_36938_, _14625_, _13994_);
  and (_36939_, _36875_, _06367_);
  and (_36940_, _36939_, _36938_);
  or (_36941_, _36940_, _06533_);
  or (_36943_, _36941_, _36937_);
  nand (_36944_, _11215_, _07907_);
  and (_36945_, _36944_, _36870_);
  or (_36946_, _36945_, _07216_);
  and (_36947_, _36946_, _07213_);
  and (_36948_, _36947_, _36943_);
  or (_36949_, _14623_, _13994_);
  and (_36950_, _36875_, _06366_);
  and (_36951_, _36950_, _36949_);
  or (_36952_, _36951_, _06541_);
  or (_36954_, _36952_, _36948_);
  nor (_36955_, _36868_, _07210_);
  nand (_36956_, _36955_, _36944_);
  and (_36957_, _36956_, _07231_);
  and (_36958_, _36957_, _36954_);
  or (_36959_, _36933_, _08302_);
  and (_36960_, _36875_, _06383_);
  and (_36961_, _36960_, _36959_);
  or (_36962_, _36961_, _06528_);
  or (_36963_, _36962_, _36958_);
  and (_36965_, _36963_, _36871_);
  or (_36966_, _36965_, _06563_);
  or (_36967_, _36879_, _07241_);
  and (_36968_, _36967_, _06571_);
  and (_36969_, _36968_, _36966_);
  and (_36970_, _36903_, _06199_);
  or (_36971_, _36970_, _06188_);
  or (_36972_, _36971_, _36969_);
  or (_36973_, _36868_, _06189_);
  or (_36974_, _36973_, _36877_);
  and (_36976_, _36974_, _01452_);
  and (_36977_, _36976_, _36972_);
  or (_36978_, _36977_, _36867_);
  and (_43946_, _36978_, _43223_);
  and (_36979_, _01456_, \oc8051_golden_model_1.PSW [2]);
  and (_36980_, _13994_, \oc8051_golden_model_1.PSW [2]);
  nor (_36981_, _11213_, _13994_);
  or (_36982_, _36981_, _36980_);
  and (_36983_, _36982_, _06528_);
  nor (_36984_, _13994_, _07578_);
  or (_36986_, _36984_, _36980_);
  or (_36987_, _36986_, _07188_);
  nor (_36988_, _10613_, \oc8051_golden_model_1.ACC [7]);
  not (_36989_, _10934_);
  nor (_36990_, _10612_, _36989_);
  nor (_36991_, _36990_, _36988_);
  nor (_36992_, _36991_, _10618_);
  nor (_36993_, _14174_, _10614_);
  nor (_36994_, _36993_, _36992_);
  and (_36995_, _36994_, _10676_);
  nor (_36996_, _36994_, _10676_);
  or (_36997_, _36996_, _36995_);
  and (_36998_, _36997_, _10610_);
  and (_36999_, _14712_, _07907_);
  or (_37000_, _36999_, _36980_);
  or (_37001_, _37000_, _06252_);
  and (_37002_, _07907_, \oc8051_golden_model_1.ACC [2]);
  or (_37003_, _37002_, _36980_);
  and (_37004_, _37003_, _07123_);
  and (_37005_, _07124_, \oc8051_golden_model_1.PSW [2]);
  or (_37007_, _37005_, _06251_);
  or (_37008_, _37007_, _37004_);
  and (_37009_, _37008_, _06476_);
  and (_37010_, _37009_, _37001_);
  not (_37011_, _08543_);
  and (_37012_, _37011_, \oc8051_golden_model_1.PSW [2]);
  and (_37013_, _14702_, _08543_);
  or (_37014_, _37013_, _37012_);
  and (_37015_, _37014_, _06475_);
  or (_37016_, _37015_, _06468_);
  or (_37018_, _37016_, _37010_);
  or (_37019_, _36986_, _07142_);
  and (_37020_, _37019_, _37018_);
  or (_37021_, _37020_, _06466_);
  or (_37022_, _37003_, _06801_);
  and (_37023_, _37022_, _06484_);
  and (_37024_, _37023_, _37021_);
  and (_37025_, _14706_, _08543_);
  or (_37026_, _37025_, _37012_);
  and (_37027_, _37026_, _06483_);
  or (_37029_, _37027_, _06461_);
  or (_37030_, _37029_, _37024_);
  or (_37031_, _37012_, _14739_);
  and (_37032_, _37031_, _37014_);
  or (_37033_, _37032_, _07164_);
  and (_37034_, _37033_, _09494_);
  and (_37035_, _37034_, _37030_);
  or (_37036_, _16520_, _16407_);
  or (_37037_, _37036_, _16632_);
  or (_37038_, _37037_, _16751_);
  or (_37040_, _37038_, _16869_);
  or (_37041_, _37040_, _16986_);
  or (_37042_, _37041_, _10030_);
  or (_37043_, _37042_, _17103_);
  and (_37044_, _37043_, _09487_);
  or (_37045_, _37044_, _12236_);
  or (_37046_, _37045_, _37035_);
  not (_37047_, _10801_);
  nor (_37048_, _10529_, _10459_);
  or (_37049_, _10459_, _08004_);
  and (_37051_, _37049_, _08506_);
  or (_37052_, _37051_, _37048_);
  and (_37053_, _37052_, _14162_);
  nor (_37054_, _37052_, _14162_);
  nor (_37055_, _37054_, _37053_);
  nor (_37056_, _37055_, _37047_);
  and (_37057_, _37055_, _37047_);
  or (_37058_, _37057_, _37056_);
  or (_37059_, _37058_, _10779_);
  and (_37060_, _37059_, _10611_);
  and (_37062_, _37060_, _37046_);
  or (_37063_, _37062_, _36998_);
  and (_37064_, _37063_, _06516_);
  nor (_37065_, _10550_, _14283_);
  nor (_37066_, _10551_, \oc8051_golden_model_1.ACC [7]);
  nor (_37067_, _37066_, _37065_);
  nor (_37068_, _37067_, _10556_);
  nor (_37069_, _14003_, _10552_);
  or (_37070_, _37069_, _37068_);
  nand (_37071_, _37070_, _10605_);
  or (_37073_, _37070_, _10605_);
  and (_37074_, _37073_, _06510_);
  and (_37075_, _37074_, _37071_);
  or (_37076_, _37075_, _10542_);
  or (_37077_, _37076_, _37064_);
  not (_37078_, _10941_);
  nor (_37079_, _10812_, _37078_);
  nor (_37080_, _10813_, \oc8051_golden_model_1.ACC [7]);
  nor (_37081_, _37080_, _37079_);
  not (_37082_, _37081_);
  or (_37084_, _37082_, _14187_);
  nand (_37085_, _37082_, _14187_);
  and (_37086_, _37085_, _37084_);
  and (_37087_, _37086_, _10874_);
  nor (_37088_, _37086_, _10874_);
  or (_37089_, _37088_, _37087_);
  or (_37090_, _37089_, _10543_);
  and (_37091_, _37090_, _06242_);
  and (_37092_, _37091_, _37077_);
  or (_37093_, _37012_, _14703_);
  and (_37095_, _37093_, _06241_);
  and (_37096_, _37095_, _37014_);
  or (_37097_, _37096_, _07187_);
  or (_37098_, _37097_, _37092_);
  and (_37099_, _37098_, _36987_);
  or (_37100_, _37099_, _07182_);
  and (_37101_, _09251_, _07907_);
  or (_37102_, _36980_, _07183_);
  or (_37103_, _37102_, _37101_);
  and (_37104_, _37103_, _06336_);
  and (_37106_, _37104_, _37100_);
  and (_37107_, _14808_, _07907_);
  or (_37108_, _37107_, _36980_);
  and (_37109_, _37108_, _05968_);
  or (_37110_, _37109_, _10046_);
  or (_37111_, _37110_, _37106_);
  nand (_37112_, _10065_, _10058_);
  nand (_37113_, _37112_, _10046_);
  and (_37114_, _37113_, _37111_);
  and (_37115_, _37114_, _07198_);
  and (_37117_, _07907_, _08945_);
  or (_37118_, _37117_, _36980_);
  and (_37119_, _37118_, _06371_);
  or (_37120_, _37119_, _06367_);
  or (_37121_, _37120_, _37115_);
  and (_37122_, _14824_, _07907_);
  or (_37123_, _37122_, _36980_);
  or (_37124_, _37123_, _07218_);
  and (_37125_, _37124_, _07216_);
  and (_37126_, _37125_, _37121_);
  and (_37128_, _11214_, _07907_);
  or (_37129_, _37128_, _36980_);
  and (_37130_, _37129_, _06533_);
  or (_37131_, _37130_, _37126_);
  and (_37132_, _37131_, _07213_);
  or (_37133_, _36980_, _08397_);
  and (_37134_, _37118_, _06366_);
  and (_37135_, _37134_, _37133_);
  or (_37136_, _37135_, _37132_);
  and (_37137_, _37136_, _07210_);
  and (_37139_, _37003_, _06541_);
  and (_37140_, _37139_, _37133_);
  or (_37141_, _37140_, _06383_);
  or (_37142_, _37141_, _37137_);
  and (_37143_, _14821_, _07907_);
  or (_37144_, _37143_, _36980_);
  or (_37145_, _37144_, _07231_);
  and (_37146_, _37145_, _07229_);
  and (_37147_, _37146_, _37142_);
  nor (_37148_, _37147_, _36983_);
  nor (_37150_, _10692_, _05915_);
  and (_37151_, _07492_, _06380_);
  or (_37152_, _37151_, _37150_);
  nor (_37153_, _37152_, _37148_);
  nor (_37154_, _10530_, _05915_);
  nor (_37155_, _37052_, _14242_);
  nor (_37156_, _37155_, _37048_);
  and (_37157_, _37156_, _10521_);
  and (_37158_, _37048_, _10518_);
  or (_37159_, _37158_, _37157_);
  and (_37161_, _37159_, _37152_);
  or (_37162_, _37161_, _37154_);
  or (_37163_, _37162_, _37153_);
  not (_37164_, _37154_);
  or (_37165_, _37159_, _37164_);
  and (_37166_, _37165_, _11022_);
  and (_37167_, _37166_, _37163_);
  not (_37168_, _36991_);
  nor (_37169_, _37168_, _14249_);
  nor (_37170_, _37169_, _36990_);
  and (_37172_, _37170_, _11046_);
  and (_37173_, _36990_, _11043_);
  or (_37174_, _37173_, _37172_);
  and (_37175_, _37174_, _10452_);
  or (_37176_, _37175_, _11052_);
  or (_37177_, _37176_, _37167_);
  nor (_37178_, _37066_, _14254_);
  nor (_37179_, _37178_, _37065_);
  and (_37180_, _37179_, _11076_);
  and (_37181_, _37065_, _11073_);
  or (_37183_, _37181_, _37180_);
  or (_37184_, _37183_, _06538_);
  nor (_37185_, _37082_, _14260_);
  nor (_37186_, _37185_, _37079_);
  and (_37187_, _37186_, _11106_);
  and (_37188_, _37079_, _11103_);
  or (_37189_, _37188_, _37187_);
  or (_37190_, _37189_, _11082_);
  and (_37191_, _37190_, _12103_);
  and (_37192_, _37191_, _37184_);
  and (_37194_, _37192_, _37177_);
  or (_37195_, _11149_, _10915_);
  nand (_37196_, _11149_, _10529_);
  and (_37197_, _37196_, _37195_);
  and (_37198_, _37197_, _12104_);
  or (_37199_, _37198_, _17443_);
  or (_37200_, _37199_, _37194_);
  nand (_37201_, _11192_, _36989_);
  or (_37202_, _11192_, _10933_);
  and (_37203_, _37202_, _37201_);
  or (_37205_, _37203_, _17444_);
  and (_37206_, _37205_, _37200_);
  or (_37207_, _37206_, _17442_);
  or (_37208_, _37203_, _17700_);
  and (_37209_, _37208_, _37207_);
  and (_37210_, _37209_, _12963_);
  or (_37211_, _11232_, _08508_);
  and (_37212_, _37211_, _14285_);
  and (_37213_, _11270_, _37078_);
  or (_37214_, _37213_, _14290_);
  nand (_37216_, _37214_, _07241_);
  or (_37217_, _37216_, _37212_);
  or (_37218_, _37217_, _37210_);
  or (_37219_, _37000_, _07241_);
  and (_37220_, _37219_, _06571_);
  and (_37221_, _37220_, _37218_);
  and (_37222_, _37026_, _06199_);
  or (_37223_, _37222_, _06188_);
  or (_37224_, _37223_, _37221_);
  and (_37225_, _14884_, _07907_);
  or (_37227_, _36980_, _06189_);
  or (_37228_, _37227_, _37225_);
  and (_37229_, _37228_, _01452_);
  and (_37230_, _37229_, _37224_);
  or (_37231_, _37230_, _36979_);
  and (_43947_, _37231_, _43223_);
  nor (_37232_, _01452_, _07728_);
  nor (_37233_, _07907_, _07728_);
  nor (_37234_, _13994_, _07713_);
  or (_37235_, _37234_, _37233_);
  or (_37237_, _37235_, _07188_);
  or (_37238_, _37235_, _07142_);
  and (_37239_, _14898_, _07907_);
  or (_37240_, _37239_, _37233_);
  or (_37241_, _37240_, _06252_);
  and (_37242_, _07907_, \oc8051_golden_model_1.ACC [3]);
  or (_37243_, _37242_, _37233_);
  and (_37244_, _37243_, _07123_);
  nor (_37245_, _07123_, _07728_);
  or (_37246_, _37245_, _06251_);
  or (_37248_, _37246_, _37244_);
  and (_37249_, _37248_, _06476_);
  and (_37250_, _37249_, _37241_);
  nor (_37251_, _08543_, _07728_);
  and (_37252_, _14906_, _08543_);
  or (_37253_, _37252_, _37251_);
  and (_37254_, _37253_, _06475_);
  or (_37255_, _37254_, _06468_);
  or (_37256_, _37255_, _37250_);
  and (_37257_, _37256_, _37238_);
  or (_37259_, _37257_, _06466_);
  or (_37260_, _37243_, _06801_);
  and (_37261_, _37260_, _06484_);
  and (_37262_, _37261_, _37259_);
  and (_37263_, _14904_, _08543_);
  or (_37264_, _37263_, _37251_);
  and (_37265_, _37264_, _06483_);
  or (_37266_, _37265_, _06461_);
  or (_37267_, _37266_, _37262_);
  or (_37268_, _37251_, _14931_);
  and (_37270_, _37268_, _37253_);
  or (_37271_, _37270_, _07164_);
  and (_37272_, _37271_, _06242_);
  and (_37273_, _37272_, _37267_);
  or (_37274_, _37251_, _14947_);
  and (_37275_, _37274_, _06241_);
  and (_37276_, _37275_, _37253_);
  or (_37277_, _37276_, _07187_);
  or (_37278_, _37277_, _37273_);
  and (_37279_, _37278_, _37237_);
  or (_37281_, _37279_, _07182_);
  and (_37282_, _09205_, _07907_);
  or (_37283_, _37282_, _07183_);
  or (_37284_, _37283_, _37233_);
  and (_37285_, _37284_, _06336_);
  and (_37286_, _37285_, _37281_);
  and (_37287_, _15003_, _07907_);
  or (_37288_, _37287_, _37233_);
  and (_37289_, _37288_, _05968_);
  or (_37290_, _37289_, _06371_);
  or (_37292_, _37290_, _37286_);
  and (_37293_, _07907_, _08872_);
  or (_37294_, _37293_, _37233_);
  or (_37295_, _37294_, _07198_);
  and (_37296_, _37295_, _37292_);
  or (_37297_, _37296_, _06367_);
  and (_37298_, _15018_, _07907_);
  or (_37299_, _37298_, _37233_);
  or (_37300_, _37299_, _07218_);
  and (_37301_, _37300_, _07216_);
  and (_37303_, _37301_, _37297_);
  and (_37304_, _12523_, _07907_);
  or (_37305_, _37304_, _37233_);
  and (_37306_, _37305_, _06533_);
  or (_37307_, _37306_, _37303_);
  and (_37308_, _37307_, _07213_);
  or (_37309_, _37233_, _08257_);
  and (_37310_, _37294_, _06366_);
  and (_37311_, _37310_, _37309_);
  or (_37312_, _37311_, _37308_);
  and (_37314_, _37312_, _07210_);
  and (_37315_, _37243_, _06541_);
  and (_37316_, _37315_, _37309_);
  or (_37317_, _37316_, _06383_);
  or (_37318_, _37317_, _37314_);
  and (_37319_, _15015_, _07907_);
  or (_37320_, _37233_, _07231_);
  or (_37321_, _37320_, _37319_);
  and (_37322_, _37321_, _07229_);
  and (_37323_, _37322_, _37318_);
  nor (_37325_, _11211_, _13994_);
  or (_37326_, _37325_, _37233_);
  and (_37327_, _37326_, _06528_);
  or (_37328_, _37327_, _06563_);
  or (_37329_, _37328_, _37323_);
  or (_37330_, _37240_, _07241_);
  and (_37331_, _37330_, _06571_);
  and (_37332_, _37331_, _37329_);
  and (_37333_, _37264_, _06199_);
  or (_37334_, _37333_, _06188_);
  or (_37336_, _37334_, _37332_);
  and (_37337_, _15075_, _07907_);
  or (_37338_, _37233_, _06189_);
  or (_37339_, _37338_, _37337_);
  and (_37340_, _37339_, _01452_);
  and (_37341_, _37340_, _37336_);
  or (_37342_, _37341_, _37232_);
  and (_43948_, _37342_, _43223_);
  and (_37343_, _01456_, \oc8051_golden_model_1.PSW [4]);
  and (_37344_, _13994_, \oc8051_golden_model_1.PSW [4]);
  nor (_37346_, _08494_, _13994_);
  or (_37347_, _37346_, _37344_);
  or (_37348_, _37347_, _07188_);
  and (_37349_, _37011_, \oc8051_golden_model_1.PSW [4]);
  and (_37350_, _15089_, _08543_);
  or (_37351_, _37350_, _37349_);
  and (_37352_, _37351_, _06483_);
  or (_37353_, _37347_, _07142_);
  and (_37354_, _15108_, _07907_);
  or (_37355_, _37354_, _37344_);
  or (_37357_, _37355_, _06252_);
  and (_37358_, _07907_, \oc8051_golden_model_1.ACC [4]);
  or (_37359_, _37358_, _37344_);
  and (_37360_, _37359_, _07123_);
  and (_37361_, _07124_, \oc8051_golden_model_1.PSW [4]);
  or (_37362_, _37361_, _06251_);
  or (_37363_, _37362_, _37360_);
  and (_37364_, _37363_, _06476_);
  and (_37365_, _37364_, _37357_);
  and (_37366_, _15091_, _08543_);
  or (_37368_, _37366_, _37349_);
  and (_37369_, _37368_, _06475_);
  or (_37370_, _37369_, _06468_);
  or (_37371_, _37370_, _37365_);
  and (_37372_, _37371_, _37353_);
  or (_37373_, _37372_, _06466_);
  or (_37374_, _37359_, _06801_);
  and (_37375_, _37374_, _06484_);
  and (_37376_, _37375_, _37373_);
  or (_37377_, _37376_, _37352_);
  and (_37379_, _37377_, _07164_);
  or (_37380_, _37349_, _15125_);
  and (_37381_, _37380_, _06461_);
  and (_37382_, _37381_, _37368_);
  or (_37383_, _37382_, _37379_);
  and (_37384_, _37383_, _06242_);
  or (_37385_, _37349_, _15141_);
  and (_37386_, _37385_, _06241_);
  and (_37387_, _37386_, _37368_);
  or (_37388_, _37387_, _07187_);
  or (_37390_, _37388_, _37384_);
  and (_37391_, _37390_, _37348_);
  or (_37392_, _37391_, _07182_);
  and (_37393_, _09159_, _07907_);
  or (_37394_, _37344_, _07183_);
  or (_37395_, _37394_, _37393_);
  and (_37396_, _37395_, _06336_);
  and (_37397_, _37396_, _37392_);
  and (_37398_, _15198_, _07907_);
  or (_37399_, _37398_, _37344_);
  and (_37401_, _37399_, _05968_);
  or (_37402_, _37401_, _06371_);
  or (_37403_, _37402_, _37397_);
  and (_37404_, _08892_, _07907_);
  or (_37405_, _37404_, _37344_);
  or (_37406_, _37405_, _07198_);
  and (_37407_, _37406_, _37403_);
  or (_37408_, _37407_, _06367_);
  and (_37409_, _15214_, _07907_);
  or (_37410_, _37409_, _37344_);
  or (_37412_, _37410_, _07218_);
  and (_37413_, _37412_, _07216_);
  and (_37414_, _37413_, _37408_);
  and (_37415_, _11209_, _07907_);
  or (_37416_, _37415_, _37344_);
  and (_37417_, _37416_, _06533_);
  or (_37418_, _37417_, _37414_);
  and (_37419_, _37418_, _07213_);
  or (_37420_, _37344_, _08497_);
  and (_37421_, _37405_, _06366_);
  and (_37423_, _37421_, _37420_);
  or (_37424_, _37423_, _37419_);
  and (_37425_, _37424_, _07210_);
  and (_37426_, _37359_, _06541_);
  and (_37427_, _37426_, _37420_);
  or (_37428_, _37427_, _06383_);
  or (_37429_, _37428_, _37425_);
  and (_37430_, _15211_, _07907_);
  or (_37431_, _37344_, _07231_);
  or (_37432_, _37431_, _37430_);
  and (_37434_, _37432_, _07229_);
  and (_37435_, _37434_, _37429_);
  nor (_37436_, _11208_, _13994_);
  or (_37437_, _37436_, _37344_);
  and (_37438_, _37437_, _06528_);
  or (_37439_, _37438_, _06563_);
  or (_37440_, _37439_, _37435_);
  or (_37441_, _37355_, _07241_);
  and (_37442_, _37441_, _06571_);
  and (_37443_, _37442_, _37440_);
  and (_37445_, _37351_, _06199_);
  or (_37446_, _37445_, _06188_);
  or (_37447_, _37446_, _37443_);
  and (_37448_, _15280_, _07907_);
  or (_37449_, _37344_, _06189_);
  or (_37450_, _37449_, _37448_);
  and (_37451_, _37450_, _01452_);
  and (_37452_, _37451_, _37447_);
  or (_37453_, _37452_, _37343_);
  and (_43949_, _37453_, _43223_);
  and (_37455_, _01456_, \oc8051_golden_model_1.PSW [5]);
  and (_37456_, _13994_, \oc8051_golden_model_1.PSW [5]);
  nor (_37457_, _08209_, _13994_);
  or (_37458_, _37457_, _37456_);
  or (_37459_, _37458_, _07188_);
  or (_37460_, _37458_, _07142_);
  and (_37461_, _15311_, _07907_);
  or (_37462_, _37461_, _37456_);
  or (_37463_, _37462_, _06252_);
  and (_37464_, _07907_, \oc8051_golden_model_1.ACC [5]);
  or (_37466_, _37464_, _37456_);
  and (_37467_, _37466_, _07123_);
  and (_37468_, _07124_, \oc8051_golden_model_1.PSW [5]);
  or (_37469_, _37468_, _06251_);
  or (_37470_, _37469_, _37467_);
  and (_37471_, _37470_, _06476_);
  and (_37472_, _37471_, _37463_);
  and (_37473_, _37011_, \oc8051_golden_model_1.PSW [5]);
  and (_37474_, _15296_, _08543_);
  or (_37475_, _37474_, _37473_);
  and (_37477_, _37475_, _06475_);
  or (_37478_, _37477_, _06468_);
  or (_37479_, _37478_, _37472_);
  and (_37480_, _37479_, _37460_);
  or (_37481_, _37480_, _06466_);
  or (_37482_, _37466_, _06801_);
  and (_37483_, _37482_, _06484_);
  and (_37484_, _37483_, _37481_);
  and (_37485_, _15294_, _08543_);
  or (_37486_, _37485_, _37473_);
  and (_37488_, _37486_, _06483_);
  or (_37489_, _37488_, _06461_);
  or (_37490_, _37489_, _37484_);
  or (_37491_, _37473_, _15328_);
  and (_37492_, _37491_, _37475_);
  or (_37493_, _37492_, _07164_);
  and (_37494_, _37493_, _06242_);
  and (_37495_, _37494_, _37490_);
  or (_37496_, _37473_, _15344_);
  and (_37497_, _37496_, _06241_);
  and (_37499_, _37497_, _37475_);
  or (_37500_, _37499_, _07187_);
  or (_37501_, _37500_, _37495_);
  and (_37502_, _37501_, _37459_);
  or (_37503_, _37502_, _07182_);
  and (_37504_, _09113_, _07907_);
  or (_37505_, _37456_, _07183_);
  or (_37506_, _37505_, _37504_);
  and (_37507_, _37506_, _37503_);
  or (_37508_, _37507_, _05968_);
  and (_37510_, _15400_, _07907_);
  or (_37511_, _37456_, _06336_);
  or (_37512_, _37511_, _37510_);
  and (_37513_, _37512_, _07198_);
  and (_37514_, _37513_, _37508_);
  and (_37515_, _08888_, _07907_);
  or (_37516_, _37515_, _37456_);
  and (_37517_, _37516_, _06371_);
  or (_37518_, _37517_, _06367_);
  or (_37519_, _37518_, _37514_);
  and (_37521_, _15416_, _07907_);
  or (_37522_, _37521_, _37456_);
  or (_37523_, _37522_, _07218_);
  and (_37524_, _37523_, _07216_);
  and (_37525_, _37524_, _37519_);
  and (_37526_, _11205_, _07907_);
  or (_37527_, _37526_, _37456_);
  and (_37528_, _37527_, _06533_);
  or (_37529_, _37528_, _37525_);
  and (_37530_, _37529_, _07213_);
  or (_37532_, _37456_, _08212_);
  and (_37533_, _37516_, _06366_);
  and (_37534_, _37533_, _37532_);
  or (_37535_, _37534_, _37530_);
  and (_37536_, _37535_, _07210_);
  and (_37537_, _37466_, _06541_);
  and (_37538_, _37537_, _37532_);
  or (_37539_, _37538_, _06383_);
  or (_37540_, _37539_, _37536_);
  and (_37541_, _15413_, _07907_);
  or (_37543_, _37456_, _07231_);
  or (_37544_, _37543_, _37541_);
  and (_37545_, _37544_, _07229_);
  and (_37546_, _37545_, _37540_);
  nor (_37547_, _11204_, _13994_);
  or (_37548_, _37547_, _37456_);
  and (_37549_, _37548_, _06528_);
  or (_37550_, _37549_, _06563_);
  or (_37551_, _37550_, _37546_);
  or (_37552_, _37462_, _07241_);
  and (_37554_, _37552_, _06571_);
  and (_37555_, _37554_, _37551_);
  and (_37556_, _37486_, _06199_);
  or (_37557_, _37556_, _06188_);
  or (_37558_, _37557_, _37555_);
  and (_37559_, _15477_, _07907_);
  or (_37560_, _37456_, _06189_);
  or (_37561_, _37560_, _37559_);
  and (_37562_, _37561_, _01452_);
  and (_37563_, _37562_, _37558_);
  or (_37565_, _37563_, _37455_);
  and (_43951_, _37565_, _43223_);
  nor (_37566_, _01452_, _18097_);
  or (_37567_, _11097_, _10810_);
  and (_37568_, _37567_, _11050_);
  and (_37569_, _06380_, _06817_);
  not (_37570_, _37150_);
  or (_37571_, _10512_, _10456_);
  or (_37572_, _37571_, _37570_);
  nor (_37573_, _07907_, _18097_);
  nor (_37575_, _08106_, _13994_);
  or (_37576_, _37575_, _37573_);
  or (_37577_, _37576_, _07188_);
  nor (_37578_, _08543_, _18097_);
  and (_37579_, _15499_, _08543_);
  or (_37580_, _37579_, _37578_);
  or (_37581_, _37578_, _15529_);
  and (_37582_, _37581_, _37580_);
  or (_37583_, _37582_, _07164_);
  or (_37584_, _37576_, _07142_);
  and (_37586_, _15512_, _07907_);
  or (_37587_, _37586_, _37573_);
  or (_37588_, _37587_, _06252_);
  and (_37589_, _07907_, \oc8051_golden_model_1.ACC [6]);
  or (_37590_, _37589_, _37573_);
  and (_37591_, _37590_, _07123_);
  nor (_37592_, _07123_, _18097_);
  or (_37593_, _37592_, _06251_);
  or (_37594_, _37593_, _37591_);
  and (_37595_, _37594_, _06476_);
  and (_37597_, _37595_, _37588_);
  and (_37598_, _37580_, _06475_);
  or (_37599_, _37598_, _06468_);
  or (_37600_, _37599_, _37597_);
  and (_37601_, _37600_, _37584_);
  or (_37602_, _37601_, _06466_);
  or (_37603_, _37590_, _06801_);
  and (_37604_, _37603_, _06484_);
  and (_37605_, _37604_, _37602_);
  and (_37606_, _15497_, _08543_);
  or (_37608_, _37606_, _37578_);
  and (_37609_, _37608_, _06483_);
  or (_37610_, _37609_, _06461_);
  or (_37611_, _37610_, _37605_);
  and (_37612_, _37611_, _37583_);
  and (_37613_, _37612_, _10779_);
  or (_37614_, _10456_, _10610_);
  or (_37615_, _37614_, _10794_);
  and (_37616_, _37615_, _12582_);
  or (_37617_, _37616_, _37613_);
  or (_37619_, _10629_, _10611_);
  or (_37620_, _37619_, _10668_);
  and (_37621_, _37620_, _37617_);
  or (_37622_, _37621_, _12589_);
  or (_37623_, _10547_, _06516_);
  or (_37624_, _37623_, _10598_);
  or (_37625_, _10810_, _10543_);
  or (_37626_, _37625_, _10864_);
  and (_37627_, _37626_, _06242_);
  and (_37628_, _37627_, _37624_);
  and (_37630_, _37628_, _37622_);
  or (_37631_, _37578_, _15545_);
  and (_37632_, _37631_, _06241_);
  and (_37633_, _37632_, _37580_);
  or (_37634_, _37633_, _07187_);
  or (_37635_, _37634_, _37630_);
  and (_37636_, _37635_, _37577_);
  or (_37637_, _37636_, _07182_);
  and (_37638_, _09067_, _07907_);
  or (_37639_, _37573_, _07183_);
  or (_37641_, _37639_, _37638_);
  and (_37642_, _37641_, _06336_);
  and (_37643_, _37642_, _37637_);
  and (_37644_, _15601_, _07907_);
  or (_37645_, _37644_, _37573_);
  and (_37646_, _37645_, _05968_);
  or (_37647_, _37646_, _06371_);
  or (_37648_, _37647_, _37643_);
  and (_37649_, _15608_, _07907_);
  or (_37650_, _37649_, _37573_);
  or (_37652_, _37650_, _07198_);
  and (_37653_, _37652_, _37648_);
  or (_37654_, _37653_, _06367_);
  and (_37655_, _15618_, _07907_);
  or (_37656_, _37655_, _37573_);
  or (_37657_, _37656_, _07218_);
  and (_37658_, _37657_, _07216_);
  and (_37659_, _37658_, _37654_);
  and (_37660_, _11202_, _07907_);
  or (_37661_, _37660_, _37573_);
  and (_37663_, _37661_, _06533_);
  or (_37664_, _37663_, _37659_);
  and (_37665_, _37664_, _07213_);
  or (_37666_, _37573_, _08109_);
  and (_37667_, _37650_, _06366_);
  and (_37668_, _37667_, _37666_);
  or (_37669_, _37668_, _37665_);
  and (_37670_, _37669_, _07210_);
  and (_37671_, _37590_, _06541_);
  and (_37672_, _37671_, _37666_);
  or (_37674_, _37672_, _06383_);
  or (_37675_, _37674_, _37670_);
  and (_37676_, _15615_, _07907_);
  or (_37677_, _37676_, _37573_);
  or (_37678_, _37677_, _07231_);
  and (_37679_, _37678_, _37675_);
  or (_37680_, _37679_, _06528_);
  nor (_37681_, _11201_, _13994_);
  or (_37682_, _37681_, _37573_);
  nor (_37683_, _37682_, _07229_);
  nor (_37685_, _37683_, _37151_);
  and (_37686_, _37685_, _37680_);
  and (_37687_, _37571_, _37151_);
  or (_37688_, _37687_, _37150_);
  or (_37689_, _37688_, _37686_);
  and (_37690_, _37689_, _37572_);
  or (_37691_, _37690_, _37569_);
  not (_37692_, _37569_);
  nor (_37693_, _37571_, _37692_);
  nor (_37694_, _37693_, _10522_);
  and (_37696_, _37694_, _37691_);
  and (_37697_, _37571_, _10522_);
  or (_37698_, _37697_, _10452_);
  or (_37699_, _37698_, _37696_);
  or (_37700_, _10629_, _11022_);
  or (_37701_, _37700_, _11037_);
  and (_37702_, _37701_, _37699_);
  or (_37703_, _37702_, _06537_);
  or (_37704_, _10547_, _06538_);
  or (_37705_, _37704_, _11067_);
  and (_37707_, _37705_, _11082_);
  and (_37708_, _37707_, _37703_);
  or (_37709_, _37708_, _37568_);
  and (_37710_, _37709_, _12103_);
  and (_37711_, _12104_, _11142_);
  or (_37712_, _37711_, _11156_);
  or (_37713_, _37712_, _37710_);
  or (_37714_, _11186_, _11160_);
  and (_37715_, _37714_, _06295_);
  and (_37716_, _37715_, _37713_);
  or (_37718_, _11225_, _10450_);
  and (_37719_, _37718_, _12964_);
  or (_37720_, _37719_, _37716_);
  or (_37721_, _11263_, _10451_);
  and (_37722_, _37721_, _07241_);
  and (_37723_, _37722_, _37720_);
  and (_37724_, _37587_, _06563_);
  or (_37725_, _37724_, _37723_);
  and (_37726_, _37725_, _06571_);
  and (_37727_, _37608_, _06199_);
  or (_37729_, _37727_, _06188_);
  or (_37730_, _37729_, _37726_);
  and (_37731_, _15676_, _07907_);
  or (_37732_, _37573_, _06189_);
  or (_37733_, _37732_, _37731_);
  and (_37734_, _37733_, _01452_);
  and (_37735_, _37734_, _37730_);
  or (_37736_, _37735_, _37566_);
  and (_43952_, _37736_, _43223_);
  and (_37737_, _05906_, op0_cnst);
  or (_00001_, _37737_, rst);
  and (_37739_, inst_finished_r, op0_cnst);
  not (_37740_, word_in[3]);
  and (_37741_, _37740_, word_in[2]);
  not (_37742_, _37741_);
  not (_37743_, word_in[1]);
  and (_37744_, _37743_, word_in[0]);
  and (_37745_, _37744_, \oc8051_golden_model_1.IRAM[5] [0]);
  nor (_37746_, _37743_, word_in[0]);
  and (_37747_, _37746_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_37749_, _37747_, _37745_);
  nor (_37750_, word_in[1], word_in[0]);
  and (_37751_, _37750_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_37752_, word_in[1], word_in[0]);
  and (_37753_, _37752_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_37754_, _37753_, _37751_);
  and (_37755_, _37754_, _37749_);
  nor (_37756_, _37755_, _37742_);
  nor (_37757_, _37740_, word_in[2]);
  not (_37758_, _37757_);
  and (_37760_, _37744_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_37761_, _37746_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor (_37762_, _37761_, _37760_);
  and (_37763_, _37750_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_37764_, _37752_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor (_37765_, _37764_, _37763_);
  and (_37766_, _37765_, _37762_);
  nor (_37767_, _37766_, _37758_);
  nor (_37768_, _37767_, _37756_);
  nor (_37769_, word_in[3], word_in[2]);
  not (_37771_, _37769_);
  and (_37772_, _37744_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_37773_, _37746_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_37774_, _37773_, _37772_);
  and (_37775_, _37750_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_37776_, _37752_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor (_37777_, _37776_, _37775_);
  and (_37778_, _37777_, _37774_);
  nor (_37779_, _37778_, _37771_);
  and (_37780_, word_in[3], word_in[2]);
  not (_37782_, _37780_);
  and (_37783_, _37744_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_37784_, _37746_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor (_37785_, _37784_, _37783_);
  and (_37786_, _37750_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_37787_, _37752_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_37788_, _37787_, _37786_);
  and (_37789_, _37788_, _37785_);
  nor (_37790_, _37789_, _37782_);
  nor (_37791_, _37790_, _37779_);
  and (_37793_, _37791_, _37768_);
  and (_37794_, _37746_, _37741_);
  and (_37795_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37796_, _37744_, _37741_);
  and (_37797_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_37798_, _37797_, _37795_);
  and (_37799_, _37757_, _37744_);
  and (_37800_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_37801_, _37769_, _37746_);
  and (_37802_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_37804_, _37802_, _37800_);
  and (_37805_, _37804_, _37798_);
  and (_37806_, _37757_, _37752_);
  and (_37807_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_37808_, _37757_, _37750_);
  and (_37809_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_37810_, _37809_, _37807_);
  and (_37811_, _37780_, _37750_);
  and (_37812_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_37813_, _37769_, _37752_);
  and (_37815_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_37816_, _37815_, _37812_);
  and (_37817_, _37816_, _37810_);
  and (_37818_, _37817_, _37805_);
  and (_37819_, _37780_, _37746_);
  and (_37820_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_37821_, _37780_, _37744_);
  and (_37822_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_37823_, _37822_, _37820_);
  and (_37824_, _37752_, _37741_);
  and (_37826_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37827_, _37750_, _37741_);
  and (_37828_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_37829_, _37828_, _37826_);
  and (_37830_, _37829_, _37823_);
  and (_37831_, _37757_, _37746_);
  and (_37832_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37833_, _37769_, _37744_);
  and (_37834_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37835_, _37834_, _37832_);
  and (_37837_, _37780_, _37752_);
  and (_37838_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_37839_, _37769_, _37750_);
  and (_37840_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_37841_, _37840_, _37838_);
  and (_37842_, _37841_, _37835_);
  and (_37843_, _37842_, _37830_);
  and (_37844_, _37843_, _37818_);
  nand (_37845_, _37844_, _37793_);
  or (_37846_, _37844_, _37793_);
  and (_37848_, _37846_, _37845_);
  and (_37849_, _37744_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_37850_, _37746_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor (_37851_, _37850_, _37849_);
  and (_37852_, _37750_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_37853_, _37752_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor (_37854_, _37853_, _37852_);
  and (_37855_, _37854_, _37851_);
  nor (_37856_, _37855_, _37771_);
  and (_37857_, _37744_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_37859_, _37746_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor (_37860_, _37859_, _37857_);
  and (_37861_, _37750_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_37862_, _37752_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_37863_, _37862_, _37861_);
  and (_37864_, _37863_, _37860_);
  nor (_37865_, _37864_, _37782_);
  nor (_37866_, _37865_, _37856_);
  and (_37867_, _37744_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_37868_, _37746_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_37870_, _37868_, _37867_);
  and (_37871_, _37750_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_37872_, _37752_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_37873_, _37872_, _37871_);
  and (_37874_, _37873_, _37870_);
  nor (_37875_, _37874_, _37742_);
  and (_37876_, _37744_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_37877_, _37746_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor (_37878_, _37877_, _37876_);
  and (_37879_, _37750_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_37881_, _37752_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor (_37882_, _37881_, _37879_);
  and (_37883_, _37882_, _37878_);
  nor (_37884_, _37883_, _37758_);
  nor (_37885_, _37884_, _37875_);
  and (_37886_, _37885_, _37866_);
  not (_37887_, _37886_);
  and (_37888_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_37889_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_37890_, _37889_, _37888_);
  and (_37892_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_37893_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_37894_, _37893_, _37892_);
  and (_37895_, _37894_, _37890_);
  and (_37896_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_37897_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_37898_, _37897_, _37896_);
  and (_37899_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_37900_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_37901_, _37900_, _37899_);
  and (_37903_, _37901_, _37898_);
  and (_37904_, _37903_, _37895_);
  and (_37905_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_37906_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_37907_, _37906_, _37905_);
  and (_37908_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37909_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_37910_, _37909_, _37908_);
  and (_37911_, _37910_, _37907_);
  and (_37912_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_37914_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_37915_, _37914_, _37912_);
  and (_37916_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_37917_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37918_, _37917_, _37916_);
  and (_37919_, _37918_, _37915_);
  and (_37920_, _37919_, _37911_);
  and (_37921_, _37920_, _37904_);
  nor (_37922_, _37921_, _37887_);
  and (_37923_, _37921_, _37887_);
  or (_37925_, _37923_, _37922_);
  or (_37926_, _37925_, _37848_);
  and (_37927_, _37744_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_37928_, _37746_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_37929_, _37928_, _37927_);
  and (_37930_, _37750_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_37931_, _37752_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_37932_, _37931_, _37930_);
  and (_37933_, _37932_, _37929_);
  nor (_37934_, _37933_, _37742_);
  and (_37936_, _37744_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_37937_, _37746_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_37938_, _37937_, _37936_);
  and (_37939_, _37750_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_37940_, _37752_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_37941_, _37940_, _37939_);
  and (_37942_, _37941_, _37938_);
  nor (_37943_, _37942_, _37782_);
  nor (_37944_, _37943_, _37934_);
  and (_37945_, _37744_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_37947_, _37746_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_37948_, _37947_, _37945_);
  and (_37949_, _37750_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_37950_, _37752_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor (_37951_, _37950_, _37949_);
  and (_37952_, _37951_, _37948_);
  nor (_37953_, _37952_, _37771_);
  and (_37954_, _37744_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_37955_, _37746_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor (_37956_, _37955_, _37954_);
  and (_37958_, _37750_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_37959_, _37752_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor (_37960_, _37959_, _37958_);
  and (_37961_, _37960_, _37956_);
  nor (_37962_, _37961_, _37758_);
  nor (_37963_, _37962_, _37953_);
  and (_37964_, _37963_, _37944_);
  and (_37965_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_37966_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_37967_, _37966_, _37965_);
  and (_37969_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_37970_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_37971_, _37970_, _37969_);
  and (_37972_, _37971_, _37967_);
  and (_37973_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_37974_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_37975_, _37974_, _37973_);
  and (_37976_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_37977_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_37978_, _37977_, _37976_);
  and (_37980_, _37978_, _37975_);
  and (_37981_, _37980_, _37972_);
  and (_37982_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_37983_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_37984_, _37983_, _37982_);
  and (_37985_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_37986_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_37987_, _37986_, _37985_);
  and (_37988_, _37987_, _37984_);
  and (_37989_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_37991_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_37992_, _37991_, _37989_);
  and (_37993_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_37994_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_37995_, _37994_, _37993_);
  and (_37996_, _37995_, _37992_);
  and (_37997_, _37996_, _37988_);
  and (_37998_, _37997_, _37981_);
  nand (_37999_, _37998_, _37964_);
  or (_38000_, _37998_, _37964_);
  and (_38002_, _38000_, _37999_);
  and (_38003_, _37744_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_38004_, _37746_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor (_38005_, _38004_, _38003_);
  and (_38006_, _37750_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_38007_, _37752_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor (_38008_, _38007_, _38006_);
  and (_38009_, _38008_, _38005_);
  nor (_38010_, _38009_, _37771_);
  and (_38011_, _37744_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_38013_, _37746_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor (_38014_, _38013_, _38011_);
  and (_38015_, _37750_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_38016_, _37752_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_38017_, _38016_, _38015_);
  and (_38018_, _38017_, _38014_);
  nor (_38019_, _38018_, _37782_);
  nor (_38020_, _38019_, _38010_);
  and (_38021_, _37744_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_38022_, _37746_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_38024_, _38022_, _38021_);
  and (_38025_, _37750_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_38026_, _37752_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_38027_, _38026_, _38025_);
  and (_38028_, _38027_, _38024_);
  nor (_38029_, _38028_, _37742_);
  and (_38030_, _37744_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_38031_, _37746_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor (_38032_, _38031_, _38030_);
  and (_38033_, _37750_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_38035_, _37752_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_38036_, _38035_, _38033_);
  and (_38037_, _38036_, _38032_);
  nor (_38038_, _38037_, _37758_);
  nor (_38039_, _38038_, _38029_);
  and (_38040_, _38039_, _38020_);
  and (_38041_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_38042_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_38043_, _38042_, _38041_);
  and (_38044_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_38046_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_38047_, _38046_, _38044_);
  and (_38048_, _38047_, _38043_);
  and (_38049_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_38050_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_38051_, _38050_, _38049_);
  and (_38052_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_38053_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_38054_, _38053_, _38052_);
  and (_38055_, _38054_, _38051_);
  and (_38057_, _38055_, _38048_);
  and (_38058_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_38059_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_38060_, _38059_, _38058_);
  and (_38061_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_38062_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_38063_, _38062_, _38061_);
  and (_38064_, _38063_, _38060_);
  and (_38065_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_38066_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_38068_, _38066_, _38065_);
  and (_38069_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_38070_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_38071_, _38070_, _38069_);
  and (_38072_, _38071_, _38068_);
  and (_38073_, _38072_, _38064_);
  and (_38074_, _38073_, _38057_);
  nand (_38075_, _38074_, _38040_);
  or (_38076_, _38074_, _38040_);
  and (_38077_, _38076_, _38075_);
  or (_38079_, _38077_, _38002_);
  or (_38080_, _38079_, _37926_);
  and (_38081_, _37744_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_38082_, _37746_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor (_38083_, _38082_, _38081_);
  and (_38084_, _37750_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_38085_, _37752_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor (_38086_, _38085_, _38084_);
  and (_38087_, _38086_, _38083_);
  nor (_38088_, _38087_, _37771_);
  and (_38090_, _37744_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_38091_, _37746_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_38092_, _38091_, _38090_);
  and (_38093_, _37750_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_38094_, _37752_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor (_38095_, _38094_, _38093_);
  and (_38096_, _38095_, _38092_);
  nor (_38097_, _38096_, _37782_);
  nor (_38098_, _38097_, _38088_);
  and (_38099_, _37744_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_38101_, _37746_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor (_38102_, _38101_, _38099_);
  and (_38103_, _37750_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_38104_, _37752_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor (_38105_, _38104_, _38103_);
  and (_38106_, _38105_, _38102_);
  nor (_38107_, _38106_, _37742_);
  and (_38108_, _37744_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_38109_, _37746_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor (_38110_, _38109_, _38108_);
  and (_38112_, _37750_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_38113_, _37752_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_38114_, _38113_, _38112_);
  and (_38115_, _38114_, _38110_);
  nor (_38116_, _38115_, _37758_);
  nor (_38117_, _38116_, _38107_);
  and (_38118_, _38117_, _38098_);
  and (_38119_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_38120_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_38121_, _38120_, _38119_);
  and (_38123_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_38124_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_38125_, _38124_, _38123_);
  and (_38126_, _38125_, _38121_);
  and (_38127_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_38128_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_38129_, _38128_, _38127_);
  and (_38130_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_38131_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_38132_, _38131_, _38130_);
  and (_38134_, _38132_, _38129_);
  and (_38135_, _38134_, _38126_);
  and (_38136_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_38137_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_38138_, _38137_, _38136_);
  and (_38139_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_38140_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_38141_, _38140_, _38139_);
  and (_38142_, _38141_, _38138_);
  and (_38143_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_38145_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_38146_, _38145_, _38143_);
  and (_38147_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_38148_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_38149_, _38148_, _38147_);
  and (_38150_, _38149_, _38146_);
  and (_38151_, _38150_, _38142_);
  and (_38152_, _38151_, _38135_);
  nand (_38153_, _38152_, _38118_);
  or (_38154_, _38152_, _38118_);
  and (_38156_, _38154_, _38153_);
  and (_38157_, _37744_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_38158_, _37746_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor (_38159_, _38158_, _38157_);
  and (_38160_, _37750_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_38161_, _37752_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor (_38162_, _38161_, _38160_);
  and (_38163_, _38162_, _38159_);
  nor (_38164_, _38163_, _37771_);
  and (_38165_, _37744_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_38167_, _37746_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_38168_, _38167_, _38165_);
  and (_38169_, _37750_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_38170_, _37752_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_38171_, _38170_, _38169_);
  and (_38172_, _38171_, _38168_);
  nor (_38173_, _38172_, _37758_);
  nor (_38174_, _38173_, _38164_);
  and (_38175_, _37744_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_38176_, _37746_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor (_38178_, _38176_, _38175_);
  and (_38179_, _37750_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_38180_, _37752_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor (_38181_, _38180_, _38179_);
  and (_38182_, _38181_, _38178_);
  nor (_38183_, _38182_, _37742_);
  and (_38184_, _37744_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_38185_, _37746_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_38186_, _38185_, _38184_);
  and (_38187_, _37750_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_38189_, _37752_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_38190_, _38189_, _38187_);
  and (_38191_, _38190_, _38186_);
  nor (_38192_, _38191_, _37782_);
  nor (_38193_, _38192_, _38183_);
  and (_38194_, _38193_, _38174_);
  not (_38195_, _38194_);
  and (_38196_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_38197_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_38198_, _38197_, _38196_);
  and (_38200_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38201_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_38202_, _38201_, _38200_);
  and (_38203_, _38202_, _38198_);
  and (_38204_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_38205_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_38206_, _38205_, _38204_);
  and (_38207_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_38208_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_38209_, _38208_, _38207_);
  and (_38211_, _38209_, _38206_);
  and (_38212_, _38211_, _38203_);
  and (_38213_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_38214_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_38215_, _38214_, _38213_);
  and (_38216_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_38217_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_38218_, _38217_, _38216_);
  and (_38219_, _38218_, _38215_);
  and (_38220_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_38222_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_38223_, _38222_, _38220_);
  and (_38224_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_38225_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_38226_, _38225_, _38224_);
  and (_38227_, _38226_, _38223_);
  and (_38228_, _38227_, _38219_);
  and (_38229_, _38228_, _38212_);
  nor (_38230_, _38229_, _38195_);
  and (_38231_, _38229_, _38195_);
  or (_38233_, _38231_, _38230_);
  or (_38234_, _38233_, _38156_);
  and (_38235_, _37744_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_38236_, _37746_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor (_38237_, _38236_, _38235_);
  and (_38238_, _37750_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_38239_, _37752_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor (_38240_, _38239_, _38238_);
  and (_38241_, _38240_, _38237_);
  nor (_38242_, _38241_, _37771_);
  and (_38244_, _37744_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_38245_, _37746_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor (_38246_, _38245_, _38244_);
  and (_38247_, _37750_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_38248_, _37752_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor (_38249_, _38248_, _38247_);
  and (_38250_, _38249_, _38246_);
  nor (_38251_, _38250_, _37758_);
  nor (_38252_, _38251_, _38242_);
  and (_38253_, _37744_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_38255_, _37746_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor (_38256_, _38255_, _38253_);
  and (_38257_, _37750_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_38258_, _37752_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor (_38259_, _38258_, _38257_);
  and (_38260_, _38259_, _38256_);
  nor (_38261_, _38260_, _37742_);
  and (_38262_, _37744_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_38263_, _37746_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_38264_, _38263_, _38262_);
  and (_38266_, _37750_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_38267_, _37752_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_38268_, _38267_, _38266_);
  and (_38269_, _38268_, _38264_);
  nor (_38270_, _38269_, _37782_);
  nor (_38271_, _38270_, _38261_);
  and (_38272_, _38271_, _38252_);
  and (_38273_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_38274_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_38275_, _38274_, _38273_);
  and (_38277_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_38278_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_38279_, _38278_, _38277_);
  and (_38280_, _38279_, _38275_);
  and (_38281_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_38282_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_38283_, _38282_, _38281_);
  and (_38284_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_38285_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_38286_, _38285_, _38284_);
  and (_38288_, _38286_, _38283_);
  and (_38289_, _38288_, _38280_);
  and (_38290_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_38291_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_38292_, _38291_, _38290_);
  and (_38293_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_38294_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_38295_, _38294_, _38293_);
  and (_38296_, _38295_, _38292_);
  and (_38297_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_38299_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_38300_, _38299_, _38297_);
  and (_38301_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_38302_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_38303_, _38302_, _38301_);
  and (_38304_, _38303_, _38300_);
  and (_38305_, _38304_, _38296_);
  and (_38306_, _38305_, _38289_);
  nand (_38307_, _38306_, _38272_);
  or (_38308_, _38306_, _38272_);
  and (_38310_, _38308_, _38307_);
  and (_38311_, _37744_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_38312_, _37746_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_38313_, _38312_, _38311_);
  and (_38314_, _37750_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_38315_, _37752_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor (_38316_, _38315_, _38314_);
  and (_38317_, _38316_, _38313_);
  nor (_38318_, _38317_, _37742_);
  and (_38319_, _37744_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_38321_, _37746_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_38322_, _38321_, _38319_);
  and (_38323_, _37750_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_38324_, _37752_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_38325_, _38324_, _38323_);
  and (_38326_, _38325_, _38322_);
  nor (_38327_, _38326_, _37782_);
  nor (_38328_, _38327_, _38318_);
  and (_38329_, _37744_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_38330_, _37746_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor (_38332_, _38330_, _38329_);
  and (_38333_, _37750_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_38334_, _37752_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor (_38335_, _38334_, _38333_);
  and (_38336_, _38335_, _38332_);
  nor (_38337_, _38336_, _37771_);
  and (_38338_, _37744_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_38339_, _37746_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor (_38340_, _38339_, _38338_);
  and (_38341_, _37750_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_38343_, _37752_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor (_38344_, _38343_, _38341_);
  and (_38345_, _38344_, _38340_);
  nor (_38346_, _38345_, _37758_);
  nor (_38347_, _38346_, _38337_);
  and (_38348_, _38347_, _38328_);
  and (_38349_, _37799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_38350_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_38351_, _38350_, _38349_);
  and (_38352_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_38354_, _37796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_38355_, _38354_, _38352_);
  and (_38356_, _38355_, _38351_);
  and (_38357_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_38358_, _37808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_38359_, _38358_, _38357_);
  and (_38360_, _37811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_38361_, _37813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_38362_, _38361_, _38360_);
  and (_38363_, _38362_, _38359_);
  and (_38365_, _38363_, _38356_);
  and (_38366_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_38367_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_38368_, _38367_, _38366_);
  and (_38369_, _37827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_38370_, _37839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_38371_, _38370_, _38369_);
  and (_38372_, _38371_, _38368_);
  and (_38373_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_38374_, _37833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_38376_, _38374_, _38373_);
  and (_38377_, _37837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_38378_, _37821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_38379_, _38378_, _38377_);
  and (_38380_, _38379_, _38376_);
  and (_38381_, _38380_, _38372_);
  and (_38382_, _38381_, _38365_);
  not (_38383_, _38382_);
  nor (_38384_, _38383_, _38348_);
  and (_38385_, _38383_, _38348_);
  or (_38387_, _38385_, _38384_);
  or (_38388_, _38387_, _38310_);
  or (_38389_, _38388_, _38234_);
  or (_38390_, _38389_, _38080_);
  and (property_invalid_iram, _38390_, _37739_);
  nor (_38391_, _10165_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_38392_, _10165_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_38393_, _38392_, _38391_);
  nand (_38394_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38395_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38397_, _38395_, _38394_);
  or (_38398_, _38397_, _38393_);
  and (_38399_, _05937_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38400_, _05937_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38401_, _38400_, _38399_);
  and (_38402_, _05997_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_38403_, \oc8051_golden_model_1.ACC [0], _39465_);
  or (_38404_, _38403_, _38402_);
  or (_38405_, _38404_, _38401_);
  or (_38406_, _38405_, _38398_);
  or (_38408_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38409_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38410_, _38409_, _38408_);
  or (_38411_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38412_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38413_, _38412_, _38411_);
  or (_38414_, _38413_, _38410_);
  nand (_38415_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_38416_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_38417_, _38416_, _38415_);
  and (_38419_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_38420_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38421_, _38420_, _38419_);
  or (_38422_, _38421_, _38417_);
  or (_38423_, _38422_, _38414_);
  or (_38424_, _38423_, _38406_);
  and (property_invalid_acc, _38424_, _37739_);
  and (_38425_, _37737_, _01452_);
  nor (_38426_, _25627_, _01660_);
  and (_38427_, _25627_, _01660_);
  or (_38429_, _38427_, _38426_);
  and (_38430_, _27379_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_38431_, _26002_, _01655_);
  and (_38432_, _26002_, _01655_);
  or (_38433_, _38432_, _38431_);
  nor (_38434_, _27379_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_38435_, _26686_, _01644_);
  and (_38436_, _26686_, _01644_);
  or (_38437_, _38436_, _38435_);
  and (_38438_, _28693_, _38915_);
  nor (_38440_, _28693_, _38915_);
  or (_38441_, _38440_, _38438_);
  nor (_38442_, _29329_, _38921_);
  or (_38443_, _38442_, _38441_);
  nor (_38444_, _27733_, _01620_);
  and (_38445_, _27733_, _01620_);
  or (_38446_, _38445_, _38444_);
  or (_38447_, _38446_, _38443_);
  and (_38448_, _26349_, _01649_);
  nor (_38449_, _26349_, _01649_);
  or (_38451_, _38449_, _38448_);
  and (_38452_, _29329_, _38921_);
  and (_38453_, _29940_, _38892_);
  nor (_38454_, _29940_, _38892_);
  or (_38455_, _38454_, _38453_);
  or (_38456_, _38455_, _38452_);
  nor (_38457_, _27035_, _01635_);
  and (_38458_, _27035_, _01635_);
  or (_38459_, _38458_, _38457_);
  and (_38460_, _28058_, _38904_);
  nor (_38462_, _28058_, _38904_);
  or (_38463_, _38462_, _38460_);
  nor (_38464_, _28385_, _38910_);
  and (_38465_, _28385_, _38910_);
  or (_38466_, _38465_, _38464_);
  nor (_38467_, _13031_, _38888_);
  and (_38468_, _13031_, _38888_);
  and (_38469_, _29636_, _38896_);
  and (_38470_, _29013_, _38900_);
  nor (_38471_, _29013_, _38900_);
  or (_38473_, _38471_, _38470_);
  nor (_38474_, _29636_, _38896_);
  or (_38475_, _25230_, _02059_);
  nand (_38476_, _25230_, _02059_);
  and (_38477_, _38476_, _38475_);
  or (_38478_, _38477_, _38474_);
  or (_38479_, _38478_, _38473_);
  or (_38480_, _38479_, _38469_);
  or (_38481_, _38480_, _38468_);
  or (_38482_, _38481_, _38467_);
  or (_38484_, _38482_, _38466_);
  or (_38485_, _38484_, _38463_);
  or (_38486_, _38485_, _38459_);
  or (_38487_, _38486_, _38456_);
  or (_38488_, _38487_, _38451_);
  or (_38489_, _38488_, _38447_);
  or (_38490_, _38489_, _38437_);
  or (_38491_, _38490_, _38434_);
  or (_38492_, _38491_, _38433_);
  or (_38493_, _38492_, _38430_);
  or (_38495_, _38493_, _38429_);
  and (property_invalid_pc, _38495_, _38425_);
  buf (_00550_, _43226_);
  buf (_05062_, _43223_);
  buf (_05113_, _43223_);
  buf (_05165_, _43223_);
  buf (_05217_, _43223_);
  buf (_05268_, _43223_);
  buf (_05320_, _43223_);
  buf (_05371_, _43223_);
  buf (_05423_, _43223_);
  buf (_05474_, _43223_);
  buf (_05526_, _43223_);
  buf (_05578_, _43223_);
  buf (_05631_, _43223_);
  buf (_05684_, _43223_);
  buf (_05737_, _43223_);
  buf (_05790_, _43223_);
  buf (_05843_, _43223_);
  buf (_39350_, _39249_);
  buf (_39352_, _39251_);
  buf (_39365_, _39249_);
  buf (_39366_, _39251_);
  buf (_39680_, _39269_);
  buf (_39681_, _39270_);
  buf (_39682_, _39272_);
  buf (_39683_, _39273_);
  buf (_39684_, _39274_);
  buf (_39685_, _39275_);
  buf (_39686_, _39276_);
  buf (_39687_, _39278_);
  buf (_39688_, _39279_);
  buf (_39689_, _39280_);
  buf (_39690_, _39281_);
  buf (_39691_, _39282_);
  buf (_39692_, _39284_);
  buf (_39693_, _39285_);
  buf (_39745_, _39269_);
  buf (_39746_, _39270_);
  buf (_39747_, _39272_);
  buf (_39748_, _39273_);
  buf (_39749_, _39274_);
  buf (_39750_, _39275_);
  buf (_39751_, _39276_);
  buf (_39752_, _39278_);
  buf (_39753_, _39279_);
  buf (_39755_, _39280_);
  buf (_39756_, _39281_);
  buf (_39757_, _39282_);
  buf (_39758_, _39284_);
  buf (_39759_, _39285_);
  buf (_40289_, _40063_);
  buf (_40451_, _40063_);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _05066_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _05070_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _05074_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _05077_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _05081_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _05085_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _05089_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _05059_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _05062_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _05117_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _05121_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _05125_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _05129_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _05133_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _05137_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _05141_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _05110_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _05113_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _05582_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _05586_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _05590_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _05594_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _05598_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _05602_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _05606_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _05575_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _05578_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _05635_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _05639_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _05643_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _05647_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _05651_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _05655_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _05659_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _05628_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _05631_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _05688_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _05692_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _05696_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _05700_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _05704_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _05708_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _05712_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _05681_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _05684_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _05741_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _05745_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _05749_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _05753_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _05757_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _05761_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _05765_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _05734_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _05737_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _05794_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _05798_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _05802_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _05806_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _05810_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _05814_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _05818_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _05787_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _05790_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _05847_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _05851_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _05855_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _05859_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _05863_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _05867_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _05871_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _05840_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _05843_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _05169_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _05173_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _05177_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _05181_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _05185_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _05188_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _05192_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _05162_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _05165_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _05220_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _05224_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _05228_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _05232_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _05236_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _05240_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _05244_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _05214_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _05217_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _05272_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _05276_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _05280_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _05284_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _05288_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _05292_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _05295_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _05265_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _05268_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _05324_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _05328_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _05331_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _05335_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _05339_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _05343_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _05347_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _05317_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _05320_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _05375_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _05379_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _05383_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _05387_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _05391_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _05395_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _05399_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _05368_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _05371_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _05427_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _05431_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _05435_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _05439_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _05442_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _05446_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _05450_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _05420_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _05423_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _05478_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _05482_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _05486_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _05490_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _05494_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _05498_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _05502_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _05472_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _05474_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _05530_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _05534_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _05538_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _05542_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _05546_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _05549_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _05553_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _05523_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _05526_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _41399_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _41400_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _41401_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _41403_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _41404_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _41405_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _41406_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _41177_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _41388_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _41389_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _41390_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _41391_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _41392_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _41393_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _41394_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _41395_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _41376_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _41377_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _41378_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _41379_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _41381_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _41382_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _41383_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _41384_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _41364_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _41365_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _41366_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _41367_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _41369_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _41370_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _41371_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _41372_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _41351_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _41353_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _41354_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _41355_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _41356_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _41357_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _41359_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _41360_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _41339_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _41341_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _41342_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _41343_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _41344_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _41345_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _41347_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _41348_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _41327_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _41328_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _41330_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _41331_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _41332_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _41333_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _41334_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _41336_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _41315_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _41316_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _41318_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _41319_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _41320_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _41321_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _41322_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _41324_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _41302_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _41304_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _41305_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _41306_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _41307_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _41308_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _41310_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _41311_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _41289_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _41292_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _41293_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _41294_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _41295_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _41296_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _41298_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _41299_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _41277_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _41278_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _41281_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _41282_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _41283_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _41284_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _41285_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _41287_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _41266_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _41267_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _41269_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _41270_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _41271_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _41272_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _41273_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _41275_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _41255_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _41256_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _41257_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _41258_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _41259_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _41260_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _41262_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _41263_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _41244_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _41245_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _41247_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _41248_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _41249_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _41250_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _41251_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _41253_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _41230_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _41233_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _41234_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _41235_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _41236_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _41237_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _41239_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _41240_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _41219_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _41220_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _41221_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _41222_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _41223_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _41225_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _41226_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _41227_);
  dff (\oc8051_golden_model_1.B [0], _43761_);
  dff (\oc8051_golden_model_1.B [1], _43762_);
  dff (\oc8051_golden_model_1.B [2], _43763_);
  dff (\oc8051_golden_model_1.B [3], _43764_);
  dff (\oc8051_golden_model_1.B [4], _43765_);
  dff (\oc8051_golden_model_1.B [5], _43767_);
  dff (\oc8051_golden_model_1.B [6], _43768_);
  dff (\oc8051_golden_model_1.B [7], _41178_);
  dff (\oc8051_golden_model_1.ACC [0], _43769_);
  dff (\oc8051_golden_model_1.ACC [1], _43771_);
  dff (\oc8051_golden_model_1.ACC [2], _43772_);
  dff (\oc8051_golden_model_1.ACC [3], _43773_);
  dff (\oc8051_golden_model_1.ACC [4], _43774_);
  dff (\oc8051_golden_model_1.ACC [5], _43775_);
  dff (\oc8051_golden_model_1.ACC [6], _43776_);
  dff (\oc8051_golden_model_1.ACC [7], _41179_);
  dff (\oc8051_golden_model_1.PCON [0], _43778_);
  dff (\oc8051_golden_model_1.PCON [1], _43779_);
  dff (\oc8051_golden_model_1.PCON [2], _43780_);
  dff (\oc8051_golden_model_1.PCON [3], _43781_);
  dff (\oc8051_golden_model_1.PCON [4], _43782_);
  dff (\oc8051_golden_model_1.PCON [5], _43783_);
  dff (\oc8051_golden_model_1.PCON [6], _43784_);
  dff (\oc8051_golden_model_1.PCON [7], _41180_);
  dff (\oc8051_golden_model_1.TMOD [0], _43786_);
  dff (\oc8051_golden_model_1.TMOD [1], _43787_);
  dff (\oc8051_golden_model_1.TMOD [2], _43788_);
  dff (\oc8051_golden_model_1.TMOD [3], _43790_);
  dff (\oc8051_golden_model_1.TMOD [4], _43791_);
  dff (\oc8051_golden_model_1.TMOD [5], _43792_);
  dff (\oc8051_golden_model_1.TMOD [6], _43793_);
  dff (\oc8051_golden_model_1.TMOD [7], _41181_);
  dff (\oc8051_golden_model_1.DPL [0], _43795_);
  dff (\oc8051_golden_model_1.DPL [1], _43796_);
  dff (\oc8051_golden_model_1.DPL [2], _43797_);
  dff (\oc8051_golden_model_1.DPL [3], _43798_);
  dff (\oc8051_golden_model_1.DPL [4], _43799_);
  dff (\oc8051_golden_model_1.DPL [5], _43800_);
  dff (\oc8051_golden_model_1.DPL [6], _43801_);
  dff (\oc8051_golden_model_1.DPL [7], _41182_);
  dff (\oc8051_golden_model_1.DPH [0], _43803_);
  dff (\oc8051_golden_model_1.DPH [1], _43804_);
  dff (\oc8051_golden_model_1.DPH [2], _43805_);
  dff (\oc8051_golden_model_1.DPH [3], _43806_);
  dff (\oc8051_golden_model_1.DPH [4], _43807_);
  dff (\oc8051_golden_model_1.DPH [5], _43809_);
  dff (\oc8051_golden_model_1.DPH [6], _43810_);
  dff (\oc8051_golden_model_1.DPH [7], _41185_);
  dff (\oc8051_golden_model_1.TL1 [0], _43811_);
  dff (\oc8051_golden_model_1.TL1 [1], _43813_);
  dff (\oc8051_golden_model_1.TL1 [2], _43814_);
  dff (\oc8051_golden_model_1.TL1 [3], _43815_);
  dff (\oc8051_golden_model_1.TL1 [4], _43816_);
  dff (\oc8051_golden_model_1.TL1 [5], _43817_);
  dff (\oc8051_golden_model_1.TL1 [6], _43818_);
  dff (\oc8051_golden_model_1.TL1 [7], _41186_);
  dff (\oc8051_golden_model_1.TL0 [0], _43820_);
  dff (\oc8051_golden_model_1.TL0 [1], _43821_);
  dff (\oc8051_golden_model_1.TL0 [2], _43822_);
  dff (\oc8051_golden_model_1.TL0 [3], _43823_);
  dff (\oc8051_golden_model_1.TL0 [4], _43824_);
  dff (\oc8051_golden_model_1.TL0 [5], _43825_);
  dff (\oc8051_golden_model_1.TL0 [6], _43826_);
  dff (\oc8051_golden_model_1.TL0 [7], _41187_);
  dff (\oc8051_golden_model_1.TCON [0], _43828_);
  dff (\oc8051_golden_model_1.TCON [1], _43829_);
  dff (\oc8051_golden_model_1.TCON [2], _43830_);
  dff (\oc8051_golden_model_1.TCON [3], _43832_);
  dff (\oc8051_golden_model_1.TCON [4], _43833_);
  dff (\oc8051_golden_model_1.TCON [5], _43834_);
  dff (\oc8051_golden_model_1.TCON [6], _43835_);
  dff (\oc8051_golden_model_1.TCON [7], _41188_);
  dff (\oc8051_golden_model_1.TH1 [0], _43837_);
  dff (\oc8051_golden_model_1.TH1 [1], _43838_);
  dff (\oc8051_golden_model_1.TH1 [2], _43839_);
  dff (\oc8051_golden_model_1.TH1 [3], _43840_);
  dff (\oc8051_golden_model_1.TH1 [4], _43841_);
  dff (\oc8051_golden_model_1.TH1 [5], _43842_);
  dff (\oc8051_golden_model_1.TH1 [6], _43843_);
  dff (\oc8051_golden_model_1.TH1 [7], _41189_);
  dff (\oc8051_golden_model_1.TH0 [0], _43845_);
  dff (\oc8051_golden_model_1.TH0 [1], _43846_);
  dff (\oc8051_golden_model_1.TH0 [2], _43847_);
  dff (\oc8051_golden_model_1.TH0 [3], _43848_);
  dff (\oc8051_golden_model_1.TH0 [4], _43849_);
  dff (\oc8051_golden_model_1.TH0 [5], _43851_);
  dff (\oc8051_golden_model_1.TH0 [6], _43852_);
  dff (\oc8051_golden_model_1.TH0 [7], _41191_);
  dff (\oc8051_golden_model_1.PC [0], _43854_);
  dff (\oc8051_golden_model_1.PC [1], _43855_);
  dff (\oc8051_golden_model_1.PC [2], _43856_);
  dff (\oc8051_golden_model_1.PC [3], _43858_);
  dff (\oc8051_golden_model_1.PC [4], _43859_);
  dff (\oc8051_golden_model_1.PC [5], _43860_);
  dff (\oc8051_golden_model_1.PC [6], _43861_);
  dff (\oc8051_golden_model_1.PC [7], _43862_);
  dff (\oc8051_golden_model_1.PC [8], _43863_);
  dff (\oc8051_golden_model_1.PC [9], _43864_);
  dff (\oc8051_golden_model_1.PC [10], _43865_);
  dff (\oc8051_golden_model_1.PC [11], _43866_);
  dff (\oc8051_golden_model_1.PC [12], _43867_);
  dff (\oc8051_golden_model_1.PC [13], _43869_);
  dff (\oc8051_golden_model_1.PC [14], _43870_);
  dff (\oc8051_golden_model_1.PC [15], _41192_);
  dff (\oc8051_golden_model_1.P2 [0], _43871_);
  dff (\oc8051_golden_model_1.P2 [1], _43873_);
  dff (\oc8051_golden_model_1.P2 [2], _43874_);
  dff (\oc8051_golden_model_1.P2 [3], _43875_);
  dff (\oc8051_golden_model_1.P2 [4], _43876_);
  dff (\oc8051_golden_model_1.P2 [5], _43877_);
  dff (\oc8051_golden_model_1.P2 [6], _43878_);
  dff (\oc8051_golden_model_1.P2 [7], _41193_);
  dff (\oc8051_golden_model_1.P3 [0], _43880_);
  dff (\oc8051_golden_model_1.P3 [1], _43881_);
  dff (\oc8051_golden_model_1.P3 [2], _43882_);
  dff (\oc8051_golden_model_1.P3 [3], _43883_);
  dff (\oc8051_golden_model_1.P3 [4], _43884_);
  dff (\oc8051_golden_model_1.P3 [5], _43885_);
  dff (\oc8051_golden_model_1.P3 [6], _43886_);
  dff (\oc8051_golden_model_1.P3 [7], _41194_);
  dff (\oc8051_golden_model_1.P0 [0], _43888_);
  dff (\oc8051_golden_model_1.P0 [1], _43889_);
  dff (\oc8051_golden_model_1.P0 [2], _43890_);
  dff (\oc8051_golden_model_1.P0 [3], _43892_);
  dff (\oc8051_golden_model_1.P0 [4], _43893_);
  dff (\oc8051_golden_model_1.P0 [5], _43894_);
  dff (\oc8051_golden_model_1.P0 [6], _43895_);
  dff (\oc8051_golden_model_1.P0 [7], _41195_);
  dff (\oc8051_golden_model_1.P1 [0], _43897_);
  dff (\oc8051_golden_model_1.P1 [1], _43898_);
  dff (\oc8051_golden_model_1.P1 [2], _43899_);
  dff (\oc8051_golden_model_1.P1 [3], _43900_);
  dff (\oc8051_golden_model_1.P1 [4], _43901_);
  dff (\oc8051_golden_model_1.P1 [5], _43902_);
  dff (\oc8051_golden_model_1.P1 [6], _43903_);
  dff (\oc8051_golden_model_1.P1 [7], _41197_);
  dff (\oc8051_golden_model_1.IP [0], _43904_);
  dff (\oc8051_golden_model_1.IP [1], _43905_);
  dff (\oc8051_golden_model_1.IP [2], _43906_);
  dff (\oc8051_golden_model_1.IP [3], _43907_);
  dff (\oc8051_golden_model_1.IP [4], _43908_);
  dff (\oc8051_golden_model_1.IP [5], _43910_);
  dff (\oc8051_golden_model_1.IP [6], _43911_);
  dff (\oc8051_golden_model_1.IP [7], _41198_);
  dff (\oc8051_golden_model_1.IE [0], _43912_);
  dff (\oc8051_golden_model_1.IE [1], _43913_);
  dff (\oc8051_golden_model_1.IE [2], _43914_);
  dff (\oc8051_golden_model_1.IE [3], _43915_);
  dff (\oc8051_golden_model_1.IE [4], _43916_);
  dff (\oc8051_golden_model_1.IE [5], _43917_);
  dff (\oc8051_golden_model_1.IE [6], _43918_);
  dff (\oc8051_golden_model_1.IE [7], _41199_);
  dff (\oc8051_golden_model_1.SCON [0], _43920_);
  dff (\oc8051_golden_model_1.SCON [1], _43921_);
  dff (\oc8051_golden_model_1.SCON [2], _43922_);
  dff (\oc8051_golden_model_1.SCON [3], _43923_);
  dff (\oc8051_golden_model_1.SCON [4], _43924_);
  dff (\oc8051_golden_model_1.SCON [5], _43925_);
  dff (\oc8051_golden_model_1.SCON [6], _43926_);
  dff (\oc8051_golden_model_1.SCON [7], _41200_);
  dff (\oc8051_golden_model_1.SP [0], _43928_);
  dff (\oc8051_golden_model_1.SP [1], _43929_);
  dff (\oc8051_golden_model_1.SP [2], _43930_);
  dff (\oc8051_golden_model_1.SP [3], _43932_);
  dff (\oc8051_golden_model_1.SP [4], _43933_);
  dff (\oc8051_golden_model_1.SP [5], _43934_);
  dff (\oc8051_golden_model_1.SP [6], _43935_);
  dff (\oc8051_golden_model_1.SP [7], _41201_);
  dff (\oc8051_golden_model_1.SBUF [0], _43937_);
  dff (\oc8051_golden_model_1.SBUF [1], _43938_);
  dff (\oc8051_golden_model_1.SBUF [2], _43939_);
  dff (\oc8051_golden_model_1.SBUF [3], _43940_);
  dff (\oc8051_golden_model_1.SBUF [4], _43941_);
  dff (\oc8051_golden_model_1.SBUF [5], _43942_);
  dff (\oc8051_golden_model_1.SBUF [6], _43943_);
  dff (\oc8051_golden_model_1.SBUF [7], _41202_);
  dff (\oc8051_golden_model_1.PSW [0], _43945_);
  dff (\oc8051_golden_model_1.PSW [1], _43946_);
  dff (\oc8051_golden_model_1.PSW [2], _43947_);
  dff (\oc8051_golden_model_1.PSW [3], _43948_);
  dff (\oc8051_golden_model_1.PSW [4], _43949_);
  dff (\oc8051_golden_model_1.PSW [5], _43951_);
  dff (\oc8051_golden_model_1.PSW [6], _43952_);
  dff (\oc8051_golden_model_1.PSW [7], _41203_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02843_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02854_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02876_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02902_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02927_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00953_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02938_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00924_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02951_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02963_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02975_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02988_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03000_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03011_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03024_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00973_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02346_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22107_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02538_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02716_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02889_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03129_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03335_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03513_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03714_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03913_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04014_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04110_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04209_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04309_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04408_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04502_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04600_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24267_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _39261_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _39263_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _39264_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _39265_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _39266_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _39267_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _39268_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _39248_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _39269_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _39270_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _39272_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _39273_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _39274_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _39275_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _39276_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _39249_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _39278_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _39279_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _39280_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _39281_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _39282_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _39284_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _39285_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _39251_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34167_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34170_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09667_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34172_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34174_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09670_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34176_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09673_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34178_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34180_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34182_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09676_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34184_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09679_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _09682_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09741_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09743_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09646_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09746_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09749_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09649_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _09752_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _09652_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _09755_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _09758_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09761_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09764_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09767_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09770_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09773_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _09655_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09658_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34165_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09664_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09776_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09661_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _40063_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _40162_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _40163_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _40164_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _40165_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _40166_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _40167_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _40168_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _40064_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _40169_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _40170_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _40171_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _40173_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _40174_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _40175_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _40176_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _40065_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _40177_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _40178_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _40179_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _40180_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _40181_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _40182_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _40184_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _40066_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _40185_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _40186_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _40187_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _40188_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _40189_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _40190_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _40191_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _40068_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _40192_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _40193_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _40195_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _40196_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _40197_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _40198_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _40199_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _40069_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _40200_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _40201_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _40202_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _40203_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _40204_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _40206_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _40207_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _40070_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _40208_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _40209_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _40210_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _40211_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _40212_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _40213_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _40214_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _40071_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _40215_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _40217_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _40218_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _40219_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _40220_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _40221_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _40222_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _40072_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39633_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39634_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39635_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39636_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39421_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39422_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39423_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39425_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39429_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39430_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39432_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39433_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39310_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39441_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39442_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39446_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39448_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39450_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39452_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39453_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39454_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39455_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39456_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39311_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39637_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39638_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39639_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39640_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39642_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39644_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39646_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39648_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39649_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39650_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39653_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39654_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39656_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39657_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39658_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39659_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39660_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39661_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39662_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39664_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39665_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39666_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39667_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39668_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39373_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39346_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39671_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39673_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39674_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39675_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39676_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39677_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39349_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39680_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39681_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39682_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39683_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39685_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39686_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39690_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39693_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39353_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39694_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39696_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39698_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39700_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39702_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39704_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39714_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39716_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39718_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39722_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39727_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39728_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39729_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39734_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39359_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39736_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39737_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39738_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39740_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39741_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39363_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39742_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39744_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39364_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39745_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39746_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39748_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39365_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39756_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39758_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39366_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _39367_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39760_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39762_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39764_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39766_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39368_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _39370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39371_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39768_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39770_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39372_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39772_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39774_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39778_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39780_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39782_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39784_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39786_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39788_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39790_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39794_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39796_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39800_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39802_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39804_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39374_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39808_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39810_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39811_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39375_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39378_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39814_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39818_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39822_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39379_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39381_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39382_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39830_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39832_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39834_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39836_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39838_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39840_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39844_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39383_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39384_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _40449_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _40469_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _40470_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _40471_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _40472_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _40473_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _40474_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _40475_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _40450_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _40451_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _40476_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _40478_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _40452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _03002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02560_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _40283_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _40369_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _40370_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _40371_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _40285_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _40286_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _40287_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _40373_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _40374_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _40375_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _40376_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _40377_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _40378_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _40379_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _40288_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _40289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19775_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19787_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19798_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08865_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08876_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08887_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08898_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06613_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13611_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13676_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12685_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _43228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _43226_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _43223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _43220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _43218_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _43216_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _43214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _43174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _43172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _43170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _43168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _43165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00176_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00177_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00179_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _43163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00183_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00185_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00187_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00188_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00190_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00192_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _43160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40913_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40915_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40923_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40931_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40938_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31040_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40944_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40946_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40948_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40952_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31062_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40962_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40963_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40965_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17370_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17381_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09470_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10669_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10713_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09491_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _41415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _41418_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41932_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41936_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41938_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _41421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41944_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41946_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41948_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41949_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41951_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41953_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _41424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _41427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _41430_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41955_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41957_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41959_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41961_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41963_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41965_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41967_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _41433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41968_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41970_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41972_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41976_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _41436_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _41439_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41982_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41984_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41989_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41991_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41993_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _41441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02129_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01627_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02171_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02175_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02177_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02179_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01642_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01226_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01230_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01232_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00574_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00552_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00558_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00563_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00566_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01238_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01240_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00568_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01244_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00576_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00579_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00582_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00584_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01260_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01262_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01268_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01285_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01287_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01291_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01304_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00598_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1071 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1071 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1071 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1071 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1073 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1075 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1075 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1076 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1076 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1077 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1077 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1078 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1078 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1079 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1079 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1080 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1080 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1081 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1118 , \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.n1146 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1147 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1147 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1147 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1147 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1147 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1147 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1148 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1148 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1148 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1148 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1148 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1148 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1149 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1149 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1149 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1149 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1149 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1149 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1149 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1150 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1151 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1152 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1152 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1152 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1153 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1154 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1154 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1155 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1155 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1155 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1155 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1155 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1155 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1181 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1181 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1181 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1181 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1181 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1181 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1181 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1181 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1181 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1181 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1181 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1181 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1181 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1183 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1183 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1183 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1183 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1183 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1183 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1185 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1185 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1185 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1185 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1185 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1185 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1185 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1189 [8], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1190 , \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1191 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1191 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1191 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1191 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1192 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1192 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1192 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1196 [4], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1197 , \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1198 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1198 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1198 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1198 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1198 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1198 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1198 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1198 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1198 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1206 , \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.n1207 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1207 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1207 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1207 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1207 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1212 , \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1217 [4], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1218 , \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1226 , \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.n1227 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1227 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1227 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1227 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1227 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1229 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1229 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1229 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1229 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1229 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1229 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1229 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1229 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1229 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1231 [8], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1232 , \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1233 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1233 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1233 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1233 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1234 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1234 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1234 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1236 [4], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1249 [8], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1257 , \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.n1258 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1258 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1258 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1258 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1258 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1260 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1262 [8], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1276 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1278 [4], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1279 , \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1280 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1280 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1280 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1280 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1280 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1280 [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1282 [8], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1290 , \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1291 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1291 [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1291 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1291 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1291 [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1292 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1292 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1292 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1292 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1292 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1295 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1295 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1295 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1295 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1295 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1295 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1295 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1295 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1295 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1296 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1296 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1296 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1296 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1296 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1296 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1297 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1297 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1297 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1297 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1297 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1297 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1297 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1297 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1298 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1299 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1299 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1299 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1299 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1299 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1299 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1299 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1299 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1300 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1300 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1303 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1305 [8], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1306 , \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1307 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1307 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1309 [4], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1310 , \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.n1318 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1318 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1318 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1318 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1318 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1322 [8], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1323 , \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.n1334 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1334 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1334 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1334 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1334 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1338 [8], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1339 , \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1350 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1350 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1354 [8], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1357 [4], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1358 , \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1365 , \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1520 , \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1521 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1521 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1521 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1521 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1521 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1521 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1521 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1680 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1683 , \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.n1691 , \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.n1692 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1692 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1692 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1692 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1692 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1696 , \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.n1698 , \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1709 , \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.n1711 , \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.n1717 , \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.n1718 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1718 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1718 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1718 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1718 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 , \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.n1724 , \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.n1730 , \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1733 , \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.n1734 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1734 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1734 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1734 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1734 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1734 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1734 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1739 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1739 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1739 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1739 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1739 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1739 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1739 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1739 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1739 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1745 , \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.n1746 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1746 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1746 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1746 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1746 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1746 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1746 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1749 , \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.n1750 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1750 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1750 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1750 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1750 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1750 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1750 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1765 , \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.n1766 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1766 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1766 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1766 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1766 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1766 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1766 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1771 , \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.n1772 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1772 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1772 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1772 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1772 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1772 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1772 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.n1778 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1778 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1778 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1778 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1778 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1778 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1778 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1783 , \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.n1784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1791 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1791 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1791 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1791 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1791 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1791 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1792 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1792 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1792 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1792 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1793 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1793 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1793 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1793 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1793 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1793 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1828 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1828 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1828 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1828 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1828 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1828 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1828 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1828 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1847 , \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.n1848 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1848 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1848 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1848 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1848 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1848 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1848 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1852 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1854 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1854 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1854 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1854 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
