
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire [15:0] _26812_;
  wire _26813_;
  wire [7:0] _26814_;
  wire [7:0] _26815_;
  wire [7:0] _26816_;
  wire [7:0] _26817_;
  wire [7:0] _26818_;
  wire [7:0] _26819_;
  wire [7:0] _26820_;
  wire [7:0] _26821_;
  wire [7:0] _26822_;
  wire [7:0] _26823_;
  wire [7:0] _26824_;
  wire [7:0] _26825_;
  wire [7:0] _26826_;
  wire [7:0] _26827_;
  wire [7:0] _26828_;
  wire [7:0] _26829_;
  wire _26830_;
  wire [7:0] _26831_;
  wire [2:0] _26832_;
  wire [2:0] _26833_;
  wire [1:0] _26834_;
  wire [7:0] _26835_;
  wire _26836_;
  wire [1:0] _26837_;
  wire [1:0] _26838_;
  wire [2:0] _26839_;
  wire [2:0] _26840_;
  wire [1:0] _26841_;
  wire [3:0] _26842_;
  wire [1:0] _26843_;
  wire _26844_;
  wire [7:0] _26845_;
  wire [7:0] _26846_;
  wire [7:0] _26847_;
  wire [7:0] _26848_;
  wire [7:0] _26849_;
  wire [7:0] _26850_;
  wire [7:0] _26851_;
  wire [7:0] _26852_;
  wire [15:0] _26853_;
  wire [15:0] _26854_;
  wire _26855_;
  wire [4:0] _26856_;
  wire [7:0] _26857_;
  wire [7:0] _26858_;
  wire _26859_;
  wire _26860_;
  wire [15:0] _26861_;
  wire [15:0] _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire [7:0] _26866_;
  wire [2:0] _26867_;
  wire [7:0] _26868_;
  wire _26869_;
  wire [7:0] _26870_;
  wire _26871_;
  wire _26872_;
  wire [3:0] _26873_;
  wire [31:0] _26874_;
  wire [31:0] _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire [15:0] _26879_;
  wire _26880_;
  wire _26881_;
  wire [7:0] _26882_;
  wire _26883_;
  wire [2:0] _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire [7:0] _27321_;
  wire _27322_;
  wire [3:0] _27323_;
  wire _27324_;
  wire _27325_;
  wire [7:0] _27326_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_22773_, rst);
  and (_22774_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_22775_, _22774_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_22776_, _22775_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_22778_, _22776_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_22779_, _22778_);
  not (_22780_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_22781_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_22782_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _22781_);
  and (_22783_, _22782_, _22780_);
  and (_22784_, _22783_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not (_22785_, _22784_);
  nor (_22786_, _22776_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_22787_, _22786_, _22785_);
  and (_22789_, _22787_, _22779_);
  not (_22790_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_22791_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _22781_);
  and (_22792_, _22791_, _22790_);
  and (_22793_, _22792_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22794_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_22795_, _22794_, _22789_);
  and (_22796_, _22792_, _22780_);
  and (_22797_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_22798_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  nor (_22799_, _22798_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22800_, _22799_, _22782_);
  and (_22801_, _22800_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_22802_, _22801_, _22797_);
  and (_22803_, _22791_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_22804_, _22803_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22805_, _22798_, _22782_);
  and (_22806_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_22807_, _22806_, _22804_);
  and (_22808_, _22807_, _22802_);
  and (_22809_, _22808_, _22795_);
  and (_22810_, _22778_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_22811_, _22810_);
  nor (_22812_, _22778_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_22813_, _22812_, _22785_);
  and (_22814_, _22813_, _22811_);
  not (_22815_, _22814_);
  and (_22816_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_22817_, _22816_, _22804_);
  and (_22818_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_22819_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor (_22820_, _22819_, _22818_);
  and (_22821_, _22820_, _22817_);
  and (_22822_, _22821_, _22815_);
  and (_22823_, _22822_, _22809_);
  and (_22824_, _22810_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_22825_, _22824_);
  nor (_22826_, _22810_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_22827_, _22826_, _22785_);
  and (_22828_, _22827_, _22825_);
  not (_22829_, _22828_);
  and (_22831_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_22832_, _22831_, _22804_);
  and (_22834_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_22835_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_22836_, _22835_, _22834_);
  and (_22837_, _22836_, _22832_);
  and (_22838_, _22837_, _22829_);
  or (_22839_, _22824_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_22840_, _22824_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_22841_, _22840_, _22784_);
  and (_22842_, _22841_, _22839_);
  not (_22844_, _22842_);
  and (_22845_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_22848_, _22845_);
  not (_22849_, _22804_);
  and (_22850_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_22851_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_22852_, _22851_, _22850_);
  and (_22853_, _22852_, _22849_);
  and (_22854_, _22853_, _22848_);
  nand (_22855_, _22854_, _22844_);
  and (_22856_, _22855_, _22838_);
  and (_22857_, _22856_, _22823_);
  and (_22859_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_22860_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_22861_, _22860_, _22859_);
  and (_22862_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not (_22863_, _22862_);
  not (_22864_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_22865_, _22784_, _22864_);
  and (_22866_, _22800_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_22867_, _22866_, _22865_);
  and (_22868_, _22867_, _22863_);
  and (_22869_, _22868_, _22861_);
  not (_22870_, _22869_);
  nor (_22871_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_22872_, _22871_, _22774_);
  and (_22873_, _22872_, _22784_);
  and (_22874_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_22875_, _22874_, _22873_);
  and (_22876_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_22877_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_22878_, _22800_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_22879_, _22878_, _22877_);
  nor (_22880_, _22879_, _22876_);
  and (_22881_, _22880_, _22875_);
  and (_22882_, _22881_, _22870_);
  nor (_22883_, _22774_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_22884_, _22883_, _22775_);
  and (_22885_, _22884_, _22784_);
  and (_22886_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_22887_, _22886_, _22885_);
  and (_22888_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_22889_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_22890_, _22800_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_22891_, _22890_, _22889_);
  nor (_22892_, _22891_, _22888_);
  and (_22894_, _22892_, _22887_);
  and (_22895_, _22894_, _22882_);
  not (_22896_, _22776_);
  nor (_22897_, _22775_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_22898_, _22785_, _22897_);
  and (_22899_, _22898_, _22896_);
  not (_22900_, _22899_);
  and (_22901_, _22800_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_22902_, _22805_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_22903_, _22902_, _22901_);
  and (_22904_, _22793_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_22905_, _22796_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_22906_, _22905_, _22904_);
  and (_22907_, _22906_, _22903_);
  and (_22908_, _22907_, _22900_);
  not (_22910_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_22912_, \oc8051_top_1.oc8051_decoder1.wr , _22781_);
  not (_22913_, _22912_);
  nor (_22914_, _22913_, _22783_);
  and (_22915_, _22914_, _22910_);
  not (_22917_, _22915_);
  nor (_22918_, _22917_, _22908_);
  and (_22920_, _22918_, _22895_);
  and (_22922_, _22920_, _22857_);
  or (_22923_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_22924_, _22923_, _22773_);
  not (_22926_, _22908_);
  and (_22927_, _22895_, _22926_);
  and (_22928_, _22857_, _22915_);
  and (_22930_, _22928_, _22927_);
  not (_22931_, _22930_);
  and (_22932_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22781_);
  and (_22933_, _22932_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_22935_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _22781_);
  and (_22937_, _22935_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_22938_, _22937_, _22933_);
  not (_22939_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_22940_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_22941_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_22942_, _22941_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_22943_, _22942_, _22940_);
  or (_22944_, _22943_, _22939_);
  nor (_22945_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_22946_, _22945_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_22947_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_22948_, _22947_, _22944_);
  nor (_22949_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_22950_, _22949_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_22951_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  not (_22952_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_22953_, _22942_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_22954_, _22953_, _22952_);
  and (_22955_, _22954_, _22951_);
  and (_22956_, _22955_, _22948_);
  nand (_22957_, _22949_, _22941_);
  not (_22958_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_22959_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _22958_);
  or (_22960_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  not (_22961_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_22962_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _22961_);
  and (_22963_, _22962_, _22960_);
  or (_22964_, _22963_, _22959_);
  nand (_22965_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _22958_);
  or (_22966_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_22967_, _22966_, _22964_);
  or (_22968_, _22967_, _22957_);
  and (_22969_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_22970_, _22969_, _22940_);
  nand (_22971_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_22972_, _22969_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_22973_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_22974_, _22973_, _22971_);
  and (_22975_, _22974_, _22968_);
  and (_22976_, _22975_, _22956_);
  not (_22977_, _22976_);
  or (_22978_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_22979_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _22961_);
  and (_22980_, _22979_, _22978_);
  or (_22981_, _22980_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_22982_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  or (_22983_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_22984_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _22961_);
  and (_22986_, _22984_, _22983_);
  or (_22987_, _22986_, _22982_);
  not (_22988_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_22989_, _22988_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_22990_, _22989_, _22987_);
  nand (_22991_, _22990_, _22981_);
  not (_22992_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_22993_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _22992_);
  or (_22994_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_22995_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _22961_);
  and (_22996_, _22995_, _22994_);
  nand (_22997_, _22996_, _22982_);
  or (_22998_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_22999_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _22961_);
  and (_23000_, _22999_, _22998_);
  nand (_23002_, _23000_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23003_, _23002_, _22997_);
  nand (_23004_, _23003_, _22993_);
  or (_23005_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_23006_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _22961_);
  and (_23007_, _23006_, _23005_);
  not (_23008_, _23007_);
  and (_23009_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_23010_, _23009_, _22982_);
  or (_23011_, _23010_, _23008_);
  or (_23012_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_23013_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _22961_);
  and (_23014_, _23013_, _23012_);
  nor (_23015_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23016_, _23015_, _22982_);
  nand (_23017_, _23016_, _23014_);
  and (_23019_, _23017_, _23011_);
  and (_23020_, _23015_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23021_, _23020_, _22963_);
  or (_23023_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or (_23024_, _22961_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_23025_, _23024_, _23023_);
  not (_23026_, _23025_);
  nand (_23028_, _23009_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  or (_23029_, _23028_, _23026_);
  and (_23030_, _23029_, _23021_);
  and (_23032_, _23030_, _23019_);
  and (_23033_, _23032_, _23004_);
  nand (_23034_, _23033_, _22991_);
  nand (_23035_, _23034_, _22965_);
  and (_23036_, _22959_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_23037_, _23036_);
  and (_23038_, _23037_, _23035_);
  and (_23039_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_23040_, _23039_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_23041_, _23040_, _23038_);
  not (_23043_, _23040_);
  and (_23044_, _23043_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_23045_, _23044_);
  and (_23046_, _23045_, _23041_);
  and (_23047_, _23046_, _22977_);
  nand (_23048_, _23045_, _23041_);
  or (_23050_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_23051_, _23050_, _22967_);
  and (_23053_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nand (_23054_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_23055_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_23056_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_23057_, _23056_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_23058_, _23057_, _23055_);
  and (_23059_, _23058_, _23054_);
  nand (_23060_, _23059_, _23051_);
  and (_23061_, _23060_, _23048_);
  or (_23062_, _23061_, _23047_);
  and (_23063_, _23062_, _22938_);
  not (_23064_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23065_, _22932_, _23064_);
  and (_23067_, _23065_, _22937_);
  nand (_23068_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_23071_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_23073_, _22943_, _23071_);
  and (_23074_, _23073_, _23068_);
  nand (_23076_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand (_23077_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_23079_, _23077_, _23076_);
  and (_23080_, _23079_, _23074_);
  or (_23082_, _23007_, _22959_);
  or (_23083_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_23084_, _23083_, _23082_);
  or (_23085_, _23084_, _22957_);
  not (_23086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_23087_, _22953_, _23086_);
  nand (_23088_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_23089_, _23088_, _23087_);
  and (_23090_, _23089_, _23085_);
  and (_23091_, _23090_, _23080_);
  not (_23092_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_23093_, _22943_, _23092_);
  and (_23094_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_23095_, _23094_, _23093_);
  and (_23096_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not (_23097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_23098_, _22953_, _23097_);
  nor (_23099_, _23098_, _23096_);
  and (_23100_, _23099_, _23095_);
  or (_23101_, _23014_, _22959_);
  or (_23102_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_23103_, _23102_, _23101_);
  or (_23104_, _23103_, _22957_);
  and (_23105_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_23106_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_23107_, _23106_, _23105_);
  and (_23108_, _23107_, _23104_);
  and (_23109_, _23108_, _23100_);
  nand (_23110_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand (_23111_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_23112_, _23111_, _23110_);
  not (_23114_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_23115_, _22943_, _23114_);
  nand (_23116_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_23117_, _23116_, _23115_);
  and (_23118_, _23117_, _23112_);
  or (_23119_, _22980_, _22959_);
  or (_23120_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_23121_, _23120_, _23119_);
  or (_23122_, _23121_, _22957_);
  not (_23123_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_23124_, _22953_, _23123_);
  nand (_23125_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_23126_, _23125_, _23124_);
  and (_23127_, _23126_, _23122_);
  nand (_23128_, _23127_, _23118_);
  not (_23129_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_23130_, _22943_, _23129_);
  nand (_23131_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_23132_, _23131_, _23130_);
  not (_23133_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_23134_, _22953_, _23133_);
  nand (_23135_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_23136_, _23135_, _23134_);
  and (_23137_, _23136_, _23132_);
  or (_23138_, _22996_, _22959_);
  or (_23139_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_23140_, _23139_, _23138_);
  or (_23142_, _23140_, _22957_);
  nand (_23143_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand (_23144_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_23145_, _23144_, _23143_);
  and (_23146_, _23145_, _23142_);
  nand (_23147_, _23146_, _23137_);
  nor (_23148_, _23147_, _23128_);
  and (_23149_, _23148_, _23109_);
  and (_23150_, _23149_, _23091_);
  nand (_23151_, _23150_, _23048_);
  not (_23152_, _23091_);
  not (_23153_, _23109_);
  and (_23154_, _23147_, _23153_);
  and (_23155_, _23154_, _23128_);
  and (_23156_, _23155_, _23152_);
  nand (_23157_, _23156_, _23046_);
  and (_23158_, _23157_, _23151_);
  or (_23159_, _23158_, _22976_);
  nand (_23160_, _23158_, _22976_);
  and (_23161_, _23160_, _23159_);
  and (_23162_, _23161_, _23067_);
  nor (_23163_, _23162_, _23063_);
  not (_23164_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not (_23165_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_23166_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _22781_);
  and (_23167_, _23166_, _23165_);
  and (_23168_, _23167_, _23164_);
  and (_23169_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _22781_);
  nor (_23170_, _23166_, _22935_);
  and (_23171_, _23170_, _23169_);
  nor (_23172_, _23169_, _22932_);
  and (_23173_, _23172_, _23170_);
  or (_23174_, _23173_, _23171_);
  nor (_23175_, _23174_, _23168_);
  and (_23176_, _22937_, _23164_);
  not (_23177_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23178_, _22935_, _23177_);
  and (_23179_, _23178_, _22932_);
  nor (_23180_, _23179_, _23176_);
  and (_23181_, _23180_, _23175_);
  nor (_23182_, _23181_, _22976_);
  not (_23183_, _23182_);
  and (_23184_, _23178_, _23172_);
  and (_23185_, _23059_, _23051_);
  nor (_23186_, _23185_, _22976_);
  and (_23187_, _23185_, _22976_);
  nor (_23188_, _23187_, _23186_);
  and (_23189_, _23188_, _23184_);
  not (_23190_, _23189_);
  and (_23191_, _23169_, _23164_);
  and (_23192_, _23178_, _23191_);
  not (_23193_, _23192_);
  nor (_23194_, _23193_, _23187_);
  not (_23195_, _23194_);
  and (_23196_, _23167_, _22933_);
  and (_23197_, _23196_, _23186_);
  and (_23198_, _23167_, _23065_);
  and (_23199_, _23198_, _22976_);
  nor (_23200_, _23199_, _23197_);
  and (_23201_, _23200_, _23195_);
  and (_23202_, _23201_, _23190_);
  and (_23204_, _23202_, _23183_);
  nand (_23205_, _23204_, _23163_);
  or (_23206_, _23205_, _22931_);
  and (_22846_, _23206_, _22924_);
  not (_23207_, _22894_);
  and (_23208_, _23207_, _22882_);
  and (_23209_, _23208_, _22918_);
  and (_23210_, _23209_, _22857_);
  not (_23211_, _23210_);
  or (_23212_, _23121_, _23050_);
  nand (_23213_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_23214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_23215_, _23057_, _23214_);
  and (_23216_, _23215_, _23213_);
  nand (_23217_, _23216_, _23212_);
  and (_23218_, _23217_, _22938_);
  nor (_23219_, _23154_, _23048_);
  not (_23220_, _23147_);
  and (_23221_, _23220_, _23109_);
  nor (_23222_, _23221_, _23046_);
  nor (_23223_, _23222_, _23219_);
  nand (_23224_, _23223_, _23128_);
  or (_23225_, _23223_, _23128_);
  and (_23226_, _23225_, _23067_);
  and (_23228_, _23226_, _23224_);
  nor (_23229_, _23228_, _23218_);
  not (_23230_, _23181_);
  and (_23231_, _23230_, _23128_);
  not (_23232_, _23231_);
  and (_23233_, _23217_, _23128_);
  nor (_23234_, _23217_, _23128_);
  nor (_23235_, _23234_, _23233_);
  and (_23236_, _23235_, _23184_);
  not (_23237_, _23236_);
  nor (_23238_, _23234_, _23193_);
  not (_23239_, _23238_);
  and (_23240_, _23233_, _23196_);
  not (_23241_, _23128_);
  and (_23242_, _23198_, _23241_);
  nor (_23243_, _23242_, _23240_);
  and (_23244_, _23243_, _23239_);
  and (_23245_, _23244_, _23237_);
  and (_23246_, _23245_, _23232_);
  nand (_23247_, _23246_, _23229_);
  or (_23248_, _23247_, _23211_);
  nor (_23249_, _22881_, _22869_);
  and (_23250_, _23249_, _22894_);
  and (_23251_, _23250_, _22918_);
  and (_23252_, _23251_, _22857_);
  not (_23253_, _23252_);
  not (_23254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  not (_23255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_23256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_23257_, _23256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not (_23258_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_23259_, t1_i);
  and (_23260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _23259_);
  nor (_23261_, _23260_, _23258_);
  not (_23262_, _23261_);
  not (_23263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_23264_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _23263_);
  nor (_23265_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_23266_, _23265_);
  and (_23267_, _23266_, _23264_);
  and (_23268_, _23267_, _23262_);
  and (_23269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_23270_, _23269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_23271_, _23270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_23272_, _23271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_23273_, _23272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_23274_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_23275_, _23274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_23276_, _23275_, _23268_);
  and (_23277_, _23276_, _23257_);
  and (_23278_, _23277_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_23279_, _23268_, _23256_);
  not (_23280_, _23257_);
  and (_23281_, _23272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_23282_, _23281_, _23280_);
  and (_23283_, _23282_, _23279_);
  nor (_23284_, _23283_, _23278_);
  nor (_23285_, _23284_, _23255_);
  nor (_23286_, _23285_, _23254_);
  and (_23287_, _23285_, _23254_);
  or (_23288_, _23287_, _23286_);
  or (_23289_, _23210_, _23288_);
  and (_23290_, _23289_, _23253_);
  and (_23291_, _23290_, _23248_);
  and (_23292_, _23252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_23293_, _23292_, _23291_);
  and (_23069_, _23293_, _22773_);
  or (_23294_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_23295_, _23294_, _22773_);
  not (_23296_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_23297_, _22943_, _23296_);
  nand (_23298_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_23299_, _23298_, _23297_);
  not (_23300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_23301_, _22953_, _23300_);
  nand (_23302_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_23303_, _23302_, _23301_);
  and (_23304_, _23303_, _23299_);
  or (_23305_, _23000_, _22959_);
  or (_23306_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_23307_, _23306_, _23305_);
  or (_23308_, _23307_, _22957_);
  nand (_23309_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_23310_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_23311_, _23310_, _23309_);
  and (_23312_, _23311_, _23308_);
  nand (_23313_, _23312_, _23304_);
  not (_23314_, _23313_);
  and (_23315_, _23314_, _23046_);
  not (_23316_, _22938_);
  or (_23317_, _23307_, _23050_);
  nand (_23318_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not (_23319_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_23321_, _23057_, _23319_);
  and (_23322_, _23321_, _23318_);
  and (_23323_, _23322_, _23317_);
  and (_23324_, _23323_, _23048_);
  or (_23325_, _23324_, _23316_);
  nor (_23326_, _23325_, _23315_);
  and (_23327_, _23156_, _22977_);
  nor (_23328_, _23327_, _23048_);
  and (_23330_, _23150_, _22976_);
  nor (_23331_, _23330_, _23046_);
  nor (_23332_, _23331_, _23328_);
  nor (_23333_, _23332_, _23313_);
  not (_23335_, _23067_);
  and (_23336_, _23332_, _23313_);
  or (_23337_, _23336_, _23335_);
  nor (_23338_, _23337_, _23333_);
  nor (_23340_, _23338_, _23326_);
  and (_23341_, _23313_, _23230_);
  not (_23342_, _23341_);
  nand (_23343_, _23322_, _23317_);
  and (_23344_, _23313_, _23343_);
  nor (_23345_, _23313_, _23343_);
  nor (_23346_, _23345_, _23344_);
  and (_23347_, _23346_, _23184_);
  not (_23348_, _23347_);
  nor (_23349_, _23345_, _23193_);
  not (_23350_, _23349_);
  and (_23351_, _23344_, _23196_);
  and (_23352_, _23314_, _23198_);
  nor (_23353_, _23352_, _23351_);
  and (_23354_, _23353_, _23350_);
  and (_23355_, _23354_, _23348_);
  and (_23356_, _23355_, _23342_);
  and (_23357_, _23356_, _23340_);
  nand (_23359_, _23357_, _22930_);
  and (_26609_, _23359_, _23295_);
  and (_23360_, _23275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_23361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_23362_, _23361_, _23268_);
  and (_23363_, _23362_, _23360_);
  nand (_23364_, _23363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_23365_, _23363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_23366_, _23365_, _23257_);
  and (_23367_, _23366_, _23364_);
  and (_23368_, _23281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_23370_, _23368_, _23268_);
  and (_23371_, _23370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_23372_, _23371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_23373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not (_23374_, _23373_);
  and (_23375_, _23371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_23376_, _23375_, _23374_);
  and (_23377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_23378_, _23377_, _23376_);
  and (_23379_, _23378_, _23372_);
  or (_23380_, _23379_, _23367_);
  or (_23381_, _23380_, _23210_);
  or (_23383_, _23084_, _23050_);
  nand (_23384_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not (_23385_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_23386_, _23057_, _23385_);
  and (_23387_, _23386_, _23384_);
  nand (_23388_, _23387_, _23383_);
  and (_23389_, _23388_, _22938_);
  or (_23390_, _23149_, _23046_);
  or (_23391_, _23155_, _23048_);
  and (_23392_, _23391_, _23390_);
  nand (_23393_, _23392_, _23152_);
  or (_23394_, _23392_, _23152_);
  and (_23395_, _23394_, _23067_);
  and (_23396_, _23395_, _23393_);
  nor (_23397_, _23396_, _23389_);
  and (_23398_, _23387_, _23383_);
  nor (_23399_, _23398_, _23091_);
  and (_23400_, _23399_, _23196_);
  and (_23401_, _23198_, _23091_);
  nor (_23402_, _23401_, _23400_);
  nor (_23403_, _23181_, _23091_);
  and (_23404_, _23398_, _23091_);
  nor (_23405_, _23404_, _23193_);
  not (_23406_, _23184_);
  or (_23407_, _23399_, _23404_);
  nor (_23408_, _23407_, _23406_);
  or (_23409_, _23408_, _23405_);
  nor (_23411_, _23409_, _23403_);
  and (_23412_, _23411_, _23402_);
  nand (_23413_, _23412_, _23397_);
  or (_23414_, _23413_, _23211_);
  and (_23415_, _23414_, _23381_);
  or (_23416_, _23415_, _23252_);
  or (_23417_, _23253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_23418_, _23417_, _22773_);
  and (_00001_, _23418_, _23416_);
  nor (_23419_, _22855_, _22910_);
  and (_23420_, _23419_, _22926_);
  nor (_23421_, _22869_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23422_, _23421_, _23420_);
  and (_23423_, _22853_, _22912_);
  not (_23424_, _23423_);
  nor (_23425_, _23424_, _23422_);
  not (_23426_, _22809_);
  and (_23427_, _23419_, _23426_);
  nor (_23428_, _22881_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23429_, _23428_, _23427_);
  nor (_23431_, _23429_, _23424_);
  and (_23432_, _23431_, _23425_);
  not (_23433_, _22838_);
  and (_23434_, _23419_, _23433_);
  nor (_23435_, _23419_, _22908_);
  nor (_23436_, _23435_, _23434_);
  nor (_23437_, _23436_, _23424_);
  not (_23439_, _22822_);
  and (_23440_, _23419_, _23439_);
  nor (_23441_, _22894_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23442_, _23441_, _23440_);
  and (_23443_, _23442_, _23437_);
  and (_23444_, _23443_, _23432_);
  nor (_23445_, _23419_, _23439_);
  nor (_23446_, _23445_, _23424_);
  nor (_23447_, _23419_, _22809_);
  not (_23448_, _23447_);
  and (_23449_, _23448_, _23446_);
  nor (_23450_, _22855_, _23433_);
  nor (_23451_, _23450_, _23419_);
  not (_23452_, _23451_);
  and (_23453_, _23452_, _23449_);
  and (_23454_, _23453_, _23444_);
  and (_23455_, _22982_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23456_, _23455_, _22989_);
  and (_23458_, _23170_, _23065_);
  not (_23459_, _23458_);
  not (_23460_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_23461_, _22943_, _23460_);
  nand (_23462_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_23463_, _23462_, _23461_);
  not (_23464_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or (_23465_, _22953_, _23464_);
  nand (_23466_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_23467_, _23466_, _23465_);
  and (_23468_, _23467_, _23463_);
  or (_23469_, _23025_, _22959_);
  or (_23470_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_23471_, _23470_, _23469_);
  or (_23472_, _23471_, _22957_);
  nand (_23474_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand (_23475_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_23476_, _23475_, _23474_);
  and (_23478_, _23476_, _23472_);
  and (_23479_, _23478_, _23468_);
  or (_23480_, _23471_, _23050_);
  and (_23481_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_23482_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_23483_, _23057_, _23482_);
  nor (_23484_, _23483_, _23481_);
  and (_23485_, _23484_, _23480_);
  not (_23487_, _23485_);
  and (_23488_, _23487_, _23479_);
  nor (_23489_, _23485_, _23479_);
  and (_23490_, _23485_, _23479_);
  nor (_23492_, _23490_, _23489_);
  not (_23493_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_23494_, _22943_, _23493_);
  nand (_23495_, _22946_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_23496_, _23495_, _23494_);
  nand (_23497_, _22950_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_23498_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_23499_, _22953_, _23498_);
  and (_23501_, _23499_, _23497_);
  and (_23502_, _23501_, _23496_);
  or (_23503_, _22986_, _22959_);
  or (_23504_, _22965_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_23505_, _23504_, _23503_);
  or (_23506_, _23505_, _22957_);
  nand (_23507_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_23508_, _22972_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_23509_, _23508_, _23507_);
  and (_23510_, _23509_, _23506_);
  and (_23511_, _23510_, _23502_);
  or (_23512_, _23505_, _23050_);
  nand (_23513_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_23514_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_23515_, _23057_, _23514_);
  and (_23516_, _23515_, _23513_);
  nand (_23518_, _23516_, _23512_);
  nor (_23519_, _23518_, _23511_);
  not (_23520_, _23518_);
  nor (_23521_, _23520_, _23511_);
  and (_23522_, _23520_, _23511_);
  nor (_23523_, _23522_, _23521_);
  and (_23524_, _23313_, _23323_);
  and (_23525_, _23060_, _22976_);
  nor (_23526_, _23346_, _23525_);
  nor (_23527_, _23526_, _23524_);
  nor (_23528_, _23527_, _23523_);
  nor (_23529_, _23528_, _23519_);
  and (_23530_, _23527_, _23523_);
  nor (_23531_, _23530_, _23528_);
  not (_23532_, _23531_);
  and (_23533_, _23346_, _23525_);
  nor (_23534_, _23533_, _23526_);
  not (_23535_, _23534_);
  not (_23536_, _23188_);
  not (_23537_, _23407_);
  and (_23538_, _23216_, _23212_);
  and (_23539_, _23538_, _23128_);
  or (_23540_, _23140_, _23050_);
  nand (_23541_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not (_23542_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_23543_, _23057_, _23542_);
  and (_23544_, _23543_, _23541_);
  nand (_23545_, _23544_, _23540_);
  and (_23546_, _23545_, _23147_);
  nor (_23547_, _23545_, _23147_);
  nor (_23548_, _23547_, _23546_);
  or (_23549_, _23103_, _23050_);
  nand (_23550_, _23053_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not (_23551_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_23552_, _23057_, _23551_);
  and (_23553_, _23552_, _23550_);
  nand (_23554_, _23553_, _23549_);
  and (_23555_, _23554_, _23109_);
  nor (_23557_, _23555_, _23548_);
  not (_23558_, _23545_);
  and (_23559_, _23558_, _23147_);
  nor (_23560_, _23559_, _23557_);
  nor (_23561_, _23560_, _23235_);
  nor (_23562_, _23561_, _23539_);
  nor (_23563_, _23562_, _23537_);
  and (_23564_, _23562_, _23537_);
  nor (_23565_, _23564_, _23563_);
  not (_23566_, _23565_);
  and (_23567_, _23560_, _23235_);
  nor (_23568_, _23567_, _23561_);
  not (_23569_, _23568_);
  not (_23570_, _23554_);
  nor (_23571_, _23570_, _23109_);
  and (_23572_, _23570_, _23109_);
  nor (_23573_, _23572_, _23571_);
  not (_23575_, _23573_);
  and (_23576_, _23575_, _23048_);
  and (_23577_, _23555_, _23548_);
  nor (_23578_, _23577_, _23557_);
  not (_23579_, _23578_);
  and (_23580_, _23579_, _23576_);
  and (_23581_, _23580_, _23569_);
  and (_23582_, _23581_, _23566_);
  or (_23583_, _23388_, _23091_);
  and (_23584_, _23388_, _23091_);
  or (_23585_, _23562_, _23584_);
  and (_23586_, _23585_, _23583_);
  or (_23587_, _23586_, _23582_);
  and (_23588_, _23587_, _23536_);
  and (_23589_, _23588_, _23535_);
  and (_23590_, _23589_, _23532_);
  nor (_23591_, _23590_, _23529_);
  nor (_23593_, _23591_, _23492_);
  nor (_23594_, _23593_, _23488_);
  nor (_23595_, _23594_, _23459_);
  not (_23596_, _23595_);
  and (_23597_, _23191_, _23170_);
  not (_23598_, _23597_);
  not (_23599_, _23489_);
  not (_23600_, _23235_);
  and (_23601_, _23571_, _23548_);
  nor (_23602_, _23601_, _23546_);
  nor (_23603_, _23602_, _23600_);
  nor (_23604_, _23603_, _23233_);
  nor (_23605_, _23604_, _23537_);
  and (_23606_, _23604_, _23537_);
  nor (_23607_, _23606_, _23605_);
  and (_23608_, _23573_, _23048_);
  and (_23610_, _23608_, _23548_);
  and (_23611_, _23602_, _23600_);
  nor (_23612_, _23611_, _23603_);
  and (_23613_, _23612_, _23610_);
  not (_23614_, _23613_);
  nor (_23615_, _23614_, _23607_);
  nor (_23616_, _23604_, _23404_);
  or (_23617_, _23616_, _23399_);
  or (_23618_, _23617_, _23615_);
  and (_23620_, _23618_, _23188_);
  and (_23621_, _23620_, _23346_);
  not (_23622_, _23523_);
  and (_23623_, _23346_, _23186_);
  nor (_23624_, _23623_, _23344_);
  nor (_23625_, _23624_, _23622_);
  and (_23626_, _23624_, _23622_);
  nor (_23627_, _23626_, _23625_);
  and (_23628_, _23627_, _23621_);
  not (_23629_, _23628_);
  nor (_23630_, _23625_, _23521_);
  and (_23631_, _23630_, _23629_);
  or (_23632_, _23631_, _23490_);
  and (_23633_, _23632_, _23599_);
  nor (_23634_, _23633_, _23598_);
  and (_23635_, _23178_, _22933_);
  not (_23636_, _23479_);
  and (_23637_, _23636_, _23635_);
  not (_23638_, _23637_);
  and (_23639_, _23191_, _23167_);
  nor (_23640_, _23148_, _23091_);
  and (_23641_, _23640_, _23639_);
  and (_23642_, _23191_, _22937_);
  and (_23643_, _23642_, _23153_);
  nor (_23644_, _23643_, _23641_);
  and (_23645_, _23644_, _23638_);
  nand (_23647_, _23173_, _23048_);
  and (_23648_, _23647_, _23645_);
  and (_23649_, _23045_, _23038_);
  and (_23650_, _23184_, _23041_);
  nor (_23651_, _23650_, _23192_);
  nor (_23652_, _23651_, _23649_);
  and (_23653_, _23641_, _22977_);
  nor (_23654_, _23653_, _23313_);
  and (_23655_, _23654_, _23511_);
  nor (_23656_, _23655_, _23479_);
  or (_23657_, _23656_, _23048_);
  and (_23658_, _23636_, _23048_);
  not (_23659_, _23658_);
  or (_23660_, _23659_, _23655_);
  and (_23661_, _23660_, _23639_);
  and (_23662_, _23661_, _23657_);
  and (_23663_, _23172_, _22937_);
  and (_23664_, _23663_, _23038_);
  and (_23665_, _23664_, _23048_);
  and (_23666_, _23198_, _23046_);
  or (_23667_, _23666_, _23665_);
  nand (_23668_, _23037_, _23035_);
  and (_23669_, _23040_, _23668_);
  and (_23670_, _23178_, _23065_);
  and (_23671_, _23196_, _23668_);
  nor (_23672_, _23671_, _23670_);
  nor (_23673_, _23672_, _23669_);
  or (_23675_, _23673_, _23667_);
  or (_23676_, _23675_, _23662_);
  nor (_23677_, _23676_, _23652_);
  and (_23678_, _23677_, _23648_);
  not (_23679_, _23678_);
  nor (_23680_, _23679_, _23634_);
  and (_23681_, _23680_, _23596_);
  nor (_23682_, _23681_, _23456_);
  and (_23683_, _23247_, _22910_);
  and (_23685_, _23455_, _22992_);
  and (_23686_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23687_, _23455_, _23009_);
  or (_23688_, _23687_, _23686_);
  or (_23689_, _23688_, _23685_);
  and (_23690_, _23689_, _22980_);
  or (_23691_, _23690_, _23683_);
  or (_23692_, _23691_, _23682_);
  and (_23693_, _23692_, _23423_);
  and (_23694_, _23693_, _23454_);
  not (_23695_, _23454_);
  and (_23696_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or (_01943_, _23696_, _23694_);
  and (_23697_, _23429_, _23425_);
  nor (_23698_, _23442_, _23424_);
  nor (_23699_, _23698_, _23437_);
  and (_23700_, _23699_, _23697_);
  and (_23701_, _23447_, _23423_);
  and (_23702_, _23701_, _23446_);
  nor (_23703_, _23419_, _22838_);
  nor (_23704_, _22855_, _22913_);
  and (_23705_, _23704_, _23703_);
  and (_23706_, _23705_, _23702_);
  and (_23707_, _23706_, _23700_);
  not (_23708_, _23681_);
  and (_23709_, _23687_, _23708_);
  and (_23710_, _23413_, _22910_);
  and (_23711_, _23010_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23712_, _23711_, _23007_);
  or (_23713_, _23712_, _23710_);
  or (_23714_, _23713_, _23709_);
  and (_23715_, _23714_, _23423_);
  and (_23716_, _23715_, _23707_);
  not (_23717_, _23707_);
  and (_23718_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_02308_, _23718_, _23716_);
  and (_23719_, _23702_, _22856_);
  and (_23721_, _23719_, _23700_);
  and (_23722_, _23721_, _23693_);
  not (_23723_, _23721_);
  and (_23724_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_02806_, _23724_, _23722_);
  nand (_23725_, _23455_, _22993_);
  nor (_23726_, _23725_, _23681_);
  and (_23727_, _23230_, _23147_);
  and (_23728_, _23545_, _22938_);
  nor (_23729_, _23154_, _23221_);
  nand (_23730_, _23729_, _23048_);
  or (_23731_, _23729_, _23048_);
  and (_23732_, _23731_, _23067_);
  and (_23733_, _23732_, _23730_);
  nor (_23734_, _23733_, _23728_);
  and (_23735_, _23546_, _23196_);
  and (_23736_, _23198_, _23220_);
  nor (_23737_, _23736_, _23735_);
  and (_23738_, _23548_, _23184_);
  nor (_23739_, _23547_, _23193_);
  or (_23740_, _23739_, _23738_);
  not (_23741_, _23740_);
  and (_23742_, _23741_, _23737_);
  nand (_23743_, _23742_, _23734_);
  or (_23744_, _23743_, _23727_);
  and (_23745_, _23744_, _22910_);
  and (_23746_, _23455_, _22988_);
  or (_23747_, _23746_, _23688_);
  and (_23748_, _23747_, _22996_);
  or (_23749_, _23748_, _23745_);
  or (_23750_, _23749_, _23726_);
  and (_23751_, _23750_, _23423_);
  and (_23752_, _23751_, _23721_);
  and (_23753_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_03081_, _23753_, _23752_);
  and (_23754_, _23751_, _23454_);
  and (_23755_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or (_03266_, _23755_, _23754_);
  not (_23756_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_23757_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_23758_, _23757_, _23756_);
  nor (_23759_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_23760_, _23759_, _22781_);
  and (_23761_, _23760_, _23758_);
  and (_23763_, _23761_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_23764_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_23765_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_23766_, _23763_, _23765_);
  or (_23767_, _23766_, _23764_);
  and (_26853_[0], _23767_, _22773_);
  and (_23768_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_23769_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_23770_, _23763_, _23769_);
  or (_23771_, _23770_, _23768_);
  and (_26853_[1], _23771_, _22773_);
  and (_23772_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_23774_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_23775_, _23763_, _23774_);
  or (_23776_, _23775_, _23772_);
  and (_26853_[2], _23776_, _22773_);
  and (_23777_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_23778_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_23779_, _23763_, _23778_);
  or (_23780_, _23779_, _23777_);
  and (_26853_[3], _23780_, _22773_);
  and (_23781_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_23782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_23783_, _23763_, _23782_);
  or (_23784_, _23783_, _23781_);
  and (_26853_[4], _23784_, _22773_);
  and (_23785_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_23786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_23787_, _23763_, _23786_);
  or (_23788_, _23787_, _23785_);
  and (_26853_[5], _23788_, _22773_);
  and (_23789_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_23790_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_23791_, _23763_, _23790_);
  or (_23792_, _23791_, _23789_);
  and (_26853_[6], _23792_, _22773_);
  and (_23793_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_23794_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_23795_, _23763_, _23794_);
  or (_23796_, _23795_, _23793_);
  and (_26853_[7], _23796_, _22773_);
  and (_23797_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_23798_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_23799_, _23763_, _23798_);
  or (_23800_, _23799_, _23797_);
  and (_26853_[8], _23800_, _22773_);
  and (_23801_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_23802_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_23803_, _23763_, _23802_);
  or (_23804_, _23803_, _23801_);
  and (_26853_[9], _23804_, _22773_);
  and (_23805_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_23806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_23808_, _23763_, _23806_);
  or (_23809_, _23808_, _23805_);
  and (_26853_[10], _23809_, _22773_);
  and (_23810_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_23811_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_23812_, _23763_, _23811_);
  or (_23813_, _23812_, _23810_);
  and (_26853_[11], _23813_, _22773_);
  and (_23814_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_23816_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_23817_, _23763_, _23816_);
  or (_23818_, _23817_, _23814_);
  and (_26853_[12], _23818_, _22773_);
  and (_23819_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_23820_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_23821_, _23763_, _23820_);
  or (_23822_, _23821_, _23819_);
  and (_26853_[13], _23822_, _22773_);
  and (_23823_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_23824_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_23825_, _23763_, _23824_);
  or (_23827_, _23825_, _23823_);
  and (_26853_[14], _23827_, _22773_);
  and (_23828_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_23830_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23831_, _23763_, _23830_);
  or (_23832_, _23831_, _23828_);
  and (_26854_[0], _23832_, _22773_);
  and (_23833_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_23835_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_23836_, _23763_, _23835_);
  or (_23837_, _23836_, _23833_);
  and (_26854_[1], _23837_, _22773_);
  and (_23839_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_23840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_23841_, _23763_, _23840_);
  or (_23842_, _23841_, _23839_);
  and (_26854_[2], _23842_, _22773_);
  and (_23843_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_23844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_23845_, _23763_, _23844_);
  or (_23846_, _23845_, _23843_);
  and (_26854_[3], _23846_, _22773_);
  or (_23847_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand (_23848_, _23763_, _23782_);
  and (_23849_, _23848_, _22773_);
  and (_26854_[4], _23849_, _23847_);
  and (_23850_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_23851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_23852_, _23763_, _23851_);
  or (_23853_, _23852_, _23850_);
  and (_26854_[5], _23853_, _22773_);
  and (_23854_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_23855_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_23856_, _23763_, _23855_);
  or (_23858_, _23856_, _23854_);
  and (_26854_[6], _23858_, _22773_);
  and (_23859_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_23860_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_23861_, _23763_, _23860_);
  or (_23862_, _23861_, _23859_);
  and (_26854_[7], _23862_, _22773_);
  or (_23863_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand (_23864_, _23763_, _23798_);
  and (_23865_, _23864_, _22773_);
  and (_26854_[8], _23865_, _23863_);
  and (_23866_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not (_23867_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_23868_, _23763_, _23867_);
  or (_23869_, _23868_, _23866_);
  and (_26854_[9], _23869_, _22773_);
  or (_23870_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nand (_23871_, _23763_, _23806_);
  and (_23872_, _23871_, _22773_);
  and (_26854_[10], _23872_, _23870_);
  and (_23873_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_23874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_23875_, _23763_, _23874_);
  or (_23876_, _23875_, _23873_);
  and (_26854_[11], _23876_, _22773_);
  and (_23877_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  not (_23878_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_23879_, _23763_, _23878_);
  or (_23880_, _23879_, _23877_);
  and (_26854_[12], _23880_, _22773_);
  or (_23881_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nand (_23882_, _23763_, _23820_);
  and (_23883_, _23882_, _22773_);
  and (_26854_[13], _23883_, _23881_);
  and (_23884_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  not (_23885_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_23886_, _23763_, _23885_);
  or (_23887_, _23886_, _23884_);
  and (_26854_[14], _23887_, _22773_);
  nor (_23888_, _23431_, _23425_);
  and (_23889_, _23698_, _23436_);
  and (_23890_, _23889_, _23888_);
  and (_23891_, _23702_, _23452_);
  and (_23892_, _23891_, _23890_);
  nand (_23893_, _23686_, _23015_);
  nor (_23894_, _23893_, _23681_);
  and (_23895_, _23205_, _22910_);
  nand (_23896_, _22963_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23897_, _23896_, _23020_);
  or (_23898_, _23897_, _23895_);
  or (_23899_, _23898_, _23894_);
  and (_23900_, _23899_, _23423_);
  and (_23901_, _23900_, _23892_);
  not (_23902_, _23892_);
  and (_23903_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or (_22706_, _23903_, _23901_);
  and (_23904_, _23698_, _23437_);
  and (_23905_, _23904_, _23888_);
  and (_23906_, _23701_, _22822_);
  and (_23907_, _22855_, _23433_);
  and (_23909_, _23907_, _23906_);
  and (_23910_, _23909_, _23905_);
  nand (_23911_, _23686_, _22993_);
  nor (_23912_, _23911_, _23681_);
  nor (_23913_, _23357_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23914_, _22993_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_23915_, _23000_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23917_, _23915_, _23914_);
  or (_23918_, _23917_, _23913_);
  or (_23919_, _23918_, _23912_);
  and (_23920_, _23919_, _23423_);
  and (_23921_, _23920_, _23910_);
  not (_23922_, _23910_);
  and (_23923_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_22718_, _23923_, _23921_);
  and (_23924_, _23904_, _23432_);
  and (_23925_, _23924_, _23891_);
  and (_23926_, _23925_, _23920_);
  not (_23927_, _23925_);
  and (_23928_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_22733_, _23928_, _23926_);
  and (_23929_, _23431_, _23422_);
  and (_23930_, _23929_, _23443_);
  and (_23932_, _23930_, _23453_);
  and (_23933_, _23932_, _23920_);
  not (_23934_, _23932_);
  and (_23935_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_22858_, _23935_, _23933_);
  and (_23936_, _23910_, _23715_);
  and (_23937_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_22911_, _23937_, _23936_);
  and (_23938_, _23888_, _23699_);
  and (_23939_, _23938_, _23719_);
  and (_23940_, _23939_, _23693_);
  not (_23941_, _23939_);
  and (_23942_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or (_23070_, _23942_, _23940_);
  and (_23943_, _23686_, _23009_);
  and (_23944_, _23943_, _23708_);
  and (_23945_, _23511_, _23314_);
  and (_23946_, _23945_, _23330_);
  nor (_23948_, _23946_, _23046_);
  not (_23949_, _23511_);
  and (_23950_, _23327_, _23313_);
  and (_23951_, _23950_, _23949_);
  nor (_23952_, _23951_, _23048_);
  nor (_23953_, _23952_, _23948_);
  and (_23954_, _23953_, _23636_);
  not (_23955_, _23954_);
  nor (_23957_, _23953_, _23636_);
  nor (_23958_, _23957_, _23335_);
  and (_23959_, _23958_, _23955_);
  and (_23960_, _23485_, _23048_);
  not (_23961_, _23960_);
  and (_23963_, _23479_, _23046_);
  nor (_23964_, _23963_, _23316_);
  and (_23965_, _23964_, _23961_);
  nor (_23966_, _23965_, _23959_);
  and (_23967_, _23489_, _23196_);
  and (_23968_, _23479_, _23198_);
  nor (_23969_, _23968_, _23967_);
  nor (_23970_, _23479_, _23181_);
  and (_23971_, _23492_, _23184_);
  nor (_23972_, _23490_, _23193_);
  or (_23973_, _23972_, _23971_);
  nor (_23974_, _23973_, _23970_);
  and (_23975_, _23974_, _23969_);
  and (_23976_, _23975_, _23966_);
  nor (_23977_, _23976_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23978_, _23028_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23979_, _23978_, _23025_);
  nor (_23980_, _23979_, _23977_);
  not (_23981_, _23980_);
  nor (_23982_, _23981_, _23944_);
  nor (_23983_, _23982_, _23424_);
  and (_23984_, _23983_, _23932_);
  and (_23985_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_23227_, _23985_, _23984_);
  nor (_23986_, _23701_, _23446_);
  and (_23987_, _23986_, _23705_);
  and (_23988_, _23987_, _23938_);
  and (_23989_, _23988_, _23751_);
  not (_23990_, _23988_);
  and (_23991_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_24194_, _23991_, _23989_);
  nor (_23992_, _23950_, _23949_);
  not (_23993_, _23992_);
  and (_23994_, _23993_, _23952_);
  and (_23995_, _23314_, _23330_);
  nor (_23996_, _23511_, _23995_);
  nor (_23997_, _23996_, _23946_);
  nor (_23998_, _23997_, _23046_);
  nor (_23999_, _23998_, _23994_);
  nor (_24000_, _23999_, _23335_);
  and (_24002_, _23518_, _23048_);
  and (_24003_, _23949_, _23046_);
  nor (_24004_, _24003_, _24002_);
  nor (_24005_, _24004_, _23316_);
  nor (_24006_, _24005_, _24000_);
  and (_24008_, _23521_, _23196_);
  and (_24009_, _23511_, _23198_);
  nor (_24010_, _24009_, _24008_);
  nor (_24011_, _23511_, _23181_);
  and (_24012_, _23523_, _23184_);
  nor (_24013_, _23522_, _23193_);
  or (_24014_, _24013_, _24012_);
  nor (_24015_, _24014_, _24011_);
  and (_24016_, _24015_, _24010_);
  and (_24017_, _24016_, _24006_);
  nor (_24018_, _24017_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_24019_, _23686_, _22989_);
  and (_24020_, _24019_, _23708_);
  and (_24021_, _22989_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_24022_, _24021_);
  and (_24023_, _22986_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_24024_, _24023_, _24022_);
  or (_24025_, _24024_, _24020_);
  nor (_24026_, _24025_, _24018_);
  nor (_24027_, _24026_, _23424_);
  and (_24028_, _24027_, _23932_);
  and (_24029_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_24794_, _24029_, _24028_);
  and (_24030_, _23939_, _23751_);
  and (_24031_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or (_25009_, _24031_, _24030_);
  nand (_24032_, _23455_, _23015_);
  nor (_24033_, _24032_, _23681_);
  nor (_24034_, _23571_, _23406_);
  nor (_24035_, _24034_, _23192_);
  or (_24036_, _24035_, _23572_);
  and (_24037_, _23571_, _23196_);
  and (_24038_, _23198_, _23109_);
  nor (_24039_, _24038_, _24037_);
  and (_24040_, _23554_, _22938_);
  and (_24041_, _23067_, _23109_);
  nor (_24042_, _24041_, _24040_);
  nor (_24043_, _23181_, _23109_);
  not (_24044_, _24043_);
  and (_24045_, _24044_, _24042_);
  and (_24046_, _24045_, _24039_);
  and (_24047_, _24046_, _24036_);
  nor (_24048_, _24047_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_24049_, _23016_, _22910_);
  and (_24050_, _24049_, _23014_);
  or (_24051_, _24050_, _24048_);
  or (_24052_, _24051_, _24033_);
  and (_24053_, _24052_, _23423_);
  and (_24054_, _24053_, _23939_);
  and (_24055_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or (_27025_, _24055_, _24054_);
  or (_24056_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_24057_, _24056_, _22773_);
  nand (_24058_, _24017_, _22930_);
  and (_26173_, _24058_, _24057_);
  and (_24059_, _23939_, _23920_);
  and (_24060_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or (_26760_, _24060_, _24059_);
  and (_24061_, _23697_, _23443_);
  and (_24062_, _24061_, _23453_);
  and (_24063_, _24062_, _24027_);
  not (_24064_, _24062_);
  and (_24065_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_26791_, _24065_, _24063_);
  and (_24066_, _23939_, _23900_);
  and (_24067_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or (_00032_, _24067_, _24066_);
  and (_24068_, _23929_, _23699_);
  and (_24069_, _24068_, _23453_);
  and (_24071_, _24069_, _24053_);
  not (_24072_, _24069_);
  and (_24074_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or (_27194_, _24074_, _24071_);
  and (_24076_, _24062_, _23751_);
  and (_24077_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_00364_, _24077_, _24076_);
  or (_24078_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_24079_, _24078_, _22773_);
  or (_24080_, _23413_, _22931_);
  and (_00565_, _24080_, _24079_);
  and (_24081_, _24062_, _23715_);
  and (_24082_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_00705_, _24082_, _24081_);
  and (_24083_, _23423_, _22856_);
  and (_24084_, _24083_, _23449_);
  and (_24085_, _24084_, _23924_);
  not (_24086_, _24085_);
  and (_24087_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_24088_, _24085_, _23920_);
  or (_00968_, _24088_, _24087_);
  and (_24089_, _24062_, _23693_);
  and (_24090_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_01039_, _24090_, _24089_);
  and (_24091_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_24092_, _24085_, _23900_);
  or (_27024_, _24092_, _24091_);
  and (_24093_, _23932_, _23751_);
  and (_24094_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_27209_, _24094_, _24093_);
  and (_24095_, _24053_, _23932_);
  and (_24096_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_01416_, _24096_, _24095_);
  and (_24097_, _23699_, _23432_);
  and (_24098_, _24097_, _23719_);
  and (_24099_, _24098_, _23751_);
  not (_24100_, _24098_);
  and (_24101_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or (_01561_, _24101_, _24099_);
  and (_24102_, _23932_, _23715_);
  and (_24103_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_01677_, _24103_, _24102_);
  and (_24104_, _23932_, _23693_);
  and (_24105_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_01782_, _24105_, _24104_);
  and (_24106_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_24107_, _24085_, _23983_);
  or (_01850_, _24107_, _24106_);
  and (_24108_, _23888_, _23443_);
  and (_24109_, _24108_, _23987_);
  and (_24110_, _24109_, _23715_);
  not (_24111_, _24109_);
  and (_24112_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_27271_, _24112_, _24110_);
  and (_24113_, _24109_, _23693_);
  and (_24114_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or (_02078_, _24114_, _24113_);
  and (_24115_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_24116_, _24085_, _24027_);
  or (_02107_, _24116_, _24115_);
  and (_24117_, _24061_, _23987_);
  and (_24118_, _24117_, _24053_);
  not (_24119_, _24117_);
  and (_24120_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_02490_, _24120_, _24118_);
  and (_24121_, _24098_, _23900_);
  and (_24122_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or (_02511_, _24122_, _24121_);
  and (_24123_, _23929_, _23889_);
  and (_24124_, _23906_, _23705_);
  and (_24126_, _24124_, _24123_);
  and (_24127_, _24126_, _23983_);
  not (_24128_, _24126_);
  and (_24129_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_02537_, _24129_, _24127_);
  and (_24130_, _23705_, _23449_);
  and (_24131_, _24130_, _24097_);
  and (_24132_, _24131_, _23693_);
  not (_24133_, _24131_);
  and (_24134_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_02563_, _24134_, _24132_);
  and (_24135_, _24131_, _23983_);
  and (_24136_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_02600_, _24136_, _24135_);
  and (_24137_, _24130_, _23890_);
  and (_24138_, _24137_, _24053_);
  not (_24139_, _24137_);
  and (_24140_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_02665_, _24140_, _24138_);
  and (_24141_, _24137_, _23693_);
  and (_24142_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_02706_, _24142_, _24141_);
  and (_24143_, _24109_, _23983_);
  and (_24144_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or (_02787_, _24144_, _24143_);
  and (_24145_, _23929_, _23904_);
  and (_24146_, _24145_, _24084_);
  not (_24147_, _24146_);
  and (_24148_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and (_24149_, _24146_, _23983_);
  or (_02819_, _24149_, _24148_);
  and (_24150_, _24109_, _24027_);
  and (_24151_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or (_02837_, _24151_, _24150_);
  and (_24152_, _24109_, _23920_);
  and (_24153_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_27272_, _24153_, _24152_);
  or (_24154_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_24155_, _24154_, _22773_);
  nand (_24156_, _23976_, _22930_);
  and (_03200_, _24156_, _24155_);
  and (_24157_, _23889_, _23432_);
  and (_24158_, _24157_, _23987_);
  and (_24159_, _24158_, _23920_);
  not (_24160_, _24158_);
  and (_24161_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_27270_, _24161_, _24159_);
  and (_03412_, t1_i, _22773_);
  and (_24162_, _24158_, _23900_);
  and (_24163_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_27269_, _24163_, _24162_);
  and (_24164_, _24108_, _23909_);
  and (_24165_, _24164_, _24027_);
  not (_24166_, _24164_);
  and (_24167_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_03581_, _24167_, _24165_);
  and (_24168_, _24158_, _23715_);
  and (_24169_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_27268_, _24169_, _24168_);
  and (_24170_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_24171_, _24085_, _23693_);
  or (_27023_, _24171_, _24170_);
  and (_24172_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_24173_, _24085_, _23751_);
  or (_03910_, _24173_, _24172_);
  and (_24174_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_24175_, _24085_, _24053_);
  or (_03965_, _24175_, _24174_);
  and (_24176_, _24109_, _24053_);
  and (_24177_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_03991_, _24177_, _24176_);
  and (_24178_, _24158_, _23983_);
  and (_24179_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_04257_, _24179_, _24178_);
  and (_24180_, _24158_, _24027_);
  and (_24181_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_04331_, _24181_, _24180_);
  not (_24182_, _22881_);
  and (_24183_, _24182_, _22869_);
  and (_24184_, _24183_, _22894_);
  and (_24185_, _24184_, _22918_);
  and (_24186_, _24185_, _22857_);
  not (_24188_, _24186_);
  and (_24189_, _22881_, _22869_);
  and (_24190_, _24189_, _23207_);
  and (_24191_, _24190_, _22918_);
  and (_24192_, _24191_, _22857_);
  and (_24193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_24195_, _24193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_24196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_24197_, _24196_, _22773_);
  and (_24198_, _24197_, _24195_);
  not (_24199_, _24193_);
  and (_24200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_24201_, _24200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_24202_, _24201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_24203_, _24202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_24204_, _24203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_24205_, _24204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_24206_, _24205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_24207_, _24206_, _24199_);
  nand (_24209_, _24207_, _24198_);
  nor (_24210_, _24209_, _24192_);
  and (_04785_, _24210_, _24188_);
  and (_24211_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and (_24212_, _24146_, _23693_);
  or (_27022_, _24212_, _24211_);
  and (_24213_, _24137_, _23983_);
  and (_24214_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_04829_, _24214_, _24213_);
  and (_24215_, _23987_, _23444_);
  and (_24216_, _24215_, _23751_);
  not (_24217_, _24215_);
  and (_24218_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_27278_, _24218_, _24216_);
  and (_24219_, _24157_, _24124_);
  and (_24220_, _24219_, _23715_);
  not (_24221_, _24219_);
  and (_24222_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or (_04897_, _24222_, _24220_);
  and (_24223_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and (_24224_, _24146_, _23751_);
  or (_04951_, _24224_, _24223_);
  and (_24225_, _24137_, _23715_);
  and (_24226_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_26886_, _24226_, _24225_);
  and (_24227_, _24137_, _23920_);
  and (_24228_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_05034_, _24228_, _24227_);
  and (_24229_, _24158_, _23693_);
  and (_24230_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_05231_, _24230_, _24229_);
  and (_24231_, _24130_, _24068_);
  and (_24232_, _24231_, _23983_);
  not (_24233_, _24231_);
  and (_24234_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or (_05277_, _24234_, _24232_);
  and (_24235_, _23889_, _23697_);
  and (_24236_, _23907_, _23423_);
  and (_24237_, _23986_, _24236_);
  and (_24238_, _24237_, _24235_);
  and (_24239_, _24238_, _23693_);
  not (_24240_, _24238_);
  and (_24241_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or (_05315_, _24241_, _24239_);
  and (_24242_, _24235_, _24130_);
  and (_24243_, _24242_, _23900_);
  not (_24244_, _24242_);
  and (_24245_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or (_05397_, _24245_, _24243_);
  and (_24246_, _24242_, _23751_);
  and (_24247_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or (_05451_, _24247_, _24246_);
  and (_24248_, _24242_, _23693_);
  and (_24249_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or (_05580_, _24249_, _24248_);
  and (_24250_, _23987_, _23930_);
  and (_24251_, _24250_, _23900_);
  not (_24252_, _24250_);
  and (_24253_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_27277_, _24253_, _24251_);
  and (_24254_, _24250_, _23715_);
  and (_24255_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_27276_, _24255_, _24254_);
  and (_24257_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and (_24258_, _24146_, _23920_);
  or (_06151_, _24258_, _24257_);
  and (_24259_, _24250_, _23693_);
  and (_24261_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_27275_, _24261_, _24259_);
  and (_24262_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and (_24263_, _24146_, _23900_);
  or (_06564_, _24263_, _24262_);
  and (_24264_, _24250_, _23983_);
  and (_24265_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_06887_, _24265_, _24264_);
  and (_24266_, _24250_, _24027_);
  and (_24267_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_06914_, _24267_, _24266_);
  and (_24268_, _24237_, _23700_);
  and (_24269_, _24268_, _23751_);
  not (_24270_, _24268_);
  and (_24271_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or (_06973_, _24271_, _24269_);
  and (_24272_, _24250_, _23920_);
  and (_24273_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_07186_, _24273_, _24272_);
  and (_24274_, _23904_, _23697_);
  and (_24275_, _24274_, _24084_);
  not (_24276_, _24275_);
  and (_24277_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and (_24278_, _24275_, _24027_);
  or (_07594_, _24278_, _24277_);
  and (_24279_, _24117_, _23715_);
  and (_24280_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_07678_, _24280_, _24279_);
  and (_24281_, _24117_, _23920_);
  and (_24282_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_07738_, _24282_, _24281_);
  nand (_24283_, _23976_, _23252_);
  nor (_24284_, _23256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor (_24285_, _24284_, _23257_);
  nor (_24286_, _24285_, _23210_);
  not (_24287_, _24286_);
  and (_24288_, _24287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_24289_, _23274_, _23268_);
  or (_24290_, _24289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_24292_, _24285_, _23276_);
  and (_24293_, _24292_, _24290_);
  and (_24294_, _24284_, _23276_);
  and (_24295_, _24294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_24296_, _24295_, _24293_);
  nor (_24297_, _24296_, _23210_);
  or (_24298_, _24297_, _24288_);
  or (_24299_, _24298_, _23252_);
  and (_24300_, _24299_, _22773_);
  and (_07761_, _24300_, _24283_);
  and (_24301_, _24117_, _23900_);
  and (_24302_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_27273_, _24302_, _24301_);
  and (_07889_, t0_i, _22773_);
  and (_24303_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and (_24304_, _24275_, _23920_);
  or (_27020_, _24304_, _24303_);
  and (_24305_, _24237_, _24068_);
  and (_24307_, _24305_, _24053_);
  not (_24308_, _24305_);
  and (_24309_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_27046_, _24309_, _24307_);
  and (_24310_, _24117_, _23983_);
  and (_24312_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_27274_, _24312_, _24310_);
  and (_24313_, _23892_, _23715_);
  and (_24314_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or (_27223_, _24314_, _24313_);
  and (_24315_, _24250_, _24053_);
  and (_24316_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_08689_, _24316_, _24315_);
  and (_24317_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and (_24318_, _24146_, _24053_);
  or (_08895_, _24318_, _24317_);
  and (_24319_, _24097_, _23453_);
  and (_24320_, _24319_, _23900_);
  not (_24321_, _24319_);
  and (_24322_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_09009_, _24322_, _24320_);
  and (_24323_, _23708_, _23250_);
  nor (_24324_, _23249_, _23207_);
  and (_24325_, _24324_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_24326_, _24325_, _24323_);
  and (_24328_, _22838_, _23439_);
  nor (_24329_, _22809_, _22908_);
  and (_24330_, _22914_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_24331_, _24330_, _22855_);
  and (_24332_, _24331_, _24329_);
  and (_24333_, _24332_, _24328_);
  and (_24335_, _24333_, _24326_);
  not (_24336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_24337_, _24333_, _22894_);
  nor (_24338_, _24337_, _24336_);
  nor (_24339_, _22822_, _22809_);
  and (_24340_, _24339_, _22856_);
  and (_24341_, _23249_, _23207_);
  and (_24342_, _22915_, _22908_);
  and (_24343_, _24342_, _24341_);
  and (_24344_, _24343_, _24340_);
  or (_24345_, _24344_, _24338_);
  or (_24346_, _24345_, _24335_);
  not (_24347_, _24344_);
  or (_24348_, _24347_, _23413_);
  and (_24349_, _24348_, _22773_);
  and (_09255_, _24349_, _24346_);
  and (_24350_, _24333_, _24184_);
  or (_24351_, _24350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24352_, _24351_, _24347_);
  nand (_24353_, _24350_, _23681_);
  and (_24354_, _24353_, _24352_);
  and (_24355_, _24344_, _23247_);
  or (_24356_, _24355_, _24354_);
  and (_09302_, _24356_, _22773_);
  and (_24357_, _24333_, _22895_);
  or (_24358_, _24357_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24359_, _24358_, _24347_);
  nand (_24360_, _24357_, _23681_);
  and (_24361_, _24360_, _24359_);
  and (_24362_, _24344_, _23744_);
  or (_24363_, _24362_, _24361_);
  and (_09331_, _24363_, _22773_);
  nand (_24364_, _24337_, _24189_);
  nor (_24365_, _24364_, _23681_);
  and (_24366_, _24364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_24367_, _24366_, _24344_);
  or (_24368_, _24367_, _24365_);
  nand (_24369_, _24344_, _24047_);
  and (_24370_, _24369_, _22773_);
  and (_09351_, _24370_, _24368_);
  and (_24371_, _24117_, _23751_);
  and (_24372_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_09433_, _24372_, _24371_);
  and (_24373_, _24183_, _23207_);
  and (_24374_, _24373_, _24333_);
  nand (_24375_, _24374_, _23681_);
  or (_24376_, _24374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_24377_, _24376_, _24347_);
  and (_24378_, _24377_, _24375_);
  nor (_24379_, _24347_, _24017_);
  or (_24380_, _24379_, _24378_);
  and (_09536_, _24380_, _22773_);
  and (_24381_, _24333_, _23208_);
  nand (_24382_, _24381_, _23681_);
  or (_24383_, _24381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24384_, _24383_, _24347_);
  and (_24385_, _24384_, _24382_);
  nor (_24386_, _24347_, _23357_);
  or (_24387_, _24386_, _24385_);
  and (_09573_, _24387_, _22773_);
  and (_24388_, _23906_, _23452_);
  and (_24389_, _24388_, _23924_);
  and (_24390_, _24389_, _23920_);
  not (_24391_, _24389_);
  and (_24392_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_27189_, _24392_, _24390_);
  and (_24393_, _24084_, _24061_);
  not (_24394_, _24393_);
  and (_24395_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and (_24396_, _24393_, _24027_);
  or (_09661_, _24396_, _24395_);
  and (_24397_, _24235_, _23987_);
  and (_24398_, _24397_, _23983_);
  not (_24399_, _24397_);
  and (_24400_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_27261_, _24400_, _24398_);
  and (_24401_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and (_24402_, _24393_, _23920_);
  or (_27007_, _24402_, _24401_);
  and (_24403_, _23439_, _22809_);
  and (_24404_, _24403_, _22856_);
  and (_24405_, _24189_, _22894_);
  and (_24406_, _24405_, _22918_);
  and (_24407_, _24406_, _24404_);
  and (_24408_, _22809_, _22926_);
  and (_24410_, _24331_, _24328_);
  and (_24411_, _24410_, _24408_);
  and (_24412_, _24411_, _22895_);
  nand (_24413_, _24412_, _23681_);
  or (_24414_, _24412_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24415_, _24414_, _24413_);
  or (_24416_, _24415_, _24407_);
  not (_24417_, _24407_);
  or (_24418_, _24417_, _23744_);
  and (_24419_, _24418_, _22773_);
  and (_09763_, _24419_, _24416_);
  not (_24420_, _24330_);
  nor (_24421_, _24420_, _22908_);
  and (_24422_, _22855_, _22809_);
  and (_24423_, _24422_, _24421_);
  nand (_24424_, _24423_, _24328_);
  nor (_24425_, _24189_, _22894_);
  or (_24426_, _24425_, _24405_);
  or (_24427_, _24426_, _24424_);
  and (_24428_, _24427_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_24429_, _24428_, _24407_);
  and (_24431_, _24190_, _23708_);
  nor (_24432_, _24189_, _23207_);
  and (_24433_, _24432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_24434_, _24433_, _24431_);
  and (_24435_, _24434_, _24411_);
  or (_24436_, _24435_, _24429_);
  or (_24437_, _24417_, _23205_);
  and (_24438_, _24437_, _22773_);
  and (_09790_, _24438_, _24436_);
  and (_24439_, _24397_, _24027_);
  and (_24440_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or (_09808_, _24440_, _24439_);
  or (_24441_, _24424_, _23207_);
  and (_24442_, _24441_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_24443_, _24442_, _24407_);
  and (_24444_, _24324_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_24445_, _24444_, _24323_);
  and (_24446_, _24445_, _24411_);
  or (_24447_, _24446_, _24443_);
  or (_24448_, _24417_, _23413_);
  and (_24449_, _24448_, _22773_);
  and (_09826_, _24449_, _24447_);
  and (_24450_, _24411_, _24184_);
  nand (_24451_, _24450_, _23681_);
  or (_24452_, _24450_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24453_, _24452_, _24451_);
  or (_24454_, _24453_, _24407_);
  or (_24455_, _24417_, _23247_);
  and (_24456_, _24455_, _22773_);
  and (_09861_, _24456_, _24454_);
  and (_24457_, _24411_, _24405_);
  nand (_24458_, _24457_, _23681_);
  or (_24459_, _24457_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24460_, _24459_, _24458_);
  or (_24461_, _24460_, _24407_);
  nand (_24462_, _24407_, _24047_);
  and (_24463_, _24462_, _22773_);
  and (_09879_, _24463_, _24461_);
  and (_24464_, _24268_, _24053_);
  and (_24466_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or (_27044_, _24466_, _24464_);
  or (_24467_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_24468_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_24469_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_24470_, _24469_, _24468_);
  and (_24471_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not (_24472_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_24473_, _24472_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_24474_, _24473_, _24468_);
  and (_24475_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_24476_, _24475_, _24471_);
  and (_24477_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_24478_, _24477_, _24468_);
  and (_24479_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_24480_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_24481_, _24480_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_24482_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_24483_, _24482_, _24479_);
  and (_24484_, _24469_, _24468_);
  and (_24485_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_24486_, _24469_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_24487_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_24488_, _24487_, _24485_);
  and (_24489_, _24488_, _24483_);
  and (_24490_, _24489_, _24476_);
  nor (_24492_, _24490_, _24467_);
  and (_24494_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_24495_, _24494_, _24492_);
  and (_24497_, _24495_, _23761_);
  not (_24498_, _24497_);
  not (_24500_, _23758_);
  nor (_24501_, _23760_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_24502_, _24501_, _24500_);
  and (_24503_, _24502_, _24498_);
  and (_24504_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_24505_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_24506_, _24505_, _24504_);
  nand (_24507_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand (_24508_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_24509_, _24508_, _24507_);
  nand (_24510_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_24511_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_24512_, _24511_, _24510_);
  and (_24513_, _24512_, _24509_);
  and (_24514_, _24513_, _24506_);
  or (_24515_, _24514_, _24467_);
  and (_24516_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not (_24517_, _24516_);
  and (_24518_, _24517_, _24515_);
  nand (_24519_, _24518_, _23761_);
  nor (_24520_, _23760_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_24521_, _24520_, _24500_);
  and (_24522_, _24521_, _24519_);
  and (_24523_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_24524_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_24525_, _24524_, _24523_);
  nand (_24526_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nand (_24527_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_24528_, _24527_, _24526_);
  nand (_24529_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_24530_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_24531_, _24530_, _24529_);
  and (_24532_, _24531_, _24528_);
  and (_24533_, _24532_, _24525_);
  or (_24534_, _24533_, _24467_);
  and (_24535_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24536_, _24535_);
  and (_24537_, _24536_, _24534_);
  nand (_24538_, _24537_, _23761_);
  nor (_24539_, _23760_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_24540_, _24539_, _24500_);
  and (_24541_, _24540_, _24538_);
  nor (_24542_, _24541_, _24522_);
  and (_24543_, _24542_, _24503_);
  and (_24544_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_24545_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_24546_, _24545_, _24544_);
  nand (_24548_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_24549_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_24550_, _24549_, _24548_);
  nand (_24551_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand (_24553_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_24554_, _24553_, _24551_);
  and (_24555_, _24554_, _24550_);
  and (_24556_, _24555_, _24546_);
  or (_24557_, _24467_, _24556_);
  and (_24559_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  not (_24560_, _24559_);
  and (_24561_, _24560_, _24557_);
  nand (_24562_, _24561_, _23761_);
  nor (_24563_, _23760_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_24564_, _24563_, _24500_);
  and (_24565_, _24564_, _24562_);
  not (_24566_, _24565_);
  not (_24567_, _23761_);
  not (_24568_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24569_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_24570_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_24571_, _24570_, _24569_);
  and (_24572_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_24573_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_24574_, _24573_, _24572_);
  and (_24575_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_24576_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_24577_, _24576_, _24575_);
  or (_24578_, _24577_, _24574_);
  or (_24579_, _24578_, _24571_);
  and (_24580_, _24579_, _24568_);
  or (_24581_, _24580_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24582_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_24583_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _24582_);
  not (_24585_, _24583_);
  and (_24586_, _24585_, _24581_);
  or (_24588_, _24586_, _24567_);
  nor (_24589_, _23760_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_24590_, _24589_, _24500_);
  and (_24591_, _24590_, _24588_);
  and (_24592_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_24594_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_24595_, _24594_, _24592_);
  nand (_24596_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_24597_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_24598_, _24597_, _24596_);
  nand (_24599_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand (_24601_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_24602_, _24601_, _24599_);
  and (_24603_, _24602_, _24598_);
  nand (_24604_, _24603_, _24595_);
  nand (_24605_, _24604_, _24568_);
  nand (_24606_, _24605_, _24582_);
  nor (_24608_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _24582_);
  not (_24609_, _24608_);
  and (_24610_, _24609_, _24606_);
  or (_24611_, _24610_, _24567_);
  nor (_24612_, _23760_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_24613_, _24612_, _24500_);
  and (_24615_, _24613_, _24611_);
  nor (_24616_, _24615_, _24591_);
  and (_24617_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_24618_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_24619_, _24618_, _24617_);
  and (_24620_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not (_24621_, _24620_);
  and (_24622_, _24621_, _24619_);
  nand (_24623_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_24624_, _24623_, _24568_);
  and (_24625_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_24626_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_24627_, _24626_, _24625_);
  and (_24628_, _24627_, _24624_);
  and (_24629_, _24628_, _24622_);
  and (_24630_, _24629_, _24582_);
  nor (_24631_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _24582_);
  or (_24632_, _24631_, _24630_);
  and (_24633_, _24632_, _23761_);
  not (_24634_, _24633_);
  nor (_24635_, _23760_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_24636_, _24635_, _24500_);
  and (_24637_, _24636_, _24634_);
  and (_24638_, _24637_, _24616_);
  and (_24639_, _24638_, _24566_);
  and (_24640_, _24639_, _24543_);
  and (_24641_, \oc8051_top_1.oc8051_decoder1.state [1], _22781_);
  and (_24642_, _24641_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_24643_, _24642_, _24640_);
  not (_24644_, _24643_);
  or (_24646_, _23759_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_24647_, _24646_);
  and (_24648_, _24638_, _24565_);
  and (_24649_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_24650_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_24651_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_24652_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_24653_, _24652_, _24651_);
  and (_24654_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_24655_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_24657_, _24655_, _24654_);
  nand (_24658_, _24657_, _24653_);
  or (_24659_, _24658_, _24650_);
  nor (_24660_, _24659_, _24649_);
  and (_24661_, _24660_, _24568_);
  and (_24662_, _24661_, _24582_);
  nor (_24663_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _24582_);
  nor (_24664_, _24663_, _24662_);
  nor (_24665_, _24664_, _24567_);
  not (_24666_, _24665_);
  nor (_24667_, _23760_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_24668_, _24667_, _24500_);
  and (_24669_, _24668_, _24666_);
  not (_24670_, _24669_);
  not (_24671_, _24541_);
  and (_24672_, _24671_, _24522_);
  and (_24673_, _24672_, _24503_);
  and (_24674_, _24673_, _24670_);
  and (_24675_, _24674_, _24648_);
  not (_24676_, _24503_);
  and (_24677_, _24672_, _24676_);
  and (_24678_, _24677_, _24669_);
  not (_24679_, _24522_);
  and (_24680_, _24541_, _24679_);
  and (_24681_, _24680_, _24503_);
  and (_24682_, _24681_, _24669_);
  or (_24683_, _24682_, _24678_);
  and (_24684_, _24683_, _24648_);
  nor (_24685_, _24684_, _24675_);
  and (_24686_, _24541_, _24522_);
  and (_24687_, _24686_, _24676_);
  not (_24688_, _24615_);
  and (_24689_, _24637_, _24591_);
  and (_24690_, _24689_, _24688_);
  and (_24691_, _24690_, _24687_);
  and (_24693_, _24690_, _24678_);
  or (_24694_, _24693_, _24691_);
  and (_24696_, _24686_, _24503_);
  and (_24697_, _24696_, _24670_);
  and (_24698_, _24680_, _24676_);
  and (_24699_, _24698_, _24670_);
  or (_24700_, _24699_, _24697_);
  and (_24702_, _24700_, _24690_);
  not (_24703_, _24690_);
  and (_24704_, _24698_, _24669_);
  nor (_24705_, _24704_, _24543_);
  nor (_24706_, _24705_, _24703_);
  or (_24707_, _24706_, _24702_);
  nor (_24708_, _24707_, _24694_);
  and (_24709_, _24677_, _24670_);
  and (_24710_, _24709_, _24690_);
  not (_24711_, _24710_);
  and (_24712_, _24673_, _24669_);
  and (_24714_, _24712_, _24690_);
  and (_24715_, _24681_, _24670_);
  and (_24716_, _24715_, _24690_);
  nor (_24717_, _24716_, _24714_);
  and (_24718_, _24717_, _24711_);
  not (_24719_, _24640_);
  nor (_24720_, _24637_, _24565_);
  and (_24721_, _24720_, _24616_);
  and (_24722_, _24687_, _24669_);
  and (_24723_, _24722_, _24721_);
  and (_24724_, _24542_, _24676_);
  and (_24725_, _24724_, _24690_);
  nor (_24726_, _24725_, _24723_);
  and (_24727_, _24726_, _24719_);
  and (_24728_, _24727_, _24718_);
  and (_24729_, _24728_, _24708_);
  and (_24730_, _24729_, _24685_);
  nor (_24731_, _24730_, _24647_);
  not (_24732_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_24733_, _24641_, _24732_);
  and (_24735_, _24733_, _24681_);
  and (_24736_, _24735_, _24721_);
  nor (_24737_, _24736_, _24731_);
  and (_24738_, _24737_, _24644_);
  nor (_26832_[0], _24738_, rst);
  and (_24740_, _24235_, _23706_);
  and (_24741_, _24740_, _23983_);
  not (_24742_, _24740_);
  and (_24743_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_10156_, _24743_, _24741_);
  and (_24745_, _24411_, _24373_);
  or (_24746_, _24745_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_24747_, _24746_, _24417_);
  nand (_24748_, _24745_, _23681_);
  and (_24749_, _24748_, _24747_);
  nor (_24750_, _24417_, _24017_);
  or (_24751_, _24750_, _24749_);
  and (_10212_, _24751_, _22773_);
  and (_24752_, _24123_, _23987_);
  and (_24753_, _24752_, _23693_);
  not (_24754_, _24752_);
  and (_24755_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_10313_, _24755_, _24753_);
  and (_24756_, _24752_, _23751_);
  and (_24757_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_10419_, _24757_, _24756_);
  and (_24758_, _22838_, _22822_);
  and (_24759_, _24758_, _24423_);
  and (_24761_, _24759_, _24190_);
  or (_24762_, _24761_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_24763_, _24406_, _22857_);
  not (_24764_, _24763_);
  and (_24765_, _24764_, _24762_);
  nand (_24767_, _24761_, _23681_);
  and (_24768_, _24767_, _24765_);
  and (_24769_, _24763_, _23205_);
  or (_24770_, _24769_, _24768_);
  and (_10435_, _24770_, _22773_);
  and (_24772_, _24759_, _24184_);
  or (_24773_, _24772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_24774_, _24773_, _24764_);
  nand (_24775_, _24772_, _23681_);
  and (_24777_, _24775_, _24774_);
  and (_24778_, _24763_, _23247_);
  or (_24779_, _24778_, _24777_);
  and (_10451_, _24779_, _22773_);
  and (_24781_, _24759_, _24405_);
  or (_24782_, _24781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_24784_, _24782_, _24764_);
  nand (_24785_, _24781_, _23681_);
  and (_24787_, _24785_, _24784_);
  not (_24788_, _24047_);
  and (_24789_, _24763_, _24788_);
  or (_24790_, _24789_, _24787_);
  and (_10467_, _24790_, _22773_);
  and (_24791_, _24752_, _24053_);
  and (_24793_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or (_10506_, _24793_, _24791_);
  and (_24795_, _24084_, _23930_);
  not (_24796_, _24795_);
  and (_24797_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and (_24798_, _24795_, _23751_);
  or (_10593_, _24798_, _24797_);
  and (_24799_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_24801_, _24795_, _24053_);
  or (_27011_, _24801_, _24799_);
  nor (_26831_[7], _24518_, rst);
  and (_24802_, _24397_, _23751_);
  and (_24803_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_27259_, _24803_, _24802_);
  nor (_24804_, _23760_, _23464_);
  and (_24805_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_24806_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_24807_, _24806_, _24805_);
  and (_24808_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_24809_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_24810_, _24809_, _24808_);
  and (_24811_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_24812_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_24813_, _24812_, _24811_);
  and (_24814_, _24813_, _24810_);
  and (_24815_, _24814_, _24807_);
  and (_24816_, _23760_, _24568_);
  not (_24817_, _24816_);
  nor (_24818_, _24817_, _24815_);
  nor (_24819_, _24818_, _24804_);
  nor (_26858_[7], _24819_, rst);
  and (_24820_, _24397_, _24053_);
  and (_24821_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_10826_, _24821_, _24820_);
  not (_24822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_24823_, _24822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not (_24824_, _24823_);
  not (_24825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_24826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_24827_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_24828_, _24827_, _24826_);
  and (_24829_, _24828_, _24825_);
  not (_24830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_24831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_24832_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_24833_, _24832_, _24831_);
  and (_24834_, _24833_, _24830_);
  nor (_24835_, _24834_, _24829_);
  and (_24836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_24837_, _24836_, _24336_);
  not (_24838_, _24837_);
  and (_24839_, _24838_, _24835_);
  nor (_24840_, _24839_, _24824_);
  not (_24841_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_24842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24843_, _24842_, _24841_);
  not (_24844_, _24843_);
  not (_24845_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24847_, _24846_, _24845_);
  not (_24848_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24850_, _24849_, _24848_);
  nor (_24851_, _24850_, _24847_);
  and (_24852_, _24851_, _24844_);
  nor (_24853_, _24852_, _24824_);
  nor (_24854_, _24853_, _24840_);
  and (_24855_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  or (_24856_, _24855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24857_, _24856_, _24854_);
  and (_24858_, _24857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  not (_24859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_24860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_24861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _24859_);
  nor (_24862_, _24861_, _24860_);
  and (_24863_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_24864_, _24863_, _24822_);
  and (_24865_, _24842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_24866_, _24865_);
  and (_24867_, _24846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24868_, _24849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_24869_, _24868_, _24867_);
  and (_24870_, _24869_, _24866_);
  nand (_24871_, _24828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_24872_, _24833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_24873_, _24872_);
  and (_24874_, _24873_, _24871_);
  and (_24875_, _24836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_24876_, _24875_);
  and (_24877_, _24876_, _24874_);
  and (_24878_, _24877_, _24870_);
  or (_24879_, _24878_, _24864_);
  nor (_24880_, _24879_, _24855_);
  and (_24881_, _24880_, _24859_);
  or (_24882_, _24881_, _24858_);
  and (_10854_, _24882_, _22773_);
  not (_24883_, _23760_);
  and (_24884_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_24885_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24886_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_24887_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_24888_, _24887_, _24886_);
  and (_24889_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_24890_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_24891_, _24890_, _24889_);
  and (_24892_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_24893_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_24894_, _24893_, _24892_);
  and (_24895_, _24894_, _24891_);
  and (_24896_, _24895_, _24888_);
  nor (_24897_, _24896_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_24898_, _24897_, _24885_);
  nor (_24899_, _24898_, _24883_);
  nor (_24900_, _24899_, _24884_);
  nor (_26868_[7], _24900_, rst);
  and (_24901_, _24237_, _23938_);
  and (_24902_, _24901_, _23983_);
  not (_24903_, _24901_);
  and (_24904_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_10924_, _24904_, _24902_);
  and (_24905_, _24397_, _23900_);
  and (_24906_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or (_11227_, _24906_, _24905_);
  and (_24907_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and (_24908_, _24393_, _24053_);
  or (_11248_, _24908_, _24907_);
  and (_24909_, _24397_, _23715_);
  and (_24910_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_11269_, _24910_, _24909_);
  or (_24911_, _24855_, _24859_);
  or (_24912_, _24911_, _24854_);
  and (_24913_, _24912_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_24914_, _24880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24915_, _24914_, _24913_);
  and (_11290_, _24915_, _22773_);
  and (_24916_, _24397_, _23693_);
  and (_24917_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or (_27260_, _24917_, _24916_);
  not (_24918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_24919_, _24879_, _24854_);
  nor (_24920_, _24919_, _24855_);
  nor (_24921_, _24920_, _24918_);
  not (_24922_, _24855_);
  nor (_24923_, _24871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24924_, _24923_, _24875_);
  and (_24925_, _24872_, _24859_);
  or (_24926_, _24925_, _24918_);
  nand (_24927_, _24926_, _24924_);
  and (_24928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_24929_, _24928_);
  nand (_24930_, _24929_, _24875_);
  and (_24931_, _24930_, _24927_);
  or (_24932_, _24931_, _24868_);
  not (_24933_, _24867_);
  not (_24934_, _24868_);
  or (_24935_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _24859_);
  or (_24936_, _24935_, _24934_);
  and (_24937_, _24936_, _24933_);
  and (_24938_, _24937_, _24932_);
  and (_24939_, _24928_, _24867_);
  or (_24940_, _24939_, _24865_);
  or (_24941_, _24940_, _24938_);
  nor (_24942_, _24935_, _24866_);
  nor (_24943_, _24942_, _24879_);
  and (_24944_, _24943_, _24941_);
  or (_24945_, _24935_, _24844_);
  not (_24946_, _24854_);
  and (_24947_, _24879_, _24946_);
  and (_24948_, _24829_, _24859_);
  nor (_24949_, _24948_, _24837_);
  and (_24950_, _24834_, _24859_);
  or (_24951_, _24950_, _24918_);
  nand (_24952_, _24951_, _24949_);
  nand (_24953_, _24929_, _24837_);
  and (_24954_, _24953_, _24952_);
  or (_24955_, _24954_, _24850_);
  not (_24956_, _24847_);
  not (_24957_, _24850_);
  or (_24958_, _24935_, _24957_);
  and (_24959_, _24958_, _24956_);
  and (_24960_, _24959_, _24955_);
  and (_24961_, _24928_, _24847_);
  or (_24962_, _24961_, _24843_);
  or (_24963_, _24962_, _24960_);
  and (_24964_, _24963_, _24947_);
  and (_24965_, _24964_, _24945_);
  or (_24966_, _24965_, _24944_);
  and (_24967_, _24966_, _24922_);
  or (_24968_, _24967_, _24921_);
  and (_11499_, _24968_, _22773_);
  not (_24969_, _24919_);
  or (_24970_, _24969_, _24856_);
  and (_24971_, _24879_, _24922_);
  or (_24972_, _24971_, _24859_);
  and (_24973_, _24972_, _22773_);
  and (_11627_, _24973_, _24970_);
  nand (_24974_, _24192_, _23976_);
  nor (_24975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_24976_, _24975_);
  not (_24977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_24978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_24979_, _24978_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_24980_, t0_i);
  and (_24981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _24980_);
  and (_24982_, _24981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  or (_24983_, _24982_, _24979_);
  and (_24984_, _24983_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_24985_, _24984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_24986_, _24985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_24987_, _24986_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_24988_, _24987_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_24989_, _24988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand (_24990_, _24989_, _24205_);
  and (_24991_, _24990_, _24977_);
  or (_24992_, _24991_, _24976_);
  and (_24993_, _24989_, _24206_);
  nor (_24994_, _24993_, _24992_);
  and (_24995_, _24205_, _24193_);
  or (_24996_, _24995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_24997_, _24206_, _24193_);
  and (_24998_, _24997_, _24196_);
  and (_24999_, _24998_, _24996_);
  not (_25000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_25001_, _25000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_25002_, _25000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_25003_, _25002_, _25001_);
  and (_25004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_25005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_25006_, _25005_, _25004_);
  and (_25007_, _25006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_25008_, _25007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_25010_, _25008_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_25011_, _25010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_25012_, _25011_, _24984_);
  and (_25013_, _24204_, _25000_);
  and (_25014_, _25013_, _25012_);
  and (_25015_, _25014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_25016_, _25015_, _24977_);
  and (_25017_, _25015_, _24977_);
  or (_25018_, _25017_, _25016_);
  and (_25019_, _25018_, _25003_);
  or (_25020_, _25019_, _24999_);
  or (_25021_, _25020_, _24994_);
  or (_25022_, _25021_, _24192_);
  and (_25023_, _25022_, _24188_);
  and (_25024_, _25023_, _24974_);
  and (_25025_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_25026_, _25025_, _25024_);
  and (_11736_, _25026_, _22773_);
  not (_25027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_25028_, _23268_, _25027_);
  and (_25029_, _25028_, _24284_);
  or (_25030_, _25029_, _23373_);
  or (_25031_, _25028_, _23281_);
  and (_25032_, _25031_, _25030_);
  or (_25033_, _25032_, _23257_);
  and (_25034_, _25030_, _23281_);
  or (_25035_, _25034_, _23360_);
  and (_25036_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_25037_, _25036_, _23361_);
  and (_25038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_25039_, _25038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_25040_, _25039_, _25037_);
  and (_25041_, _25040_, _23268_);
  and (_25042_, _25041_, _25035_);
  or (_25043_, _25042_, _25028_);
  and (_25044_, _25043_, _25033_);
  and (_25045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_25046_, _25045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_25047_, _25046_, _24294_);
  or (_25048_, _25047_, _25044_);
  nor (_25049_, _23252_, rst);
  and (_25050_, _25049_, _23211_);
  and (_11840_, _25050_, _25048_);
  not (_25051_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_25052_, _24920_, _25051_);
  or (_25053_, _24876_, _24868_);
  and (_25054_, _25053_, _24933_);
  and (_25055_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _24859_);
  or (_25056_, _25055_, _25054_);
  and (_25057_, _24872_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25058_, _25057_, _25051_);
  nor (_25059_, _24871_, _24859_);
  nor (_25060_, _25059_, _24875_);
  and (_25061_, _25060_, _24869_);
  nand (_25062_, _25061_, _25058_);
  and (_25063_, _25062_, _25056_);
  or (_25064_, _25063_, _24865_);
  or (_25065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25066_, _24934_, _24867_);
  and (_25067_, _25066_, _24866_);
  nor (_25068_, _25067_, _25065_);
  nor (_25069_, _25068_, _24879_);
  and (_25071_, _25069_, _25064_);
  and (_25072_, _24829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25074_, _25072_, _24837_);
  and (_25075_, _24834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25076_, _25075_, _25051_);
  nand (_25077_, _25076_, _25074_);
  or (_25078_, _25055_, _24838_);
  and (_25079_, _25078_, _25077_);
  or (_25080_, _25079_, _24850_);
  or (_25081_, _25065_, _24957_);
  and (_25082_, _25081_, _24956_);
  and (_25083_, _25082_, _25080_);
  and (_25084_, _25055_, _24847_);
  or (_25085_, _25084_, _24843_);
  or (_25086_, _25085_, _25083_);
  and (_25087_, _24947_, _24844_);
  and (_25088_, _25065_, _24947_);
  or (_25089_, _25088_, _25087_);
  and (_25090_, _25089_, _25086_);
  or (_25091_, _25090_, _25071_);
  and (_25092_, _25091_, _24922_);
  or (_25093_, _25092_, _25052_);
  and (_11871_, _25093_, _22773_);
  and (_25094_, _24752_, _24027_);
  and (_25095_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or (_11983_, _25095_, _25094_);
  and (_25096_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and (_25097_, _24393_, _23715_);
  or (_12004_, _25097_, _25096_);
  and (_25098_, _24752_, _23920_);
  and (_25099_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or (_27266_, _25099_, _25098_);
  and (_25100_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  and (_25101_, _24393_, _23693_);
  or (_12219_, _25101_, _25100_);
  and (_25102_, _24855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_25103_, _25102_, _24920_);
  and (_12309_, _25103_, _22773_);
  or (_25104_, _24850_, _24837_);
  nor (_25105_, _24847_, _24843_);
  nand (_25106_, _25105_, _24823_);
  or (_25107_, _25106_, _25104_);
  nor (_25108_, _25107_, _24835_);
  and (_25109_, _25108_, _24879_);
  and (_25110_, _24855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or (_25111_, _24875_, _24855_);
  nor (_25112_, _25111_, _24864_);
  not (_25113_, _24870_);
  nor (_25114_, _24874_, _25113_);
  and (_25115_, _25114_, _25112_);
  or (_25116_, _25115_, _25110_);
  or (_25117_, _25116_, _25109_);
  and (_12333_, _25117_, _22773_);
  and (_25118_, _24835_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_25119_, _25118_, _25104_);
  and (_25120_, _25119_, _25105_);
  and (_25121_, _25120_, _24947_);
  nor (_25122_, _24867_, _24865_);
  or (_25123_, _24875_, _24868_);
  and (_25124_, _24874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_25125_, _25124_, _25123_);
  and (_25126_, _25125_, _25122_);
  nor (_25127_, _25126_, _24855_);
  nor (_25128_, _25127_, _24971_);
  or (_25129_, _25128_, _25121_);
  or (_25131_, _24922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_25132_, _25131_, _22773_);
  and (_12358_, _25132_, _25129_);
  nor (_25133_, _24834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_25134_, _25133_, _24829_);
  or (_25135_, _25134_, _24837_);
  and (_25136_, _25135_, _24957_);
  or (_25137_, _25136_, _24847_);
  and (_25138_, _25137_, _25087_);
  or (_25139_, _24872_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25140_, _25139_, _24871_);
  or (_25141_, _25140_, _24875_);
  and (_25142_, _25141_, _24934_);
  or (_25143_, _25142_, _24867_);
  nor (_25144_, _24879_, _24865_);
  and (_25145_, _25144_, _25143_);
  or (_25146_, _25145_, _24855_);
  or (_25147_, _25146_, _25138_);
  or (_25148_, _24922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25149_, _25148_, _22773_);
  and (_12399_, _25149_, _25147_);
  and (_25150_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _22773_);
  and (_12420_, _25150_, _24855_);
  and (_25151_, _24158_, _24053_);
  and (_25152_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_12621_, _25152_, _25151_);
  and (_25153_, _24108_, _24084_);
  not (_25154_, _25153_);
  and (_25155_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_25156_, _25153_, _23715_);
  or (_12759_, _25156_, _25155_);
  and (_25157_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_25158_, _25153_, _23693_);
  or (_12910_, _25158_, _25157_);
  and (_25159_, _23700_, _23453_);
  and (_25160_, _25159_, _24053_);
  not (_25161_, _25159_);
  and (_25162_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or (_27191_, _25162_, _25160_);
  nand (_25163_, _23451_, _23423_);
  and (_25164_, _23986_, _25163_);
  and (_25165_, _25164_, _23905_);
  and (_25166_, _25165_, _24053_);
  not (_25167_, _25165_);
  and (_25168_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_13221_, _25168_, _25166_);
  and (_25169_, _24068_, _23719_);
  and (_25170_, _25169_, _23715_);
  not (_25171_, _25169_);
  and (_25172_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_13520_, _25172_, _25170_);
  and (_25173_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_25174_, _25153_, _24027_);
  or (_13601_, _25174_, _25173_);
  and (_25175_, _23907_, _23449_);
  and (_25176_, _25175_, _24235_);
  and (_25177_, _25176_, _24027_);
  not (_25178_, _25176_);
  and (_25179_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or (_13792_, _25179_, _25177_);
  and (_25180_, _24388_, _24157_);
  and (_25181_, _25180_, _23900_);
  not (_25182_, _25180_);
  and (_25183_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or (_13813_, _25183_, _25181_);
  and (_25184_, _25180_, _24027_);
  and (_25185_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or (_13864_, _25185_, _25184_);
  and (_25186_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_25187_, _25153_, _23920_);
  or (_13885_, _25187_, _25186_);
  and (_25188_, _25180_, _23983_);
  and (_25189_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or (_13976_, _25189_, _25188_);
  and (_25190_, _23938_, _23453_);
  and (_25191_, _25190_, _23751_);
  not (_25192_, _25190_);
  and (_25193_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_27190_, _25193_, _25191_);
  and (_25194_, _24388_, _24108_);
  and (_25195_, _25194_, _24053_);
  not (_25196_, _25194_);
  and (_25197_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_14057_, _25197_, _25195_);
  and (_25198_, _24388_, _23890_);
  and (_25199_, _25198_, _23693_);
  not (_25200_, _25198_);
  and (_25201_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or (_14118_, _25201_, _25199_);
  and (_25202_, _24389_, _24027_);
  and (_25203_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_14209_, _25203_, _25202_);
  and (_25204_, _25198_, _23715_);
  and (_25205_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or (_14469_, _25205_, _25204_);
  and (_25206_, _25198_, _23920_);
  and (_25207_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or (_14520_, _25207_, _25206_);
  and (_25208_, _25198_, _23983_);
  and (_25209_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_14591_, _25209_, _25208_);
  and (_25210_, _24388_, _24235_);
  and (_25211_, _25210_, _23751_);
  not (_25212_, _25210_);
  and (_25213_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_14652_, _25213_, _25211_);
  and (_25214_, _25210_, _23693_);
  and (_25215_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_14743_, _25215_, _25214_);
  and (_25216_, _25210_, _23900_);
  and (_25217_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_27107_, _25217_, _25216_);
  and (_25218_, _25210_, _23920_);
  and (_25219_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_27108_, _25219_, _25218_);
  and (_25220_, _24388_, _24123_);
  and (_25221_, _25220_, _23751_);
  not (_25222_, _25220_);
  and (_25223_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_14974_, _25223_, _25221_);
  and (_25224_, _22809_, _22908_);
  and (_25225_, _25224_, _22855_);
  and (_25226_, _25225_, _24758_);
  nand (_25227_, _25226_, _22894_);
  and (_25228_, _25227_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_25229_, _24324_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_25230_, _25229_, _24323_);
  and (_25231_, _25230_, _25226_);
  or (_25232_, _25231_, _25228_);
  and (_25233_, _25232_, _24330_);
  and (_25234_, _22894_, _22908_);
  and (_25235_, _25234_, _24189_);
  and (_25236_, _25235_, _22857_);
  not (_25237_, _25236_);
  or (_25238_, _25237_, _23413_);
  or (_25239_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_25240_, _25239_, _22915_);
  and (_25241_, _25240_, _25238_);
  not (_25242_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_25243_, _22914_, _25242_);
  or (_25244_, _25243_, rst);
  or (_25245_, _25244_, _25241_);
  or (_14995_, _25245_, _25233_);
  and (_25246_, _25220_, _23715_);
  and (_25247_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_15046_, _25247_, _25246_);
  and (_25248_, _25226_, _24373_);
  nand (_25249_, _25248_, _23681_);
  or (_25250_, _25248_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25251_, _25250_, _24330_);
  and (_25252_, _25251_, _25249_);
  nand (_25253_, _25236_, _24017_);
  or (_25254_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25255_, _25254_, _22915_);
  and (_25256_, _25255_, _25253_);
  not (_25257_, _22914_);
  and (_25258_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_25259_, _25258_, rst);
  or (_25260_, _25259_, _25256_);
  or (_15092_, _25260_, _25252_);
  and (_25261_, _25226_, _23208_);
  nand (_25262_, _25261_, _23681_);
  or (_25263_, _25261_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25264_, _25263_, _24330_);
  and (_25265_, _25264_, _25262_);
  nand (_25266_, _25236_, _23357_);
  or (_25267_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25268_, _25267_, _22915_);
  and (_25269_, _25268_, _25266_);
  not (_25270_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_25271_, _22914_, _25270_);
  or (_25272_, _25271_, rst);
  or (_25273_, _25272_, _25269_);
  or (_15106_, _25273_, _25265_);
  not (_25274_, _25226_);
  or (_25275_, _25274_, _24426_);
  and (_25276_, _25275_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25277_, _24432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_25278_, _25277_, _24431_);
  and (_25279_, _25278_, _25226_);
  or (_25280_, _25279_, _25276_);
  and (_25281_, _25280_, _24330_);
  or (_25282_, _25237_, _23205_);
  or (_25283_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25284_, _25283_, _22915_);
  and (_25285_, _25284_, _25282_);
  not (_25287_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_25288_, _22914_, _25287_);
  or (_25289_, _25288_, rst);
  or (_25290_, _25289_, _25285_);
  or (_15120_, _25290_, _25281_);
  and (_25291_, _25226_, _24184_);
  or (_25292_, _25291_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25293_, _25292_, _24330_);
  nand (_25294_, _25291_, _23681_);
  and (_25295_, _25294_, _25293_);
  or (_25297_, _25237_, _23247_);
  or (_25298_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25299_, _25298_, _22915_);
  and (_25300_, _25299_, _25297_);
  and (_25301_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_25302_, _25301_, rst);
  or (_25303_, _25302_, _25300_);
  or (_15135_, _25303_, _25295_);
  and (_25304_, _25220_, _23900_);
  and (_25305_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_15235_, _25305_, _25304_);
  and (_25306_, _25220_, _23983_);
  and (_25307_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_15250_, _25307_, _25306_);
  and (_25308_, _24157_, _24084_);
  not (_25309_, _25308_);
  and (_25310_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and (_25311_, _25308_, _24027_);
  or (_15265_, _25311_, _25310_);
  and (_25312_, _25180_, _24053_);
  and (_25313_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or (_15283_, _25313_, _25312_);
  nor (_25314_, _22809_, _22926_);
  and (_25315_, _25314_, _22855_);
  and (_25316_, _25315_, _24758_);
  and (_25317_, _25316_, _24405_);
  nand (_25318_, _25317_, _23681_);
  and (_25319_, _22822_, _23426_);
  and (_25320_, _25319_, _22856_);
  and (_25321_, _25320_, _25235_);
  or (_25322_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_25323_, _25322_, _24330_);
  and (_25324_, _25323_, _25318_);
  nand (_25325_, _25321_, _24047_);
  and (_25326_, _25322_, _22915_);
  and (_25327_, _25326_, _25325_);
  not (_25328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_25329_, _22914_, _25328_);
  or (_25330_, _25329_, rst);
  or (_25331_, _25330_, _25327_);
  or (_15324_, _25331_, _25324_);
  and (_25332_, _25180_, _23693_);
  and (_25333_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or (_27137_, _25333_, _25332_);
  and (_25334_, _25180_, _23715_);
  and (_25335_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or (_15465_, _25335_, _25334_);
  and (_25336_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and (_25337_, _25308_, _23920_);
  or (_15486_, _25337_, _25336_);
  and (_25338_, _25194_, _23715_);
  and (_25339_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_15507_, _25339_, _25338_);
  and (_25340_, _25194_, _23900_);
  and (_25341_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_15748_, _25341_, _25340_);
  and (_25342_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and (_25343_, _25308_, _23900_);
  or (_15769_, _25343_, _25342_);
  and (_25344_, _25194_, _24027_);
  and (_25345_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_15790_, _25345_, _25344_);
  and (_25346_, _24388_, _24061_);
  and (_25347_, _25346_, _23693_);
  not (_25348_, _25346_);
  and (_25349_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or (_15881_, _25349_, _25347_);
  and (_25350_, _25346_, _23715_);
  and (_25351_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or (_15952_, _25351_, _25350_);
  and (_25352_, _25346_, _23920_);
  and (_25353_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or (_16003_, _25353_, _25352_);
  and (_25354_, _25346_, _23983_);
  and (_25355_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or (_27163_, _25355_, _25354_);
  and (_25356_, _24388_, _23930_);
  and (_25357_, _25356_, _23751_);
  not (_25358_, _25356_);
  and (_25359_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or (_16112_, _25359_, _25357_);
  and (_25360_, _25356_, _23715_);
  and (_25361_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or (_27165_, _25361_, _25360_);
  and (_25362_, _23920_, _23892_);
  and (_25363_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or (_16477_, _25363_, _25362_);
  and (_25364_, _23930_, _23719_);
  and (_25365_, _25364_, _23983_);
  not (_25367_, _25364_);
  and (_25368_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or (_16505_, _25368_, _25365_);
  and (_25369_, _25356_, _23920_);
  and (_25370_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or (_16999_, _25370_, _25369_);
  and (_25372_, _25356_, _24027_);
  and (_25373_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or (_17181_, _25373_, _25372_);
  nor (_25374_, _23760_, _23123_);
  and (_25375_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_25376_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_25378_, _25376_, _25375_);
  and (_25379_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_25380_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_25381_, _25380_, _25379_);
  and (_25382_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_25383_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_25384_, _25383_, _25382_);
  and (_25385_, _25384_, _25381_);
  and (_25386_, _25385_, _25378_);
  nor (_25387_, _25386_, _24817_);
  nor (_25388_, _25387_, _25374_);
  nor (_26858_[2], _25388_, rst);
  and (_25389_, _24388_, _23444_);
  and (_25390_, _25389_, _24053_);
  not (_25392_, _25389_);
  and (_25393_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_17511_, _25393_, _25390_);
  and (_25394_, _25389_, _23693_);
  and (_25395_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_17562_, _25395_, _25394_);
  and (_25396_, _25389_, _23900_);
  and (_25397_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_17583_, _25397_, _25396_);
  and (_25398_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_25399_, _25153_, _24053_);
  or (_17634_, _25399_, _25398_);
  and (_25400_, _25389_, _23920_);
  and (_25401_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_17655_, _25401_, _25400_);
  and (_25402_, _24388_, _23905_);
  and (_25403_, _25402_, _24053_);
  not (_25404_, _25402_);
  and (_25405_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_18277_, _25405_, _25403_);
  and (_25406_, _25402_, _23693_);
  and (_25407_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_27170_, _25407_, _25406_);
  and (_25408_, _25402_, _23900_);
  and (_25409_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_18497_, _25409_, _25408_);
  and (_25410_, _25364_, _23900_);
  and (_25411_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or (_19899_, _25411_, _25410_);
  and (_25412_, _25364_, _23920_);
  and (_25413_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or (_19933_, _25413_, _25412_);
  nor (_25414_, _23760_, _23133_);
  and (_25415_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_25416_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_25417_, _25416_, _25415_);
  and (_25418_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_25419_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_25420_, _25419_, _25418_);
  and (_25421_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_25422_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_25423_, _25422_, _25421_);
  and (_25424_, _25423_, _25420_);
  and (_25425_, _25424_, _25417_);
  nor (_25426_, _25425_, _24817_);
  nor (_25427_, _25426_, _25414_);
  nor (_26858_[1], _25427_, rst);
  and (_25428_, _23890_, _23453_);
  and (_25429_, _25428_, _23751_);
  not (_25430_, _25428_);
  and (_25431_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_20019_, _25431_, _25429_);
  and (_25432_, _24098_, _23920_);
  and (_25433_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or (_20200_, _25433_, _25432_);
  and (_25434_, _25402_, _23920_);
  and (_25435_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_20227_, _25435_, _25434_);
  and (_25436_, _24388_, _24274_);
  and (_25437_, _25436_, _23751_);
  not (_25438_, _25436_);
  and (_25439_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or (_27172_, _25439_, _25437_);
  and (_25440_, _24108_, _23453_);
  and (_25441_, _25440_, _23900_);
  not (_25442_, _25440_);
  and (_25443_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or (_27206_, _25443_, _25441_);
  and (_25444_, _25436_, _23715_);
  and (_25445_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or (_27173_, _25445_, _25444_);
  and (_25446_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  and (_25447_, _25308_, _23983_);
  or (_27006_, _25447_, _25446_);
  and (_25448_, _25440_, _23715_);
  and (_25449_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or (_27205_, _25449_, _25448_);
  and (_25450_, _25436_, _23900_);
  and (_25451_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or (_27174_, _25451_, _25450_);
  and (_25452_, _25436_, _23983_);
  and (_25453_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or (_27176_, _25453_, _25452_);
  and (_25454_, _24388_, _24145_);
  and (_25455_, _25454_, _24053_);
  not (_25456_, _25454_);
  and (_25457_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or (_27179_, _25457_, _25455_);
  nor (_26831_[6], _24537_, rst);
  and (_25458_, _25454_, _23693_);
  and (_25459_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or (_27180_, _25459_, _25458_);
  nor (_25460_, _23760_, _23300_);
  and (_25461_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_25462_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_25463_, _25462_, _25461_);
  and (_25464_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_25465_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_25466_, _25465_, _25464_);
  and (_25467_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_25468_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_25469_, _25468_, _25467_);
  and (_25470_, _25469_, _25466_);
  and (_25471_, _25470_, _25463_);
  nor (_25472_, _25471_, _24817_);
  nor (_25473_, _25472_, _25460_);
  nor (_26858_[5], _25473_, rst);
  and (_25474_, _25454_, _23900_);
  and (_25475_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or (_27181_, _25475_, _25474_);
  and (_25476_, _25454_, _24027_);
  and (_25477_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or (_27183_, _25477_, _25476_);
  and (_25478_, _23925_, _23715_);
  and (_25479_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_27247_, _25479_, _25478_);
  and (_25480_, _24389_, _23751_);
  and (_25481_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_27186_, _25481_, _25480_);
  and (_25482_, _24235_, _23891_);
  and (_25483_, _25482_, _23693_);
  not (_25484_, _25482_);
  and (_25485_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_27227_, _25485_, _25483_);
  and (_25486_, _24389_, _23715_);
  and (_25487_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_27187_, _25487_, _25486_);
  and (_25488_, _25165_, _23715_);
  and (_25489_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_26935_, _25489_, _25488_);
  and (_25490_, _24123_, _24084_);
  not (_25491_, _25490_);
  and (_25492_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_25493_, _25490_, _23983_);
  or (_27004_, _25493_, _25492_);
  and (_25494_, _25165_, _23693_);
  and (_25495_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_26934_, _25495_, _25494_);
  and (_25496_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_25497_, _25490_, _24027_);
  or (_27003_, _25497_, _25496_);
  and (_25499_, _25159_, _23693_);
  and (_25500_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or (_27192_, _25500_, _25499_);
  and (_25501_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_25502_, _25490_, _23920_);
  or (_27002_, _25502_, _25501_);
  and (_25503_, _25164_, _23444_);
  and (_25504_, _25503_, _23900_);
  not (_25505_, _25503_);
  and (_25506_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_26921_, _25506_, _25504_);
  and (_25507_, _25503_, _23715_);
  and (_25508_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_26920_, _25508_, _25507_);
  and (_25509_, _25503_, _23693_);
  and (_25510_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_26919_, _25510_, _25509_);
  and (_26856_[0], _24565_, _22773_);
  and (_26856_[1], _24637_, _22773_);
  and (_26856_[2], _24591_, _22773_);
  and (_25511_, _24342_, _24405_);
  and (_25512_, _25511_, _25319_);
  and (_25513_, _25512_, _23907_);
  not (_25514_, _25513_);
  and (_25515_, _25514_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_25516_, _25319_, _23907_);
  and (_25517_, _25516_, _25511_);
  and (_25518_, _25517_, _23413_);
  nor (_25519_, _25518_, _25515_);
  nor (_26856_[3], _25519_, rst);
  and (_25520_, _25503_, _23751_);
  and (_25521_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_26918_, _25521_, _25520_);
  nor (_25522_, _24477_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_25523_, _25522_, _24883_);
  nor (_25524_, _25523_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_25525_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  not (_25526_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand (_25527_, _25524_, _25526_);
  and (_25528_, _25527_, _22773_);
  and (_26874_[0], _25528_, _25525_);
  or (_25529_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  not (_25530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_25531_, _25524_, _25530_);
  and (_25532_, _25531_, _22773_);
  and (_26874_[1], _25532_, _25529_);
  or (_25533_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  not (_25534_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_25535_, _25524_, _25534_);
  and (_25536_, _25535_, _22773_);
  and (_26874_[2], _25536_, _25533_);
  or (_25537_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not (_25538_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand (_25539_, _25524_, _25538_);
  and (_25540_, _25539_, _22773_);
  and (_26874_[3], _25540_, _25537_);
  or (_25541_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not (_25542_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand (_25543_, _25524_, _25542_);
  and (_25544_, _25543_, _22773_);
  and (_26874_[4], _25544_, _25541_);
  or (_25545_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not (_25546_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_25547_, _25524_, _25546_);
  and (_25548_, _25547_, _22773_);
  and (_26874_[5], _25548_, _25545_);
  or (_25550_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  not (_25551_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_25552_, _25524_, _25551_);
  and (_25554_, _25552_, _22773_);
  and (_26874_[6], _25554_, _25550_);
  or (_25556_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  not (_25557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand (_25558_, _25524_, _25557_);
  and (_25559_, _25558_, _22773_);
  and (_26874_[7], _25559_, _25556_);
  or (_25560_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not (_25561_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_25562_, _25524_, _25561_);
  and (_25564_, _25562_, _22773_);
  and (_26874_[8], _25564_, _25560_);
  or (_25565_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  not (_25566_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_25567_, _25524_, _25566_);
  and (_25568_, _25567_, _22773_);
  and (_26874_[9], _25568_, _25565_);
  or (_25569_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  not (_25570_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_25571_, _25524_, _25570_);
  and (_25572_, _25571_, _22773_);
  and (_26874_[10], _25572_, _25569_);
  or (_25573_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  not (_25574_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_25575_, _25524_, _25574_);
  and (_25576_, _25575_, _22773_);
  and (_26874_[11], _25576_, _25573_);
  or (_25577_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  not (_25578_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand (_25579_, _25524_, _25578_);
  and (_25580_, _25579_, _22773_);
  and (_26874_[12], _25580_, _25577_);
  or (_25581_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not (_25582_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_25583_, _25524_, _25582_);
  and (_25584_, _25583_, _22773_);
  and (_26874_[13], _25584_, _25581_);
  or (_25585_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  not (_25586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_25587_, _25524_, _25586_);
  and (_25589_, _25587_, _22773_);
  and (_26874_[14], _25589_, _25585_);
  and (_25590_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not (_25591_, _25524_);
  and (_25592_, _25591_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  or (_25593_, _25592_, _25590_);
  and (_26874_[15], _25593_, _22773_);
  or (_25594_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  not (_25595_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_25596_, _25524_, _25595_);
  and (_25597_, _25596_, _22773_);
  and (_26874_[16], _25597_, _25594_);
  or (_25599_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not (_25600_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_25601_, _25524_, _25600_);
  and (_25603_, _25601_, _22773_);
  and (_26874_[17], _25603_, _25599_);
  or (_25604_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not (_25605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_25606_, _25524_, _25605_);
  and (_25607_, _25606_, _22773_);
  and (_26874_[18], _25607_, _25604_);
  or (_25608_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not (_25609_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_25610_, _25524_, _25609_);
  and (_25611_, _25610_, _22773_);
  and (_26874_[19], _25611_, _25608_);
  or (_25612_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  not (_25613_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_25614_, _25524_, _25613_);
  and (_25615_, _25614_, _22773_);
  and (_26874_[20], _25615_, _25612_);
  or (_25617_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  not (_25618_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_25619_, _25524_, _25618_);
  and (_25620_, _25619_, _22773_);
  and (_26874_[21], _25620_, _25617_);
  or (_25621_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not (_25622_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_25623_, _25524_, _25622_);
  and (_25624_, _25623_, _22773_);
  and (_26874_[22], _25624_, _25621_);
  and (_25625_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_25626_, _25591_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or (_25627_, _25626_, _25625_);
  and (_26874_[23], _25627_, _22773_);
  or (_25628_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  not (_25630_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_25631_, _25524_, _25630_);
  and (_25632_, _25631_, _22773_);
  and (_26874_[24], _25632_, _25628_);
  or (_25633_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  not (_25634_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_25635_, _25524_, _25634_);
  and (_25636_, _25635_, _22773_);
  and (_26874_[25], _25636_, _25633_);
  or (_25637_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not (_25638_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_25639_, _25524_, _25638_);
  and (_25640_, _25639_, _22773_);
  and (_26874_[26], _25640_, _25637_);
  or (_25641_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not (_25642_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_25643_, _25524_, _25642_);
  and (_25644_, _25643_, _22773_);
  and (_26874_[27], _25644_, _25641_);
  or (_25645_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  not (_25646_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_25647_, _25524_, _25646_);
  and (_25648_, _25647_, _22773_);
  and (_26874_[28], _25648_, _25645_);
  or (_25649_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not (_25650_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_25651_, _25524_, _25650_);
  and (_25652_, _25651_, _22773_);
  and (_26874_[29], _25652_, _25649_);
  or (_25653_, _25524_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not (_25654_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_25655_, _25524_, _25654_);
  and (_25656_, _25655_, _22773_);
  and (_26874_[30], _25656_, _25653_);
  and (_25657_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and (_25658_, _25308_, _23693_);
  or (_22676_, _25658_, _25657_);
  and (_25659_, _25514_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_25660_, _25517_, _23205_);
  nor (_25661_, _25660_, _25659_);
  nor (_25662_, _25661_, _22809_);
  and (_25663_, _25661_, _22809_);
  nor (_25664_, _25663_, _25662_);
  not (_25665_, _25664_);
  nor (_25666_, _25519_, _22908_);
  and (_25667_, _25519_, _22908_);
  nor (_25668_, _25667_, _25666_);
  nor (_25670_, _24565_, _22869_);
  and (_25671_, _24565_, _22869_);
  nor (_25672_, _25671_, _25670_);
  and (_25673_, _22912_, _22910_);
  not (_25674_, _25673_);
  nand (_25676_, _22894_, _22881_);
  nor (_25677_, _25676_, _25674_);
  and (_25678_, _25677_, _22822_);
  and (_25680_, _25678_, _23450_);
  and (_25681_, _25680_, _25672_);
  not (_25682_, _25681_);
  nor (_25683_, _25682_, _25668_);
  and (_25684_, _25683_, _25665_);
  not (_25685_, _25661_);
  nor (_25686_, _25519_, _24566_);
  and (_25687_, _25686_, _25685_);
  and (_25688_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_25689_, _25519_, _24565_);
  and (_25690_, _25689_, _25685_);
  and (_25691_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_25692_, _25691_, _25688_);
  and (_25693_, _25519_, _24565_);
  and (_25694_, _25693_, _25685_);
  and (_25695_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_25696_, _25693_, _25661_);
  and (_25697_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_25698_, _25697_, _25695_);
  and (_25700_, _25698_, _25692_);
  and (_25701_, _25519_, _24566_);
  and (_25702_, _25701_, _25661_);
  and (_25703_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_25704_, _25686_, _25661_);
  and (_25705_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_25706_, _25705_, _25703_);
  and (_25707_, _25689_, _25661_);
  and (_25708_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_25709_, _25701_, _25685_);
  and (_25710_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_25711_, _25710_, _25708_);
  and (_25712_, _25711_, _25706_);
  and (_25713_, _25712_, _25700_);
  nor (_25714_, _25713_, _25684_);
  and (_25715_, _25684_, _24788_);
  nor (_25716_, _25715_, _25714_);
  nor (_26857_[0], _25716_, rst);
  and (_25717_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_25718_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_25719_, _25718_, _25717_);
  and (_25720_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_25721_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_25723_, _25721_, _25720_);
  and (_25725_, _25723_, _25719_);
  and (_25726_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_25727_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_25728_, _25727_, _25726_);
  and (_25729_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_25730_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_25731_, _25730_, _25729_);
  and (_25732_, _25731_, _25728_);
  and (_25733_, _25732_, _25725_);
  nor (_25734_, _25733_, _25684_);
  and (_25735_, _25684_, _23744_);
  nor (_25736_, _25735_, _25734_);
  nor (_26857_[1], _25736_, rst);
  and (_25737_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_25738_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_25739_, _25738_, _25737_);
  and (_25740_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_25741_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_25742_, _25741_, _25740_);
  and (_25743_, _25742_, _25739_);
  and (_25744_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_25745_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_25746_, _25745_, _25744_);
  and (_25747_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_25748_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_25749_, _25748_, _25747_);
  and (_25750_, _25749_, _25746_);
  and (_25751_, _25750_, _25743_);
  nor (_25752_, _25751_, _25684_);
  and (_25753_, _25684_, _23247_);
  nor (_25754_, _25753_, _25752_);
  nor (_26857_[2], _25754_, rst);
  and (_25755_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_25756_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_25757_, _25756_, _25755_);
  and (_25758_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_25759_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_25761_, _25759_, _25758_);
  and (_25762_, _25761_, _25757_);
  and (_25763_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_25764_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_25765_, _25764_, _25763_);
  and (_25766_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_25767_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_25768_, _25767_, _25766_);
  and (_25769_, _25768_, _25765_);
  and (_25771_, _25769_, _25762_);
  nor (_25773_, _25771_, _25684_);
  and (_25774_, _25684_, _23413_);
  nor (_25775_, _25774_, _25773_);
  nor (_26857_[3], _25775_, rst);
  and (_25776_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_25777_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_25778_, _25777_, _25776_);
  and (_25779_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_25780_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_25781_, _25780_, _25779_);
  and (_25782_, _25781_, _25778_);
  and (_25784_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_25785_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_25786_, _25785_, _25784_);
  and (_25787_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_25789_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_25790_, _25789_, _25787_);
  and (_25791_, _25790_, _25786_);
  and (_25792_, _25791_, _25782_);
  nor (_25794_, _25792_, _25684_);
  and (_25795_, _25684_, _23205_);
  nor (_25796_, _25795_, _25794_);
  nor (_26857_[4], _25796_, rst);
  and (_25797_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_25798_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_25799_, _25798_, _25797_);
  and (_25800_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_25801_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_25802_, _25801_, _25800_);
  and (_25803_, _25802_, _25799_);
  and (_25804_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_25805_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_25806_, _25805_, _25804_);
  and (_25807_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_25808_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_25809_, _25808_, _25807_);
  and (_25810_, _25809_, _25806_);
  and (_25811_, _25810_, _25803_);
  nor (_25812_, _25811_, _25684_);
  not (_25813_, _23357_);
  and (_25814_, _25684_, _25813_);
  nor (_25815_, _25814_, _25812_);
  nor (_26857_[5], _25815_, rst);
  and (_25816_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_25817_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_25818_, _25817_, _25816_);
  and (_25820_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_25821_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_25822_, _25821_, _25820_);
  and (_25823_, _25822_, _25818_);
  and (_25824_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_25825_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_25826_, _25825_, _25824_);
  and (_25827_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_25828_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_25829_, _25828_, _25827_);
  and (_25830_, _25829_, _25826_);
  and (_25831_, _25830_, _25823_);
  nor (_25832_, _25831_, _25684_);
  not (_25833_, _24017_);
  and (_25835_, _25684_, _25833_);
  nor (_25836_, _25835_, _25832_);
  nor (_26857_[6], _25836_, rst);
  and (_25837_, _25190_, _24053_);
  and (_25838_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_22677_, _25838_, _25837_);
  and (_25840_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  and (_25841_, _25308_, _23751_);
  or (_22678_, _25841_, _25840_);
  and (_25842_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and (_25843_, _25308_, _24053_);
  or (_22679_, _25843_, _25842_);
  and (_25844_, _25503_, _24027_);
  and (_25845_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_22680_, _25845_, _25844_);
  and (_25846_, _25503_, _23920_);
  and (_25847_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_26922_, _25847_, _25846_);
  and (_25848_, \oc8051_top_1.oc8051_decoder1.state [0], _22781_);
  and (_25849_, _24724_, _24669_);
  and (_25850_, _25849_, _24721_);
  and (_25851_, _24721_, _24543_);
  nor (_25852_, _25851_, _25850_);
  nor (_25853_, _25852_, _25848_);
  and (_25854_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_25855_, _24688_, _24591_);
  and (_25856_, _24720_, _25855_);
  and (_25857_, _25856_, _24709_);
  and (_25858_, _25856_, _24674_);
  nor (_25859_, _25858_, _25857_);
  nor (_25860_, _25859_, _24646_);
  and (_25861_, _25859_, _24685_);
  nor (_25862_, _25861_, _24647_);
  and (_25863_, _24721_, _24680_);
  and (_25864_, _25863_, _24733_);
  or (_25865_, _25864_, _25862_);
  nor (_25866_, _25865_, _25860_);
  nor (_25867_, _25866_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_25868_, _25867_, _25854_);
  and (_25869_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_25870_, _24738_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_25871_, _25870_, _25869_);
  not (_25872_, _25871_);
  and (_25873_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_25874_, _25873_);
  and (_25875_, _24639_, _24712_);
  and (_25876_, _24687_, _24670_);
  and (_25877_, _25876_, _24639_);
  nor (_25878_, _25877_, _25875_);
  and (_25879_, _24639_, _24682_);
  and (_25880_, _24721_, _24673_);
  and (_25881_, _25880_, _24670_);
  nor (_25882_, _25881_, _25879_);
  and (_25883_, _25882_, _25878_);
  and (_25884_, _25880_, _24669_);
  not (_25885_, _25884_);
  nor (_25886_, _24637_, _24566_);
  and (_25887_, _25886_, _25855_);
  and (_25888_, _25887_, _24722_);
  and (_25889_, _25887_, _25849_);
  nor (_25890_, _25889_, _25888_);
  and (_25891_, _25887_, _24699_);
  and (_25892_, _24699_, _24638_);
  nor (_25893_, _25892_, _25891_);
  and (_25894_, _25893_, _25890_);
  and (_25895_, _25894_, _25885_);
  and (_25896_, _25895_, _25883_);
  and (_25897_, _24639_, _24678_);
  and (_25898_, _24722_, _24638_);
  and (_25899_, _25898_, _24566_);
  nor (_25900_, _25899_, _25897_);
  and (_25901_, _24639_, _24709_);
  and (_25902_, _24704_, _24638_);
  nor (_25903_, _25902_, _25901_);
  and (_25904_, _24721_, _24687_);
  and (_25905_, _24715_, _24638_);
  nor (_25906_, _25905_, _25904_);
  and (_25907_, _25887_, _24712_);
  and (_25908_, _25887_, _24678_);
  nor (_25909_, _25908_, _25907_);
  and (_25910_, _25909_, _25906_);
  and (_25911_, _25910_, _25903_);
  and (_25912_, _25911_, _25900_);
  and (_25913_, _25887_, _24715_);
  and (_25914_, _25887_, _25876_);
  nor (_25915_, _25914_, _25913_);
  not (_25916_, _25915_);
  not (_25917_, _25887_);
  nor (_25918_, _25917_, _24705_);
  nor (_25919_, _25918_, _25916_);
  and (_25920_, _24639_, _24674_);
  and (_25921_, _24690_, _24674_);
  nor (_25922_, _25921_, _25920_);
  and (_25923_, _25922_, _25919_);
  nor (_25924_, _24669_, _24688_);
  and (_25925_, _25924_, _24673_);
  and (_25926_, _25887_, _24697_);
  nor (_25928_, _25926_, _25925_);
  and (_25929_, _25887_, _24709_);
  and (_25930_, _24724_, _24670_);
  and (_25931_, _25930_, _25887_);
  nor (_25932_, _25931_, _25929_);
  and (_25933_, _25932_, _25928_);
  and (_25934_, _25852_, _24719_);
  and (_25936_, _25934_, _25933_);
  and (_25937_, _25936_, _25923_);
  and (_25938_, _25937_, _25912_);
  nand (_25939_, _25938_, _25896_);
  nand (_25940_, _25939_, _24646_);
  nor (_25941_, _25864_, _24643_);
  nand (_25942_, _25941_, _25940_);
  nand (_25943_, _25942_, _22781_);
  and (_25944_, _25943_, _25874_);
  and (_25945_, _25944_, _25872_);
  and (_25946_, _25945_, _25868_);
  not (_25947_, _25946_);
  nor (_25948_, _25947_, _25796_);
  not (_25949_, _25948_);
  nor (_25951_, _25944_, _25871_);
  and (_25952_, _25951_, _25868_);
  not (_25953_, _25952_);
  and (_25954_, _25234_, _22882_);
  and (_25955_, _25954_, _22928_);
  and (_25956_, _25955_, _23205_);
  and (_25957_, _25955_, _23247_);
  not (_25958_, _25955_);
  and (_25959_, _25958_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_25960_, _25959_, _25957_);
  and (_25961_, _25955_, _23744_);
  and (_25962_, _25958_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_25963_, _25962_, _25961_);
  or (_25964_, _25955_, _22864_);
  nand (_25965_, _25955_, _24788_);
  and (_25966_, _25965_, _25964_);
  and (_25967_, _25966_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_25968_, _25967_, _25963_);
  and (_25969_, _25968_, _25960_);
  and (_25970_, _25955_, _23413_);
  and (_25971_, _25958_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_25972_, _25971_, _25970_);
  and (_25973_, _25972_, _25969_);
  and (_25974_, _25958_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_25975_, _25974_, _25956_);
  and (_25976_, _25975_, _25973_);
  nor (_25977_, _25975_, _25973_);
  nor (_25978_, _25977_, _25976_);
  nor (_25979_, _25978_, _22784_);
  nor (_25980_, _25979_, _22789_);
  nor (_25981_, _25980_, _25955_);
  nor (_25982_, _25981_, _25956_);
  nor (_25983_, _25982_, _25953_);
  not (_25984_, _25983_);
  and (_25985_, _25871_, _25868_);
  and (_25986_, _25985_, _25944_);
  and (_25987_, _25986_, _25685_);
  not (_25988_, _25987_);
  nor (_25989_, _25944_, _25872_);
  nor (_25990_, _23760_, _22952_);
  and (_25991_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_25992_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_25993_, _25992_, _25991_);
  and (_25994_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_25995_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_25996_, _25995_, _25994_);
  and (_25997_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_25998_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_25999_, _25998_, _25997_);
  and (_26001_, _25999_, _25996_);
  and (_26002_, _26001_, _25993_);
  nor (_26003_, _26002_, _24817_);
  nor (_26004_, _26003_, _25990_);
  not (_26005_, _26004_);
  and (_26006_, _26005_, _25989_);
  not (_26007_, _25868_);
  and (_26008_, _25871_, _26007_);
  nor (_26009_, _26008_, _26006_);
  and (_26010_, _26009_, _25988_);
  and (_26012_, _26010_, _25984_);
  and (_26013_, _26012_, _25949_);
  nor (_26014_, _26013_, _22809_);
  and (_26016_, _26013_, _22809_);
  nor (_26017_, _26016_, _26014_);
  nor (_26018_, _25947_, _25815_);
  not (_26019_, _25473_);
  not (_26021_, _25944_);
  and (_26022_, _25985_, _26021_);
  and (_26023_, _26022_, _26019_);
  nor (_26024_, _26023_, _26018_);
  nor (_26025_, _25958_, _23357_);
  and (_26026_, _25958_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_26027_, _26026_, _26025_);
  and (_26028_, _26027_, _25976_);
  nor (_26030_, _26027_, _25976_);
  nor (_26031_, _26030_, _26028_);
  nor (_26032_, _26031_, _22784_);
  nor (_26033_, _26032_, _22814_);
  nor (_26034_, _26033_, _25955_);
  nor (_26035_, _26034_, _26025_);
  nor (_26036_, _26035_, _25953_);
  not (_26037_, _25989_);
  nor (_26038_, _25945_, _25868_);
  and (_26039_, _26038_, _26037_);
  nor (_26040_, _26039_, _26036_);
  and (_26041_, _26040_, _26024_);
  nor (_26042_, _26041_, _22822_);
  and (_26043_, _26041_, _22822_);
  nor (_26044_, _26043_, _26042_);
  nor (_26045_, _26044_, _26017_);
  nor (_26046_, _25947_, _25775_);
  not (_26047_, _26046_);
  nor (_26048_, _25972_, _25969_);
  nor (_26049_, _26048_, _25973_);
  nor (_26050_, _26049_, _22784_);
  nor (_26051_, _26050_, _22899_);
  nor (_26052_, _26051_, _25955_);
  nor (_26053_, _26052_, _25970_);
  not (_26054_, _26053_);
  nand (_26055_, _26054_, _25952_);
  not (_26056_, _25519_);
  and (_26057_, _25986_, _26056_);
  nor (_26058_, _23760_, _23086_);
  and (_26059_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_26060_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_26061_, _26060_, _26059_);
  and (_26062_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_26063_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_26064_, _26063_, _26062_);
  and (_26065_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_26066_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_26067_, _26066_, _26065_);
  and (_26068_, _26067_, _26064_);
  and (_26069_, _26068_, _26061_);
  nor (_26070_, _26069_, _24817_);
  nor (_26071_, _26070_, _26058_);
  not (_26072_, _26071_);
  and (_26073_, _26072_, _26022_);
  nor (_26074_, _26073_, _26057_);
  and (_26075_, _26074_, _26055_);
  and (_26076_, _26075_, _26047_);
  nor (_26077_, _26076_, _22908_);
  and (_26078_, _26076_, _22908_);
  nor (_26079_, _26078_, _26077_);
  not (_26080_, _26079_);
  nor (_26081_, _25958_, _24017_);
  and (_26082_, _25958_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_26083_, _26082_, _26081_);
  and (_26084_, _26083_, _26028_);
  nor (_26086_, _26083_, _26028_);
  nor (_26087_, _26086_, _26084_);
  nor (_26088_, _26087_, _22784_);
  nor (_26089_, _26088_, _22828_);
  nor (_26090_, _26089_, _25955_);
  nor (_26091_, _26090_, _26081_);
  nor (_26092_, _26091_, _25953_);
  nor (_26093_, _25947_, _25836_);
  nor (_26094_, _23760_, _23498_);
  and (_26095_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_26096_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_26097_, _26096_, _26095_);
  and (_26098_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_26099_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_26100_, _26099_, _26098_);
  and (_26101_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_26102_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_26103_, _26102_, _26101_);
  and (_26104_, _26103_, _26100_);
  and (_26105_, _26104_, _26097_);
  nor (_26106_, _26105_, _24817_);
  nor (_26107_, _26106_, _26094_);
  not (_26108_, _26107_);
  and (_26109_, _26108_, _25989_);
  or (_26110_, _26109_, _26093_);
  or (_26111_, _26110_, _26092_);
  nor (_26112_, _26111_, _26038_);
  nor (_26113_, _26112_, _22838_);
  and (_26114_, _26112_, _22838_);
  nor (_26116_, _26114_, _26113_);
  and (_26117_, _25955_, _23976_);
  and (_26118_, _25958_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_26119_, _26118_, _26084_);
  or (_26120_, _26118_, _26084_);
  and (_26121_, _26120_, _22785_);
  nand (_26122_, _26121_, _26119_);
  nor (_26123_, _25955_, _22842_);
  and (_26124_, _26123_, _26122_);
  nor (_26125_, _26124_, _26117_);
  nand (_26126_, _26125_, _25952_);
  not (_26127_, _25684_);
  nand (_26128_, _25707_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nand (_26129_, _25702_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_26130_, _26129_, _26128_);
  nand (_26131_, _25709_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nand (_26132_, _25687_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_26133_, _26132_, _26131_);
  and (_26134_, _26133_, _26130_);
  nand (_26135_, _25690_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand (_26136_, _25694_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_26137_, _26136_, _26135_);
  nand (_26138_, _25704_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand (_26139_, _25696_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_26140_, _26139_, _26138_);
  and (_26142_, _26140_, _26137_);
  nand (_26143_, _26142_, _26134_);
  nand (_26144_, _26143_, _26127_);
  not (_26145_, _23976_);
  nand (_26146_, _25684_, _26145_);
  nand (_26147_, _26146_, _26144_);
  nand (_26148_, _26147_, _25945_);
  not (_26149_, _24819_);
  nand (_26150_, _25989_, _26149_);
  and (_26151_, _26150_, _25868_);
  and (_26152_, _26151_, _26148_);
  nand (_26153_, _26152_, _26126_);
  and (_26154_, _26153_, _22855_);
  nor (_26155_, _26153_, _22855_);
  nor (_26156_, _26155_, _26154_);
  nor (_26157_, _26156_, _26116_);
  and (_26158_, _26157_, _26080_);
  and (_26160_, _26158_, _26045_);
  nor (_26161_, _24341_, _22917_);
  and (_26163_, _26161_, _26160_);
  and (_26164_, _26163_, _25853_);
  not (_26165_, _26164_);
  and (_26166_, _24724_, _24639_);
  and (_26167_, _25886_, _24616_);
  nor (_26168_, _26167_, _26166_);
  nor (_26169_, _26168_, _24647_);
  nor (_26170_, _23587_, _23188_);
  and (_26171_, _23587_, _23188_);
  nor (_26172_, _26171_, _26170_);
  not (_26174_, _26172_);
  nor (_26175_, _23589_, _23532_);
  nor (_26176_, _26175_, _23590_);
  and (_26177_, _26176_, _26174_);
  not (_26178_, _23492_);
  and (_26179_, _23591_, _26178_);
  nor (_26180_, _23591_, _26178_);
  nor (_26182_, _26180_, _26179_);
  nor (_26183_, _25864_, _25853_);
  nor (_26185_, _23588_, _23535_);
  nor (_26186_, _26185_, _23589_);
  nor (_26187_, _23581_, _23566_);
  nor (_26188_, _26187_, _23582_);
  and (_26189_, _23575_, _23046_);
  nor (_26190_, _26189_, _23608_);
  nor (_26191_, _23568_, _26190_);
  and (_26192_, _26191_, _26188_);
  and (_26193_, _26192_, _23579_);
  and (_26195_, _26193_, _26186_);
  nand (_26196_, _26195_, _26183_);
  nor (_26197_, _26196_, _26182_);
  and (_26198_, _26197_, _26177_);
  not (_26199_, _26198_);
  and (_26200_, _25853_, _23668_);
  not (_26201_, _26200_);
  nor (_26202_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_26204_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_26205_, _26204_, _26202_);
  nor (_26207_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_26208_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_26209_, _26208_, _26207_);
  and (_26210_, _26209_, _26205_);
  and (_26211_, _26210_, _24736_);
  not (_26212_, _25864_);
  nor (_26213_, _25853_, _24676_);
  nor (_26214_, _26213_, _26212_);
  and (_26215_, _26214_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_26216_, _26215_, _26211_);
  and (_26217_, _26216_, _26201_);
  and (_26219_, _26217_, _26199_);
  and (_26221_, _25851_, _24670_);
  not (_26222_, _26221_);
  and (_26223_, _25863_, _24670_);
  nor (_26224_, _26223_, _25850_);
  and (_26225_, _26224_, _26222_);
  not (_26226_, _26225_);
  nor (_26227_, _26226_, _26219_);
  or (_26228_, _25887_, _25856_);
  and (_26229_, _26228_, _24712_);
  nor (_26230_, _26229_, _25888_);
  and (_26231_, _24669_, _24615_);
  and (_26232_, _26231_, _24687_);
  not (_26234_, _26232_);
  and (_26236_, _26234_, _26230_);
  and (_26238_, _24712_, _24615_);
  nor (_26239_, _26238_, _24714_);
  not (_26240_, _26239_);
  not (_26241_, _24721_);
  nor (_26242_, _24704_, _24682_);
  nor (_26243_, _26242_, _26241_);
  nor (_26244_, _26243_, _26240_);
  and (_26245_, _25851_, _24669_);
  not (_26246_, _26245_);
  and (_26247_, _26246_, _26244_);
  and (_26249_, _26247_, _26236_);
  and (_26250_, _26249_, _26219_);
  nor (_26252_, _26250_, _26227_);
  and (_26253_, _24682_, _24648_);
  and (_26254_, _24721_, _24709_);
  or (_26255_, _26254_, _26253_);
  nor (_26256_, _26255_, _26252_);
  and (_26257_, _26256_, _24719_);
  nor (_26258_, _24733_, _24643_);
  nor (_26259_, _26258_, _26257_);
  nor (_26260_, _26259_, _26169_);
  not (_26261_, _24736_);
  not (_26262_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_26263_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _22781_);
  and (_26264_, _26263_, _26262_);
  not (_26265_, _26264_);
  not (_26266_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_26267_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _22781_);
  and (_26268_, _26267_, _26266_);
  and (_26269_, _24403_, _23907_);
  and (_26270_, _26269_, _25511_);
  nor (_26271_, _26270_, _26268_);
  and (_26272_, _26271_, _26265_);
  nor (_26273_, _22838_, _22822_);
  and (_26274_, _26273_, _24331_);
  and (_26275_, _26274_, _25224_);
  not (_26276_, _26275_);
  and (_26277_, _26276_, _26272_);
  nor (_26278_, _26277_, _26261_);
  nor (_26279_, _22838_, _23439_);
  and (_26281_, _26279_, _24330_);
  and (_26282_, _26281_, _25315_);
  nor (_26283_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_26284_, _26283_);
  nor (_26285_, _26284_, _26282_);
  and (_26286_, _26285_, _25514_);
  not (_26287_, _26286_);
  and (_26288_, _26287_, _26214_);
  nor (_26289_, _26288_, _26278_);
  not (_26290_, _26289_);
  nor (_26291_, _26290_, _26260_);
  not (_26292_, _26291_);
  nor (_26293_, _25947_, _25736_);
  not (_26294_, _26293_);
  and (_26295_, _25945_, _26007_);
  nor (_26296_, _25967_, _25963_);
  nor (_26297_, _26296_, _25968_);
  nor (_26298_, _26297_, _22784_);
  nor (_26300_, _26298_, _22873_);
  nor (_26301_, _26300_, _25955_);
  nor (_26302_, _26301_, _25961_);
  not (_26303_, _26302_);
  and (_26304_, _26303_, _25952_);
  or (_26305_, _26304_, _26295_);
  not (_26306_, _26305_);
  and (_26307_, _25986_, _24637_);
  not (_26308_, _25427_);
  and (_26309_, _26022_, _26308_);
  nor (_26310_, _26309_, _26307_);
  and (_26311_, _26310_, _26306_);
  and (_26312_, _26311_, _26294_);
  and (_26313_, _26312_, _24182_);
  nor (_26314_, _25947_, _25716_);
  not (_26315_, _26314_);
  and (_26317_, _25986_, _24565_);
  nor (_26318_, _25966_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_26319_, _26318_, _25967_);
  nor (_26320_, _26319_, _22784_);
  nor (_26321_, _26320_, _22865_);
  nor (_26322_, _26321_, _25955_);
  not (_26323_, _26322_);
  and (_26324_, _26323_, _25965_);
  not (_26325_, _26324_);
  and (_26326_, _26325_, _25952_);
  nor (_26327_, _23760_, _23097_);
  and (_26328_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_26329_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_26330_, _26329_, _26328_);
  and (_26331_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_26332_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_26333_, _26332_, _26331_);
  and (_26334_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_26335_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_26336_, _26335_, _26334_);
  and (_26337_, _26336_, _26333_);
  and (_26338_, _26337_, _26330_);
  nor (_26339_, _26338_, _24817_);
  nor (_26340_, _26339_, _26327_);
  not (_26341_, _26340_);
  and (_26342_, _26341_, _26022_);
  or (_26343_, _26342_, _26326_);
  nor (_26344_, _26343_, _26317_);
  and (_26345_, _26344_, _26315_);
  and (_26346_, _26345_, _22870_);
  nor (_26347_, _26312_, _24182_);
  or (_26348_, _26347_, _26346_);
  nor (_26349_, _26348_, _26313_);
  nor (_26350_, _25947_, _25754_);
  not (_26351_, _26350_);
  and (_26352_, _25986_, _24591_);
  nor (_26353_, _25968_, _25960_);
  nor (_26354_, _26353_, _25969_);
  nor (_26355_, _26354_, _22784_);
  nor (_26356_, _26355_, _22885_);
  nor (_26357_, _26356_, _25955_);
  nor (_26358_, _26357_, _25957_);
  not (_26359_, _26358_);
  and (_26360_, _26359_, _25952_);
  not (_26361_, _25388_);
  and (_26362_, _26022_, _26361_);
  or (_26363_, _26362_, _26360_);
  nor (_26364_, _26363_, _26352_);
  and (_26365_, _26364_, _26351_);
  nor (_26366_, _26365_, _23207_);
  nor (_26367_, _26366_, _25257_);
  nor (_26368_, _26345_, _22870_);
  and (_26369_, _26365_, _23207_);
  nor (_26370_, _26369_, _26368_);
  and (_26371_, _26370_, _26367_);
  and (_26372_, _26371_, _26349_);
  and (_26373_, _26372_, _26045_);
  and (_26374_, _26373_, _26158_);
  and (_26375_, _22855_, _22910_);
  and (_26376_, _26375_, _26374_);
  nor (_26377_, _26376_, _26292_);
  and (_26378_, _26377_, _26165_);
  and (_26379_, _23172_, _23167_);
  nor (_26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26381_, _26380_, _23109_);
  nor (_26382_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_26383_, _26382_, _26381_);
  and (_26384_, _23554_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_26385_, _26384_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26386_, _23520_, _23485_);
  nor (_26387_, _26386_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26388_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_26389_, _23217_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26390_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26391_, _23060_, _26390_);
  nand (_26392_, _26391_, _26389_);
  or (_26393_, _23388_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26394_, _23343_, _26390_);
  nand (_26395_, _26394_, _26393_);
  and (_26396_, _26395_, _26392_);
  or (_26397_, _23060_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26398_, _23518_, _26390_);
  nand (_26399_, _26398_, _26397_);
  or (_26400_, _23343_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26401_, _23485_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26402_, _26401_, _26400_);
  and (_26403_, _26402_, _26399_);
  nand (_26404_, _26403_, _26396_);
  and (_26405_, _26404_, _26388_);
  nor (_26406_, _26405_, _26387_);
  or (_26407_, _23545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26408_, _23388_, _26390_);
  nand (_26409_, _26408_, _26407_);
  and (_26410_, _26409_, _26388_);
  and (_26411_, _26402_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_26412_, _26411_, _26410_);
  nand (_26413_, _26380_, _23479_);
  nor (_26414_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_26415_, _26414_);
  and (_26416_, _26415_, _26413_);
  not (_26417_, _26416_);
  or (_26418_, _23554_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26419_, _23217_, _26390_);
  and (_26420_, _26419_, _26418_);
  or (_26421_, _26420_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26422_, _26399_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26423_, _26422_, _26421_);
  or (_26424_, _26423_, _26417_);
  and (_26425_, _23545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26426_, _26425_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26427_, _26395_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26428_, _26427_, _26426_);
  nand (_26429_, _26380_, _23511_);
  nor (_26430_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_26431_, _26430_);
  and (_26432_, _26431_, _26429_);
  not (_26433_, _26432_);
  or (_26434_, _26433_, _26428_);
  nand (_26435_, _26422_, _26421_);
  or (_26436_, _26435_, _26416_);
  and (_26437_, _26436_, _26424_);
  not (_26438_, _26437_);
  or (_26439_, _26438_, _26434_);
  and (_26440_, _26439_, _26424_);
  nand (_26441_, _26427_, _26426_);
  or (_26442_, _26432_, _26441_);
  and (_26443_, _26442_, _26434_);
  and (_26444_, _26443_, _26437_);
  not (_26445_, _26380_);
  or (_26446_, _26445_, _23313_);
  nor (_26447_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_26448_, _26447_);
  nand (_26449_, _26448_, _26446_);
  or (_26450_, _26384_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26451_, _26392_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26452_, _26451_, _26450_);
  or (_26453_, _26452_, _26449_);
  nor (_26454_, _26409_, _26388_);
  nand (_26455_, _26380_, _22976_);
  nor (_26456_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_26457_, _26456_);
  and (_26458_, _26457_, _26455_);
  not (_26459_, _26458_);
  or (_26460_, _26459_, _26454_);
  and (_26461_, _26448_, _26446_);
  nand (_26462_, _26451_, _26450_);
  or (_26463_, _26462_, _26461_);
  nand (_26464_, _26463_, _26453_);
  or (_26465_, _26464_, _26460_);
  nand (_26466_, _26465_, _26453_);
  nand (_26467_, _26466_, _26444_);
  and (_26468_, _26467_, _26440_);
  and (_26469_, _26420_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_26470_, _26469_);
  nand (_26471_, _26380_, _23091_);
  nor (_26472_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_26473_, _26472_);
  and (_26474_, _26473_, _26471_);
  nand (_26475_, _26474_, _26470_);
  or (_26476_, _26474_, _26470_);
  nand (_26477_, _26476_, _26475_);
  nand (_26478_, _26425_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_26479_, _26445_, _23128_);
  nor (_26480_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_26481_, _26480_);
  and (_26482_, _26481_, _26479_);
  nand (_26483_, _26482_, _26478_);
  or (_26484_, _26445_, _23147_);
  nor (_26485_, _26380_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_26486_, _26485_);
  nand (_26487_, _26486_, _26484_);
  and (_26488_, _26487_, _26385_);
  or (_26489_, _26482_, _26478_);
  nand (_26490_, _26489_, _26483_);
  or (_26491_, _26490_, _26488_);
  and (_26492_, _26491_, _26483_);
  or (_26493_, _26492_, _26477_);
  nand (_26494_, _26493_, _26475_);
  not (_26495_, _26454_);
  or (_26496_, _26458_, _26495_);
  and (_26497_, _26496_, _26460_);
  and (_26498_, _26463_, _26453_);
  and (_26499_, _26498_, _26497_);
  and (_26500_, _26499_, _26444_);
  nand (_26501_, _26500_, _26494_);
  nand (_26502_, _26501_, _26468_);
  not (_26503_, _26412_);
  and (_26504_, _26503_, _26406_);
  nand (_26505_, _26504_, _26502_);
  and (_26506_, _26505_, _26417_);
  not (_26507_, _26506_);
  and (_26508_, _26504_, _26502_);
  and (_26509_, _26452_, _26449_);
  and (_26510_, _26497_, _26494_);
  not (_26511_, _26510_);
  and (_26512_, _26511_, _26460_);
  or (_26513_, _26512_, _26509_);
  and (_26514_, _26513_, _26453_);
  not (_26515_, _26514_);
  nand (_26516_, _26515_, _26443_);
  nand (_26517_, _26516_, _26434_);
  nand (_26518_, _26517_, _26438_);
  nand (_26519_, _26518_, _26508_);
  nand (_26520_, _26519_, _26507_);
  or (_26521_, _26520_, _26412_);
  or (_26522_, _26515_, _26443_);
  nand (_26523_, _26522_, _26516_);
  nand (_26524_, _26523_, _26508_);
  and (_26525_, _26505_, _26433_);
  not (_26526_, _26525_);
  and (_26527_, _26526_, _26524_);
  nand (_26528_, _26527_, _26435_);
  and (_26529_, _26519_, _26507_);
  or (_26530_, _26529_, _26503_);
  and (_26531_, _26530_, _26521_);
  not (_26532_, _26531_);
  or (_26533_, _26532_, _26528_);
  and (_26534_, _26533_, _26521_);
  or (_26535_, _26527_, _26435_);
  and (_26536_, _26535_, _26528_);
  and (_26537_, _26536_, _26531_);
  nand (_26538_, _26464_, _26512_);
  or (_26539_, _26464_, _26512_);
  nand (_26540_, _26539_, _26538_);
  nand (_26541_, _26540_, _26508_);
  and (_26542_, _26505_, _26449_);
  not (_26543_, _26542_);
  and (_26544_, _26543_, _26541_);
  and (_26545_, _26544_, _26441_);
  nor (_26546_, _26497_, _26494_);
  nor (_26547_, _26546_, _26510_);
  nor (_26548_, _26547_, _26505_);
  and (_26549_, _26505_, _26459_);
  nor (_26550_, _26549_, _26548_);
  and (_26551_, _26550_, _26462_);
  not (_26552_, _26551_);
  nor (_26553_, _26544_, _26441_);
  or (_26554_, _26545_, _26553_);
  nor (_26555_, _26554_, _26552_);
  or (_26556_, _26555_, _26545_);
  and (_26557_, _26492_, _26477_);
  not (_26558_, _26557_);
  and (_26559_, _26558_, _26493_);
  or (_26560_, _26559_, _26505_);
  or (_26561_, _26508_, _26474_);
  and (_26562_, _26561_, _26560_);
  nor (_26563_, _26562_, _26495_);
  not (_26564_, _26563_);
  not (_26565_, _26385_);
  or (_26566_, _26505_, _26565_);
  nand (_26567_, _26566_, _26487_);
  or (_26568_, _26566_, _26487_);
  and (_26569_, _26568_, _26567_);
  nand (_26570_, _26569_, _26478_);
  or (_26571_, _26569_, _26478_);
  and (_26572_, _26571_, _26570_);
  nor (_26573_, _26565_, _26383_);
  not (_26574_, _26573_);
  nand (_26575_, _26574_, _26572_);
  and (_26576_, _26575_, _26570_);
  and (_26577_, _26490_, _26488_);
  not (_26578_, _26577_);
  and (_26579_, _26578_, _26491_);
  or (_26580_, _26579_, _26505_);
  or (_26581_, _26508_, _26482_);
  and (_26582_, _26581_, _26580_);
  nand (_26583_, _26582_, _26470_);
  or (_26584_, _26582_, _26470_);
  and (_26585_, _26584_, _26583_);
  not (_26586_, _26585_);
  or (_26587_, _26586_, _26576_);
  and (_26588_, _26562_, _26495_);
  not (_26589_, _26588_);
  and (_26590_, _26589_, _26583_);
  nand (_26591_, _26590_, _26587_);
  and (_26592_, _26591_, _26564_);
  nor (_26593_, _26550_, _26462_);
  nor (_26594_, _26593_, _26551_);
  not (_26595_, _26594_);
  nor (_26596_, _26554_, _26595_);
  and (_26597_, _26596_, _26592_);
  or (_26598_, _26597_, _26556_);
  nand (_26599_, _26598_, _26537_);
  nand (_26600_, _26599_, _26534_);
  and (_26601_, _26600_, _26406_);
  nand (_26602_, _26601_, _26385_);
  and (_26603_, _26602_, _26383_);
  nor (_26604_, _26602_, _26383_);
  or (_26605_, _26604_, _26603_);
  nand (_26606_, _26605_, _26379_);
  and (_26607_, _23170_, _22933_);
  nor (_26608_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_26610_, _26608_);
  and (_26611_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand (_26612_, _26608_, _23485_);
  not (_26613_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_26614_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _26613_);
  not (_26615_, _26614_);
  or (_26616_, _26615_, _23323_);
  not (_26617_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_26618_, _26617_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_26619_, _26618_);
  or (_26620_, _26619_, _23398_);
  and (_26621_, _26620_, _26616_);
  nor (_26622_, _26618_, _26614_);
  or (_26623_, _23545_, _26613_);
  nand (_26624_, _26623_, _26622_);
  nand (_26625_, _26624_, _26621_);
  and (_26626_, _26625_, _26612_);
  and (_26627_, _26626_, _23147_);
  or (_26628_, _26610_, _23518_);
  or (_26629_, _26615_, _23185_);
  or (_26630_, _26619_, _23538_);
  and (_26631_, _26630_, _26629_);
  or (_26632_, _23554_, _26613_);
  nand (_26633_, _26632_, _26622_);
  nand (_26634_, _26633_, _26631_);
  and (_26635_, _26634_, _26628_);
  and (_26636_, _26635_, _23128_);
  nand (_26637_, _26636_, _26627_);
  and (_26638_, _26635_, _23152_);
  nand (_26639_, _26634_, _26628_);
  or (_26640_, _26639_, _23220_);
  and (_26641_, _26626_, _23128_);
  and (_26642_, _26641_, _26640_);
  nand (_26643_, _26642_, _26638_);
  nand (_26644_, _26643_, _26637_);
  nand (_26645_, _26625_, _26612_);
  or (_26646_, _26645_, _23091_);
  or (_26647_, _26639_, _22976_);
  or (_26648_, _26647_, _26646_);
  nand (_26649_, _26647_, _26646_);
  and (_26650_, _26649_, _26648_);
  and (_26651_, _26650_, _26644_);
  and (_26652_, _26626_, _22977_);
  and (_26653_, _26652_, _26638_);
  or (_26654_, _26645_, _23314_);
  or (_26655_, _26654_, _26647_);
  and (_26656_, _26635_, _23313_);
  or (_26657_, _26656_, _26652_);
  and (_26658_, _26657_, _26655_);
  nand (_26659_, _26658_, _26653_);
  or (_26660_, _26658_, _26653_);
  and (_26661_, _26660_, _26659_);
  nand (_26662_, _26661_, _26651_);
  not (_26663_, _26654_);
  or (_26664_, _26655_, _23511_);
  and (_26665_, _26635_, _23949_);
  not (_26666_, _26665_);
  nand (_26667_, _26666_, _26655_);
  and (_26668_, _26667_, _26664_);
  nand (_26669_, _26668_, _26663_);
  or (_26670_, _26665_, _26663_);
  nand (_26671_, _26670_, _26669_);
  or (_26672_, _26671_, _26662_);
  or (_26673_, _26645_, _23109_);
  nor (_26674_, _26673_, _26640_);
  or (_26675_, _26636_, _26627_);
  and (_26676_, _26675_, _26637_);
  and (_26677_, _26676_, _26674_);
  or (_26678_, _26642_, _26638_);
  and (_26679_, _26678_, _26643_);
  and (_26680_, _26679_, _26677_);
  nand (_26681_, _26650_, _26644_);
  or (_26682_, _26650_, _26644_);
  and (_26683_, _26682_, _26681_);
  and (_26684_, _26683_, _26680_);
  or (_26685_, _26661_, _26651_);
  and (_26686_, _26685_, _26662_);
  nand (_26687_, _26686_, _26684_);
  not (_26688_, _26687_);
  and (_26689_, _26662_, _26659_);
  nand (_26690_, _26689_, _26671_);
  or (_26691_, _26689_, _26671_);
  and (_26692_, _26691_, _26690_);
  nand (_26693_, _26692_, _26688_);
  nand (_26694_, _26693_, _26672_);
  nor (_26695_, _26671_, _26659_);
  or (_26696_, _26639_, _23479_);
  or (_26697_, _26645_, _23511_);
  or (_26698_, _26697_, _26696_);
  nand (_26699_, _26697_, _26696_);
  and (_26700_, _26699_, _26698_);
  not (_26701_, _26700_);
  or (_26702_, _26701_, _26664_);
  or (_26703_, _26701_, _26669_);
  nand (_26704_, _26701_, _26669_);
  nand (_26705_, _26704_, _26703_);
  nand (_26706_, _26705_, _26664_);
  and (_26707_, _26706_, _26702_);
  nand (_26708_, _26707_, _26695_);
  or (_26709_, _26707_, _26695_);
  and (_26710_, _26709_, _26708_);
  nand (_26711_, _26710_, _26694_);
  or (_26712_, _26710_, _26694_);
  and (_26713_, _26712_, _26711_);
  nand (_26714_, _26713_, _26611_);
  or (_26715_, _26713_, _26611_);
  nand (_26716_, _26715_, _26714_);
  and (_26717_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_26718_, _26692_, _26688_);
  and (_26719_, _26718_, _26693_);
  nand (_26720_, _26719_, _26717_);
  or (_26721_, _26719_, _26717_);
  nand (_26722_, _26721_, _26720_);
  and (_26723_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or (_26724_, _26686_, _26684_);
  and (_26725_, _26724_, _26687_);
  nand (_26726_, _26725_, _26723_);
  or (_26727_, _26725_, _26723_);
  and (_26728_, _26727_, _26726_);
  and (_26729_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nand (_26730_, _26683_, _26680_);
  or (_26731_, _26683_, _26680_);
  and (_26732_, _26731_, _26730_);
  nand (_26733_, _26732_, _26729_);
  and (_26734_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nand (_26735_, _26679_, _26677_);
  or (_26736_, _26679_, _26677_);
  and (_26737_, _26736_, _26735_);
  nand (_26738_, _26737_, _26734_);
  and (_26739_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_26740_, _26676_, _26674_);
  or (_26741_, _26676_, _26674_);
  and (_26742_, _26741_, _26740_);
  and (_26743_, _26742_, _26739_);
  not (_26744_, _26743_);
  or (_26745_, _26737_, _26734_);
  nand (_26746_, _26745_, _26738_);
  or (_26747_, _26746_, _26744_);
  nand (_26748_, _26747_, _26738_);
  or (_26749_, _26732_, _26729_);
  and (_26750_, _26749_, _26733_);
  nand (_26751_, _26750_, _26748_);
  nand (_26752_, _26751_, _26733_);
  nand (_26753_, _26752_, _26728_);
  and (_26754_, _26753_, _26726_);
  or (_26755_, _26754_, _26722_);
  and (_26756_, _26755_, _26720_);
  or (_26757_, _26756_, _26716_);
  nand (_26758_, _26757_, _26714_);
  and (_26759_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  nand (_26761_, _26711_, _26708_);
  and (_26762_, _26626_, _23636_);
  and (_26763_, _26762_, _26666_);
  and (_26764_, _26702_, _26703_);
  not (_26765_, _26764_);
  nand (_26766_, _26765_, _26763_);
  or (_26767_, _26765_, _26763_);
  and (_26768_, _26767_, _26766_);
  nand (_26769_, _26768_, _26761_);
  or (_26770_, _26768_, _26761_);
  and (_26771_, _26770_, _26769_);
  nand (_26772_, _26771_, _26759_);
  or (_26773_, _26771_, _26759_);
  and (_26774_, _26773_, _26772_);
  and (_26775_, _26774_, _26758_);
  nor (_26776_, _26774_, _26758_);
  nor (_26777_, _26776_, _26775_);
  and (_26778_, _26777_, _26607_);
  and (_26779_, _23636_, _23670_);
  nor (_26780_, _23639_, _23173_);
  nor (_26781_, _26780_, _23109_);
  nor (_26782_, _26781_, _26779_);
  and (_26783_, _26782_, _24036_);
  and (_26784_, _23635_, _23048_);
  nand (_26785_, _23176_, _23147_);
  nand (_26786_, _24042_, _26785_);
  nor (_26787_, _26786_, _26784_);
  and (_26788_, _26787_, _26783_);
  nor (_26789_, _23597_, _23458_);
  not (_26790_, _26789_);
  and (_26792_, _26790_, _26190_);
  not (_26793_, _26792_);
  and (_26794_, _26793_, _24039_);
  and (_26795_, _26794_, _26788_);
  not (_26796_, _26795_);
  nor (_26797_, _26796_, _26778_);
  nand (_26798_, _26797_, _26606_);
  and (_26799_, _24733_, _26253_);
  nor (_26800_, _26799_, _26169_);
  and (_26801_, _26166_, _24646_);
  not (_26802_, _26801_);
  and (_26803_, _25851_, _24646_);
  nor (_26804_, _26803_, _24643_);
  and (_26805_, _26804_, _26802_);
  and (_26806_, _26230_, _25852_);
  nand (_26807_, _26806_, _26239_);
  nand (_26808_, _26807_, _24733_);
  nand (_26809_, _26808_, _26805_);
  not (_26810_, _24733_);
  not (_26811_, _25852_);
  nor (_00002_, _26811_, _26253_);
  nor (_00003_, _26254_, _25863_);
  and (_00004_, _00003_, _26239_);
  and (_00005_, _00004_, _00002_);
  and (_00006_, _00005_, _26236_);
  nor (_00007_, _00006_, _26810_);
  nor (_00008_, _00007_, _26809_);
  and (_00009_, _00008_, _26800_);
  or (_00010_, _00009_, _26799_);
  and (_00011_, _00010_, _26798_);
  and (_00012_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_00013_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_00014_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00015_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_00016_, _00015_, _00014_);
  and (_00017_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00018_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_00019_, _00018_, _00017_);
  and (_00020_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00021_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_00022_, _00021_, _00020_);
  and (_00023_, _00022_, _00019_);
  and (_00024_, _00023_, _00016_);
  nor (_00025_, _00024_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_00026_, _00025_, _00013_);
  nor (_00027_, _00026_, _24883_);
  nor (_00028_, _00027_, _00012_);
  and (_00029_, _00028_, _26809_);
  and (_00030_, _26808_, _26805_);
  and (_00031_, _00030_, _26340_);
  nor (_00034_, _00031_, _00029_);
  and (_00035_, _00034_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_00036_, _00034_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00037_, _00007_, _26803_);
  not (_00038_, _26800_);
  and (_00039_, _00030_, _00038_);
  nor (_00040_, _00039_, _00037_);
  nand (_00041_, _00040_, _00036_);
  nor (_00042_, _00041_, _00035_);
  nor (_00043_, _00028_, _26802_);
  and (_00044_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00045_, _00008_, _00038_);
  and (_00046_, _00045_, _26341_);
  or (_00047_, _00046_, _00044_);
  or (_00048_, _00047_, _00043_);
  or (_00049_, _00048_, _00042_);
  or (_00050_, _00049_, _00011_);
  and (_00051_, _00050_, _26378_);
  not (_00052_, _26378_);
  and (_00053_, _00052_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00054_, _00053_, _00051_);
  and (_26861_[0], _00054_, _22773_);
  nand (_00055_, _26600_, _26406_);
  or (_00056_, _26574_, _26572_);
  and (_00057_, _00056_, _26575_);
  or (_00058_, _00057_, _00055_);
  or (_00059_, _26601_, _26569_);
  and (_00060_, _00059_, _00058_);
  nand (_00061_, _00060_, _26379_);
  not (_00062_, _26772_);
  nor (_00063_, _26775_, _00062_);
  and (_00064_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and (_00065_, _26766_, _26698_);
  nand (_00066_, _00065_, _26769_);
  nand (_00067_, _00066_, _00064_);
  or (_00068_, _00066_, _00064_);
  nand (_00069_, _00068_, _00067_);
  or (_00070_, _00069_, _00063_);
  nand (_00071_, _00069_, _00063_);
  and (_00072_, _00071_, _00070_);
  nand (_00073_, _00072_, _26607_);
  nor (_00074_, _23571_, _23548_);
  or (_00075_, _00074_, _23601_);
  and (_00076_, _00075_, _23608_);
  nor (_00077_, _00075_, _23608_);
  or (_00078_, _00077_, _00076_);
  and (_00079_, _00078_, _23597_);
  nor (_00080_, _23579_, _23576_);
  nor (_00081_, _00080_, _23580_);
  nor (_00082_, _00081_, _23459_);
  nor (_00083_, _00082_, _00079_);
  not (_00084_, _23639_);
  nor (_00085_, _23640_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_00086_, _00085_, _23147_);
  nor (_00087_, _00085_, _23147_);
  nor (_00088_, _00087_, _00086_);
  nor (_00089_, _00088_, _00084_);
  not (_00090_, _00089_);
  nand (_00091_, _23176_, _23128_);
  and (_00092_, _23173_, _23147_);
  and (_00093_, _23179_, _23153_);
  nor (_00094_, _00093_, _00092_);
  and (_00095_, _00094_, _00091_);
  and (_00096_, _00095_, _23742_);
  and (_00097_, _00096_, _00090_);
  and (_00098_, _00097_, _23734_);
  and (_00099_, _00098_, _00083_);
  and (_00100_, _00099_, _00073_);
  nand (_00101_, _00100_, _00061_);
  and (_00102_, _00101_, _00010_);
  and (_00103_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_00104_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_00106_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00107_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00108_, _00107_, _00106_);
  and (_00109_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00110_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_00111_, _00110_, _00109_);
  or (_00112_, _00111_, _00108_);
  and (_00113_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00114_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00115_, _00114_, _00113_);
  or (_00116_, _00115_, _00112_);
  and (_00117_, _00116_, _24568_);
  or (_00118_, _00117_, _00104_);
  and (_00119_, _00118_, _23760_);
  nor (_00120_, _00119_, _00103_);
  or (_00121_, _00120_, _00030_);
  or (_00122_, _26809_, _25427_);
  and (_00123_, _00122_, _00121_);
  or (_00124_, _00123_, _23129_);
  nand (_00126_, _00123_, _23129_);
  and (_00127_, _00126_, _00124_);
  or (_00128_, _00127_, _00035_);
  and (_00129_, _00127_, _00035_);
  not (_00130_, _00129_);
  and (_00131_, _00130_, _00040_);
  and (_00132_, _00131_, _00128_);
  and (_00133_, _00045_, _26308_);
  nor (_00134_, _00120_, _26802_);
  and (_00135_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00136_, _00135_, _00134_);
  or (_00137_, _00136_, _00133_);
  or (_00138_, _00137_, _00132_);
  nor (_00139_, _00138_, _00102_);
  nand (_00140_, _00139_, _26378_);
  or (_00141_, _26378_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00143_, _00141_, _22773_);
  and (_26861_[1], _00143_, _00140_);
  not (_00144_, _26587_);
  and (_00145_, _26586_, _26576_);
  nor (_00146_, _00145_, _00144_);
  or (_00147_, _00146_, _00055_);
  or (_00148_, _26601_, _26582_);
  and (_00149_, _00148_, _00147_);
  nand (_00150_, _00149_, _26379_);
  and (_00151_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  nand (_00152_, _00070_, _00067_);
  nand (_00153_, _00152_, _00151_);
  or (_00154_, _00152_, _00151_);
  and (_00155_, _00154_, _00153_);
  nand (_00156_, _00155_, _26607_);
  nor (_00157_, _23580_, _23569_);
  nor (_00158_, _00157_, _23581_);
  nor (_00159_, _00158_, _23459_);
  and (_00160_, _23179_, _23147_);
  not (_00161_, _00160_);
  and (_00162_, _23173_, _23128_);
  not (_00163_, _00162_);
  not (_00165_, _23176_);
  or (_00166_, _00165_, _23091_);
  and (_00167_, _00166_, _00163_);
  and (_00168_, _00167_, _00161_);
  and (_00169_, _00168_, _23245_);
  not (_00170_, _00169_);
  nor (_00171_, _00170_, _00159_);
  nor (_00172_, _23612_, _23610_);
  nor (_00173_, _00172_, _23598_);
  and (_00174_, _00173_, _23614_);
  and (_00175_, _23148_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00176_, _00087_, _23241_);
  nor (_00177_, _00176_, _00175_);
  nor (_00178_, _00177_, _00084_);
  nor (_00179_, _00178_, _00174_);
  and (_00180_, _00179_, _00171_);
  and (_00181_, _00180_, _23229_);
  and (_00182_, _00181_, _00156_);
  nand (_00183_, _00182_, _00150_);
  and (_00184_, _00183_, _00010_);
  nand (_00185_, _00130_, _00124_);
  and (_00186_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_00187_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_00188_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00189_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00190_, _00189_, _00188_);
  and (_00191_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00192_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_00193_, _00192_, _00191_);
  or (_00194_, _00193_, _00190_);
  and (_00195_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00196_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00197_, _00196_, _00195_);
  or (_00198_, _00197_, _00194_);
  and (_00199_, _00198_, _24568_);
  or (_00200_, _00199_, _00187_);
  and (_00201_, _00200_, _23760_);
  nor (_00202_, _00201_, _00186_);
  nor (_00203_, _00202_, _00030_);
  and (_00204_, _00030_, _26361_);
  nor (_00205_, _00204_, _00203_);
  nor (_00206_, _00205_, _23114_);
  and (_00207_, _00205_, _23114_);
  nor (_00208_, _00207_, _00206_);
  and (_00209_, _00208_, _00185_);
  or (_00210_, _00208_, _00185_);
  nand (_00211_, _00210_, _00040_);
  nor (_00212_, _00211_, _00209_);
  and (_00213_, _00203_, _26169_);
  and (_00214_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_00215_, _00045_, _26361_);
  or (_00216_, _00215_, _00214_);
  or (_00217_, _00216_, _00213_);
  or (_00218_, _00217_, _00212_);
  or (_00219_, _00218_, _00184_);
  and (_00220_, _00219_, _26378_);
  not (_00221_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00222_, _25524_, _00221_);
  and (_00223_, _25524_, _00221_);
  nor (_00224_, _00223_, _00222_);
  and (_00225_, _00224_, _00052_);
  or (_00226_, _00225_, _00220_);
  and (_26861_[2], _00226_, _22773_);
  not (_00227_, _26562_);
  or (_00228_, _26601_, _00227_);
  or (_00229_, _26588_, _26563_);
  and (_00230_, _26587_, _26583_);
  and (_00231_, _00230_, _00229_);
  nor (_00232_, _00230_, _00229_);
  or (_00233_, _00232_, _00231_);
  or (_00234_, _00233_, _00055_);
  nand (_00235_, _00234_, _00228_);
  nand (_00236_, _00235_, _26379_);
  or (_00237_, _00069_, _26772_);
  nand (_00238_, _00237_, _00067_);
  and (_00239_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_00240_, _00239_, _00151_);
  and (_00241_, _00240_, _00238_);
  and (_00242_, _00068_, _00067_);
  and (_00243_, _00242_, _26774_);
  and (_00244_, _00240_, _00243_);
  and (_00245_, _00244_, _26758_);
  or (_00246_, _00245_, _00241_);
  not (_00247_, _00246_);
  not (_00248_, _00239_);
  nand (_00249_, _00248_, _00153_);
  and (_00250_, _00249_, _00247_);
  nand (_00251_, _00250_, _26607_);
  and (_00252_, _23614_, _23607_);
  or (_00253_, _00252_, _23598_);
  nor (_00254_, _00253_, _23615_);
  not (_00255_, _00254_);
  nor (_00256_, _26188_, _23459_);
  not (_00257_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00258_, _23148_, _00257_);
  nor (_00259_, _00258_, _23152_);
  and (_00260_, _23173_, _23152_);
  not (_00261_, _00260_);
  or (_00262_, _23640_, _00084_);
  and (_00263_, _00262_, _00261_);
  or (_00264_, _00263_, _00259_);
  not (_00265_, _23409_);
  and (_00266_, _23402_, _00265_);
  or (_00267_, _00165_, _22976_);
  and (_00268_, _23179_, _23128_);
  not (_00269_, _00268_);
  and (_00270_, _00269_, _00267_);
  and (_00271_, _00270_, _00266_);
  and (_00272_, _00271_, _00264_);
  nand (_00273_, _00272_, _23397_);
  nor (_00274_, _00273_, _00256_);
  and (_00275_, _00274_, _00255_);
  and (_00276_, _00275_, _00251_);
  nand (_00277_, _00276_, _00236_);
  and (_00278_, _00277_, _00010_);
  or (_00279_, _00209_, _00206_);
  and (_00280_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_00281_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_00282_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00283_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_00284_, _00283_, _00282_);
  and (_00285_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00286_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_00287_, _00286_, _00285_);
  and (_00288_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00289_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_00290_, _00289_, _00288_);
  and (_00291_, _00290_, _00287_);
  and (_00292_, _00291_, _00284_);
  nor (_00293_, _00292_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_00294_, _00293_, _00281_);
  nor (_00295_, _00294_, _24883_);
  nor (_00296_, _00295_, _00280_);
  nor (_00297_, _00296_, _00030_);
  and (_00298_, _00030_, _26072_);
  nor (_00299_, _00298_, _00297_);
  nor (_00300_, _00299_, _23071_);
  and (_00301_, _00299_, _23071_);
  nor (_00302_, _00301_, _00300_);
  or (_00303_, _00302_, _00279_);
  nand (_00304_, _00302_, _00279_);
  and (_00305_, _00304_, _00040_);
  and (_00306_, _00305_, _00303_);
  and (_00307_, _00297_, _26169_);
  and (_00308_, _00045_, _26072_);
  and (_00309_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_00310_, _00309_, _00308_);
  or (_00311_, _00310_, _00307_);
  or (_00312_, _00311_, _00306_);
  nor (_00313_, _00312_, _00278_);
  nand (_00314_, _00313_, _26378_);
  and (_00315_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not (_00316_, _00315_);
  nor (_00317_, _00316_, _25524_);
  nor (_00318_, _00222_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00319_, _00318_, _00317_);
  or (_00320_, _00319_, _26378_);
  and (_00321_, _00320_, _22773_);
  and (_26861_[3], _00321_, _00314_);
  nand (_00322_, _26594_, _26592_);
  or (_00323_, _26594_, _26592_);
  and (_00324_, _00323_, _00322_);
  or (_00325_, _00324_, _00055_);
  or (_00326_, _26601_, _26550_);
  and (_00327_, _00326_, _00325_);
  and (_00328_, _00327_, _26379_);
  and (_00329_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_00330_, _00329_, _00246_);
  nor (_00331_, _00329_, _00246_);
  nor (_00332_, _00331_, _00330_);
  and (_00333_, _00332_, _26607_);
  and (_00334_, _26172_, _23458_);
  or (_00335_, _23618_, _23188_);
  nor (_00336_, _23620_, _23598_);
  and (_00337_, _00336_, _00335_);
  or (_00338_, _23641_, _22977_);
  nor (_00339_, _23653_, _00084_);
  and (_00340_, _00339_, _00338_);
  and (_00341_, _23173_, _22977_);
  and (_00342_, _23313_, _23176_);
  and (_00343_, _23179_, _23152_);
  or (_00344_, _00343_, _00342_);
  nor (_00345_, _00344_, _00341_);
  nand (_00346_, _00345_, _23202_);
  nor (_00347_, _00346_, _00340_);
  nand (_00348_, _00347_, _23163_);
  or (_00349_, _00348_, _00337_);
  or (_00350_, _00349_, _00334_);
  or (_00351_, _00350_, _00333_);
  or (_00352_, _00351_, _00328_);
  and (_00353_, _00352_, _00010_);
  and (_00354_, _00030_, _26005_);
  and (_00355_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_00356_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_00357_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00358_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00359_, _00358_, _00357_);
  and (_00360_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00361_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_00362_, _00361_, _00360_);
  or (_00363_, _00362_, _00359_);
  and (_00365_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00366_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00367_, _00366_, _00365_);
  or (_00368_, _00367_, _00363_);
  and (_00369_, _00368_, _24568_);
  or (_00370_, _00369_, _00356_);
  and (_00371_, _00370_, _23760_);
  nor (_00372_, _00371_, _00355_);
  not (_00373_, _00372_);
  and (_00374_, _00373_, _26809_);
  nor (_00376_, _00374_, _00354_);
  or (_00377_, _00376_, _22939_);
  nand (_00378_, _00376_, _22939_);
  and (_00380_, _00378_, _00377_);
  nor (_00381_, _00300_, _00279_);
  nor (_00382_, _00381_, _00301_);
  nand (_00383_, _00382_, _00380_);
  or (_00384_, _00382_, _00380_);
  and (_00385_, _00384_, _00040_);
  and (_00386_, _00385_, _00383_);
  and (_00387_, _00045_, _26005_);
  and (_00388_, _00373_, _26801_);
  and (_00389_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00390_, _00389_, _00388_);
  or (_00391_, _00390_, _00387_);
  nor (_00392_, _00391_, _00386_);
  nand (_00393_, _00392_, _26378_);
  or (_00394_, _00393_, _00353_);
  and (_00395_, _00317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00396_, _00317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00397_, _00396_, _00395_);
  or (_00398_, _00397_, _26378_);
  and (_00399_, _00398_, _22773_);
  and (_26861_[4], _00399_, _00394_);
  and (_00400_, _00055_, _26544_);
  nand (_00401_, _00322_, _26552_);
  nor (_00402_, _00401_, _26554_);
  and (_00403_, _00401_, _26554_);
  or (_00404_, _00403_, _00402_);
  and (_00405_, _00404_, _26601_);
  or (_00406_, _00405_, _00400_);
  and (_00407_, _00406_, _26379_);
  and (_00408_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_00409_, _00408_, _00329_);
  nand (_00410_, _00409_, _00246_);
  or (_00411_, _00408_, _00330_);
  and (_00412_, _00411_, _00410_);
  and (_00413_, _00412_, _26607_);
  nor (_00414_, _26186_, _23459_);
  nor (_00415_, _23346_, _23186_);
  nor (_00416_, _00415_, _23623_);
  or (_00417_, _00416_, _23620_);
  nor (_00419_, _23621_, _23598_);
  and (_00420_, _00419_, _00417_);
  nor (_00422_, _23945_, _23479_);
  nor (_00423_, _00422_, _23641_);
  and (_00424_, _00423_, _23046_);
  and (_00425_, _00424_, _23639_);
  or (_00426_, _00425_, _23173_);
  and (_00427_, _00426_, _23313_);
  and (_00428_, _23179_, _22977_);
  nor (_00429_, _23511_, _00165_);
  nor (_00430_, _00429_, _00428_);
  nand (_00431_, _00430_, _23355_);
  and (_00432_, _23653_, _23313_);
  nor (_00433_, _00432_, _23654_);
  or (_00434_, _00424_, _00084_);
  nor (_00435_, _00434_, _00433_);
  or (_00436_, _00435_, _00431_);
  nor (_00438_, _00436_, _00427_);
  nand (_00439_, _00438_, _23340_);
  or (_00440_, _00439_, _00420_);
  or (_00441_, _00440_, _00414_);
  or (_00442_, _00441_, _00413_);
  or (_00443_, _00442_, _00407_);
  and (_00444_, _00443_, _00010_);
  nand (_00446_, _00383_, _00377_);
  and (_00447_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_00448_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_00449_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00450_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_00451_, _00450_, _00449_);
  and (_00452_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00453_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_00454_, _00453_, _00452_);
  and (_00455_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00456_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_00457_, _00456_, _00455_);
  and (_00458_, _00457_, _00454_);
  and (_00459_, _00458_, _00451_);
  nor (_00460_, _00459_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_00461_, _00460_, _00448_);
  nor (_00462_, _00461_, _24883_);
  nor (_00463_, _00462_, _00447_);
  not (_00464_, _00463_);
  and (_00465_, _00464_, _26809_);
  and (_00466_, _00030_, _26019_);
  nor (_00467_, _00466_, _00465_);
  nor (_00468_, _00467_, _23296_);
  and (_00469_, _00467_, _23296_);
  nor (_00470_, _00469_, _00468_);
  or (_00471_, _00470_, _00446_);
  and (_00472_, _00470_, _00446_);
  not (_00473_, _00472_);
  and (_00474_, _00473_, _00040_);
  and (_00475_, _00474_, _00471_);
  and (_00476_, _00045_, _26019_);
  and (_00477_, _00464_, _26801_);
  and (_00478_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00479_, _00478_, _00477_);
  or (_00480_, _00479_, _00476_);
  nor (_00481_, _00480_, _00475_);
  nand (_00482_, _00481_, _26378_);
  or (_00483_, _00482_, _00444_);
  and (_00484_, _00395_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00485_, _00395_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00486_, _00485_, _00484_);
  or (_00487_, _00486_, _26378_);
  and (_00488_, _00487_, _22773_);
  and (_26861_[5], _00488_, _00483_);
  or (_00489_, _00472_, _00468_);
  and (_00491_, _24883_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_00492_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_00493_, _24478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00494_, _24474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00495_, _00494_, _00493_);
  and (_00496_, _24486_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00497_, _24481_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_00498_, _00497_, _00496_);
  or (_00499_, _00498_, _00495_);
  and (_00500_, _24470_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00501_, _24484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00502_, _00501_, _00500_);
  or (_00503_, _00502_, _00499_);
  and (_00504_, _00503_, _24568_);
  or (_00505_, _00504_, _00492_);
  and (_00506_, _00505_, _23760_);
  nor (_00507_, _00506_, _00491_);
  and (_00508_, _00507_, _26809_);
  and (_00509_, _00030_, _26107_);
  nor (_00511_, _00509_, _00508_);
  nand (_00512_, _00511_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_00513_, _00511_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00514_, _00513_, _00512_);
  nand (_00515_, _00514_, _00489_);
  or (_00517_, _00514_, _00489_);
  and (_00518_, _00517_, _00515_);
  and (_00519_, _00518_, _00040_);
  nand (_00521_, _26598_, _26536_);
  or (_00522_, _26598_, _26536_);
  nand (_00523_, _00522_, _00521_);
  nand (_00524_, _00523_, _26601_);
  or (_00526_, _26601_, _26527_);
  and (_00527_, _00526_, _00524_);
  nand (_00528_, _00527_, _26379_);
  and (_00529_, _00409_, _00246_);
  and (_00530_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  nand (_00531_, _00530_, _00529_);
  or (_00532_, _00530_, _00529_);
  and (_00533_, _00532_, _00531_);
  nand (_00534_, _00533_, _26607_);
  nor (_00535_, _23627_, _23621_);
  nor (_00536_, _00535_, _23628_);
  and (_00538_, _00536_, _23597_);
  not (_00539_, _00538_);
  nor (_00540_, _26176_, _23459_);
  and (_00541_, _23313_, _23179_);
  not (_00542_, _00541_);
  or (_00543_, _23479_, _00165_);
  and (_00544_, _00543_, _00542_);
  and (_00545_, _23949_, _23173_);
  not (_00546_, _00545_);
  and (_00547_, _00546_, _24010_);
  nand (_00548_, _00547_, _00544_);
  not (_00549_, _23654_);
  nor (_00550_, _00424_, _00549_);
  and (_00551_, _00550_, _23949_);
  not (_00552_, _00551_);
  nor (_00553_, _00550_, _23949_);
  nor (_00554_, _00553_, _00084_);
  and (_00555_, _00554_, _00552_);
  not (_00556_, _00555_);
  nand (_00557_, _00556_, _24006_);
  or (_00558_, _00557_, _00548_);
  nor (_00559_, _00558_, _24014_);
  not (_00560_, _00559_);
  nor (_00561_, _00560_, _00540_);
  and (_00562_, _00561_, _00539_);
  and (_00563_, _00562_, _00534_);
  nand (_00564_, _00563_, _00528_);
  and (_00566_, _00564_, _00010_);
  nor (_00567_, _00507_, _26802_);
  and (_00568_, _00045_, _26108_);
  and (_00569_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00570_, _00569_, _00568_);
  or (_00571_, _00570_, _00567_);
  or (_00572_, _00571_, _00566_);
  nor (_00573_, _00572_, _00519_);
  nand (_00574_, _00573_, _26378_);
  and (_00575_, _00484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00576_, _00484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00577_, _00576_, _00575_);
  or (_00578_, _00577_, _26378_);
  and (_00579_, _00578_, _22773_);
  and (_26861_[6], _00579_, _00574_);
  or (_00580_, _26601_, _26529_);
  nand (_00581_, _00521_, _26528_);
  nand (_00582_, _00581_, _26532_);
  nand (_00583_, _00582_, _26601_);
  and (_00584_, _00583_, _00580_);
  nand (_00585_, _00584_, _26379_);
  and (_00586_, _26610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_00587_, _00586_, _00531_);
  or (_00588_, _00531_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_00589_, _00588_, _00587_);
  nand (_00590_, _00589_, _26607_);
  and (_00591_, _26182_, _23458_);
  not (_00592_, _00591_);
  nor (_00593_, _23631_, _26178_);
  and (_00594_, _23631_, _26178_);
  or (_00595_, _00594_, _00593_);
  nor (_00596_, _00595_, _23598_);
  and (_00597_, _23642_, _23048_);
  and (_00598_, _23636_, _23173_);
  and (_00599_, _23949_, _23179_);
  or (_00600_, _00599_, _00598_);
  and (_00601_, _23663_, _23153_);
  not (_00602_, _00601_);
  nand (_00603_, _00602_, _23969_);
  or (_00604_, _00603_, _00600_);
  or (_00605_, _00604_, _00597_);
  nor (_00606_, _00424_, _23655_);
  nor (_00607_, _00606_, _23479_);
  and (_00608_, _00606_, _23479_);
  nor (_00609_, _00608_, _00607_);
  nor (_00610_, _00609_, _00084_);
  not (_00611_, _00610_);
  nand (_00612_, _00611_, _23966_);
  or (_00613_, _00612_, _00605_);
  nor (_00614_, _00613_, _23973_);
  not (_00615_, _00614_);
  nor (_00616_, _00615_, _00596_);
  and (_00617_, _00616_, _00592_);
  and (_00618_, _00617_, _00590_);
  nand (_00619_, _00618_, _00585_);
  and (_00620_, _00619_, _00010_);
  nand (_00621_, _00515_, _00512_);
  nor (_00622_, _00030_, _24900_);
  and (_00623_, _00030_, _26149_);
  nor (_00624_, _00623_, _00622_);
  nor (_00625_, _00624_, _23460_);
  and (_00626_, _00624_, _23460_);
  nor (_00627_, _00626_, _00625_);
  nand (_00628_, _00627_, _00621_);
  or (_00630_, _00627_, _00621_);
  and (_00631_, _00630_, _00040_);
  and (_00632_, _00631_, _00628_);
  and (_00633_, _00045_, _26149_);
  nor (_00634_, _26802_, _24900_);
  and (_00635_, _24643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_00636_, _00635_, _00634_);
  or (_00637_, _00636_, _00633_);
  nor (_00638_, _00637_, _00632_);
  nand (_00639_, _00638_, _26378_);
  or (_00640_, _00639_, _00620_);
  nor (_00641_, _00575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_00643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_00644_, _00643_, _00642_);
  and (_00645_, _00644_, _00315_);
  not (_00646_, _00645_);
  nor (_00647_, _00646_, _25524_);
  nor (_00648_, _00647_, _00641_);
  or (_00649_, _00648_, _26378_);
  and (_00650_, _00649_, _22773_);
  and (_26861_[7], _00650_, _00640_);
  not (_00651_, _00624_);
  not (_00652_, _00626_);
  and (_00653_, _00652_, _00621_);
  or (_00654_, _00653_, _00625_);
  and (_00655_, _00654_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00656_, _00654_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00657_, _00656_, _00655_);
  or (_00658_, _00657_, _00651_);
  nand (_00659_, _00657_, _00651_);
  and (_00660_, _00659_, _00658_);
  and (_00661_, _00660_, _00040_);
  and (_00662_, _26798_, _24643_);
  and (_00663_, _26801_, _26341_);
  nor (_00664_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_00665_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00666_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _00665_);
  nor (_00667_, _00666_, _00664_);
  not (_00668_, _00667_);
  or (_00669_, _00668_, _23633_);
  and (_00670_, _00668_, _23633_);
  nor (_00671_, _00670_, _23598_);
  and (_00672_, _00671_, _00669_);
  nand (_00673_, _26601_, _26379_);
  nor (_00674_, _23963_, _23658_);
  and (_00675_, _00674_, _23953_);
  nor (_00676_, _00675_, _23554_);
  and (_00677_, _00675_, _23554_);
  or (_00678_, _00677_, _23335_);
  nor (_00679_, _00678_, _00676_);
  and (_00680_, _23554_, _23173_);
  and (_00681_, _26635_, _23153_);
  and (_00682_, _00681_, _26607_);
  and (_00683_, _23635_, _22977_);
  nor (_00684_, _23109_, _23316_);
  or (_00685_, _00684_, _00683_);
  or (_00686_, _00685_, _00682_);
  nor (_00687_, _00686_, _00680_);
  not (_00688_, _00687_);
  nor (_00689_, _00688_, _00679_);
  nand (_00690_, _00689_, _00673_);
  or (_00691_, _00690_, _00672_);
  and (_00692_, _00691_, _26799_);
  not (_00693_, _24495_);
  and (_00694_, _00045_, _00693_);
  and (_00695_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00696_, _00695_, _00694_);
  or (_00697_, _00696_, _00692_);
  or (_00698_, _00697_, _00663_);
  or (_00699_, _00698_, _00662_);
  or (_00700_, _00699_, _00661_);
  or (_00701_, _00700_, _00052_);
  and (_00702_, _00647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00703_, _00647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00704_, _00703_, _00702_);
  or (_00706_, _00704_, _26378_);
  and (_00707_, _00706_, _22773_);
  and (_26861_[8], _00707_, _00701_);
  and (_00708_, _00101_, _24643_);
  not (_00709_, _26799_);
  nor (_00710_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_00711_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00712_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _00711_);
  nor (_00713_, _00712_, _00710_);
  not (_00714_, _00713_);
  and (_00715_, _00714_, _00669_);
  not (_00716_, _00715_);
  or (_00717_, _00714_, _00669_);
  and (_00718_, _00717_, _23597_);
  and (_00719_, _00718_, _00716_);
  not (_00720_, _00719_);
  and (_00721_, _26508_, _26379_);
  not (_00722_, _00721_);
  nor (_00723_, _23570_, _23479_);
  and (_00724_, _00723_, _23951_);
  nand (_00725_, _00724_, _23046_);
  and (_00726_, _23570_, _23479_);
  and (_00727_, _00726_, _23946_);
  nand (_00728_, _00727_, _23048_);
  and (_00729_, _00728_, _00725_);
  nor (_00730_, _00729_, _23545_);
  and (_00731_, _00729_, _23545_);
  or (_00733_, _00731_, _00730_);
  and (_00734_, _00733_, _23067_);
  and (_00735_, _23545_, _23173_);
  and (_00736_, _26673_, _26640_);
  nor (_00737_, _00736_, _26674_);
  and (_00738_, _00737_, _26607_);
  and (_00739_, _23313_, _23635_);
  and (_00740_, _23147_, _22938_);
  or (_00741_, _00740_, _00739_);
  or (_00742_, _00741_, _00738_);
  nor (_00743_, _00742_, _00735_);
  not (_00744_, _00743_);
  nor (_00745_, _00744_, _00734_);
  and (_00746_, _00745_, _00722_);
  and (_00747_, _00746_, _00720_);
  nor (_00748_, _00747_, _00709_);
  and (_00749_, _26801_, _26308_);
  not (_00750_, _24537_);
  and (_00751_, _00045_, _00750_);
  and (_00752_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_00753_, _00752_, _00751_);
  or (_00754_, _00753_, _00749_);
  or (_00755_, _00754_, _00748_);
  nor (_00756_, _00755_, _00708_);
  nand (_00757_, _00756_, _26378_);
  and (_00758_, _00655_, _00624_);
  and (_00759_, _00656_, _00651_);
  nor (_00760_, _00759_, _00758_);
  nand (_00761_, _00760_, _00711_);
  or (_00762_, _00760_, _00711_);
  and (_00763_, _00762_, _00761_);
  and (_00764_, _00763_, _00040_);
  or (_00765_, _00764_, _00757_);
  and (_00766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00767_, _00766_, _00647_);
  nor (_00768_, _00702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00769_, _00768_, _00767_);
  or (_00770_, _00769_, _26378_);
  and (_00771_, _00770_, _22773_);
  and (_26861_[9], _00771_, _00765_);
  not (_00772_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00773_, _00759_, _00711_);
  and (_00774_, _00655_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00775_, _00774_, _00624_);
  nor (_00776_, _00775_, _00773_);
  nand (_00777_, _00776_, _00772_);
  or (_00778_, _00776_, _00772_);
  and (_00780_, _00778_, _00040_);
  and (_00781_, _00780_, _00777_);
  and (_00782_, _00183_, _24643_);
  nor (_00783_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00784_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _00772_);
  nor (_00785_, _00784_, _00783_);
  not (_00786_, _00785_);
  and (_00787_, _00786_, _00717_);
  not (_00788_, _00787_);
  or (_00789_, _00786_, _00717_);
  and (_00790_, _00789_, _23597_);
  and (_00791_, _00790_, _00788_);
  not (_00792_, _00791_);
  nor (_00793_, _26742_, _26739_);
  nor (_00794_, _00793_, _26743_);
  and (_00795_, _00794_, _26607_);
  and (_00796_, _23949_, _23635_);
  and (_00797_, _23217_, _23173_);
  or (_00798_, _00797_, _00796_);
  nor (_00799_, _00798_, _00795_);
  and (_00800_, _00727_, _23558_);
  and (_00801_, _00800_, _23048_);
  and (_00802_, _00724_, _23545_);
  and (_00803_, _00802_, _23046_);
  nor (_00804_, _00803_, _00801_);
  nor (_00805_, _00804_, _23538_);
  not (_00806_, _00805_);
  and (_00807_, _00804_, _23538_);
  nor (_00808_, _00807_, _23335_);
  and (_00809_, _00808_, _00806_);
  and (_00810_, _23128_, _22938_);
  and (_00811_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_00812_, _00811_, _00810_);
  nor (_00813_, _00812_, _00809_);
  and (_00814_, _00813_, _00799_);
  and (_00815_, _00814_, _00792_);
  nor (_00816_, _00815_, _00709_);
  and (_00817_, _26801_, _26361_);
  not (_00818_, _24518_);
  and (_00819_, _00045_, _00818_);
  and (_00820_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_00821_, _00820_, _00819_);
  or (_00822_, _00821_, _00817_);
  nor (_00823_, _00822_, _00816_);
  nand (_00824_, _00823_, _26378_);
  or (_00825_, _00824_, _00782_);
  or (_00826_, _00825_, _00781_);
  nor (_00827_, _00767_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00828_, _00766_, _00645_);
  and (_00829_, _00828_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00830_, _00829_, _25591_);
  nor (_00831_, _00830_, _00827_);
  or (_00832_, _00831_, _26378_);
  and (_00833_, _00832_, _22773_);
  and (_26861_[10], _00833_, _00826_);
  not (_00834_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00835_, _00656_, _00711_);
  and (_00836_, _00835_, _00772_);
  and (_00837_, _00836_, _00651_);
  and (_00838_, _00774_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00839_, _00838_, _00624_);
  nor (_00840_, _00839_, _00837_);
  nand (_00841_, _00840_, _00834_);
  or (_00842_, _00840_, _00834_);
  and (_00843_, _00842_, _00040_);
  and (_00844_, _00843_, _00841_);
  and (_00845_, _00277_, _24643_);
  nor (_00846_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00847_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _00834_);
  nor (_00848_, _00847_, _00846_);
  not (_00849_, _00848_);
  and (_00850_, _00849_, _00789_);
  nor (_00851_, _00849_, _00789_);
  nor (_00852_, _00851_, _00850_);
  and (_00853_, _00852_, _23597_);
  not (_00854_, _00853_);
  and (_00855_, _26746_, _26744_);
  not (_00856_, _00855_);
  and (_00857_, _00856_, _26747_);
  and (_00858_, _00857_, _26607_);
  not (_00859_, _00858_);
  and (_00860_, _00800_, _23538_);
  and (_00861_, _00860_, _23048_);
  and (_00862_, _00802_, _23217_);
  and (_00863_, _00862_, _23046_);
  nor (_00864_, _00863_, _00861_);
  nor (_00865_, _00864_, _23398_);
  and (_00866_, _00864_, _23398_);
  or (_00867_, _00866_, _23335_);
  nor (_00868_, _00867_, _00865_);
  and (_00869_, _23388_, _23173_);
  nor (_00870_, _23091_, _23316_);
  and (_00871_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_00872_, _00871_, _00870_);
  or (_00873_, _00872_, _23637_);
  nor (_00874_, _00873_, _00869_);
  not (_00875_, _00874_);
  nor (_00876_, _00875_, _00868_);
  and (_00877_, _00876_, _00859_);
  and (_00878_, _00877_, _00854_);
  nor (_00879_, _00878_, _00709_);
  and (_00880_, _26801_, _26072_);
  not (_00881_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_00882_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_00883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_00884_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_00885_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_00886_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_00887_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00888_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_00889_, _00888_, _00887_);
  and (_00890_, _00889_, _00886_);
  and (_00891_, _00890_, _00885_);
  and (_00892_, _00891_, _00884_);
  and (_00893_, _00892_, _00883_);
  and (_00894_, _00893_, _00882_);
  nor (_00895_, _00894_, _00881_);
  and (_00896_, _00894_, _00881_);
  nor (_00897_, _00896_, _00895_);
  not (_00898_, _00897_);
  and (_00899_, _00898_, _00045_);
  and (_00900_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_00901_, _00900_, _00899_);
  or (_00902_, _00901_, _00880_);
  nor (_00903_, _00902_, _00879_);
  nand (_00904_, _00903_, _26378_);
  or (_00905_, _00904_, _00845_);
  or (_00906_, _00905_, _00844_);
  and (_00907_, _00830_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00908_, _00830_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00909_, _00908_, _00907_);
  or (_00910_, _00909_, _26378_);
  and (_00911_, _00910_, _22773_);
  and (_26861_[11], _00911_, _00906_);
  not (_00912_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00913_, _00836_, _00834_);
  and (_00914_, _00913_, _00651_);
  and (_00915_, _00838_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00916_, _00915_, _00624_);
  nor (_00917_, _00916_, _00914_);
  nand (_00918_, _00917_, _00912_);
  or (_00920_, _00917_, _00912_);
  and (_00921_, _00920_, _00918_);
  and (_00922_, _00921_, _00040_);
  and (_00923_, _00352_, _24643_);
  nor (_00924_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00925_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _00912_);
  nor (_00926_, _00925_, _00924_);
  or (_00927_, _00926_, _00851_);
  and (_00928_, _00926_, _00851_);
  nor (_00929_, _00928_, _23598_);
  and (_00930_, _00929_, _00927_);
  or (_00931_, _26750_, _26748_);
  and (_00932_, _00931_, _26751_);
  and (_00933_, _00932_, _26607_);
  and (_00934_, _23388_, _23046_);
  and (_00935_, _00934_, _00862_);
  and (_00937_, _00860_, _23398_);
  and (_00938_, _00937_, _23048_);
  nor (_00939_, _00938_, _00935_);
  nand (_00940_, _00939_, _23185_);
  or (_00941_, _00939_, _23185_);
  and (_00942_, _00941_, _23067_);
  and (_00943_, _00942_, _00940_);
  or (_00945_, _23046_, _22977_);
  and (_00946_, _23185_, _23046_);
  nor (_00947_, _00946_, _23316_);
  and (_00948_, _00947_, _00945_);
  and (_00949_, _23635_, _23153_);
  and (_00950_, _23173_, _23060_);
  and (_00951_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_00952_, _00951_, _00950_);
  or (_00953_, _00952_, _00949_);
  or (_00955_, _00953_, _00948_);
  or (_00956_, _00955_, _00943_);
  or (_00957_, _00956_, _00933_);
  or (_00958_, _00957_, _00930_);
  and (_00959_, _00958_, _26799_);
  and (_00960_, _26801_, _26005_);
  not (_00961_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00962_, _00896_, _00961_);
  and (_00963_, _00896_, _00961_);
  or (_00964_, _00963_, _00962_);
  and (_00965_, _00964_, _00045_);
  and (_00966_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_00967_, _00966_, _00965_);
  or (_00969_, _00967_, _00960_);
  nor (_00970_, _00969_, _00959_);
  nand (_00971_, _00970_, _26378_);
  or (_00972_, _00971_, _00923_);
  or (_00973_, _00972_, _00922_);
  and (_00974_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_00975_, _00974_, _00830_);
  or (_00976_, _00907_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_00977_, _00976_, _00975_);
  or (_00978_, _00977_, _26378_);
  and (_00979_, _00978_, _22773_);
  and (_26861_[12], _00979_, _00973_);
  not (_00980_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00981_, _00913_, _00912_);
  nand (_00982_, _00981_, _00651_);
  nand (_00983_, _00915_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_00984_, _00983_, _00651_);
  and (_00985_, _00984_, _00982_);
  nand (_00986_, _00985_, _00980_);
  or (_00987_, _00985_, _00980_);
  and (_00988_, _00987_, _00986_);
  and (_00989_, _00988_, _00040_);
  and (_00990_, _00443_, _24643_);
  nor (_00991_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00992_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _00980_);
  nor (_00993_, _00992_, _00991_);
  or (_00994_, _00993_, _00928_);
  nand (_00995_, _00993_, _00928_);
  and (_00996_, _00995_, _23597_);
  and (_00997_, _00996_, _00994_);
  or (_00998_, _26752_, _26728_);
  and (_00999_, _00998_, _26753_);
  and (_01001_, _00999_, _26607_);
  and (_01002_, _00937_, _23185_);
  nor (_01003_, _01002_, _00935_);
  nor (_01004_, _01003_, _00946_);
  or (_01005_, _01004_, _23343_);
  nand (_01006_, _01004_, _23343_);
  and (_01007_, _01006_, _23067_);
  and (_01008_, _01007_, _01005_);
  and (_01009_, _23313_, _23048_);
  and (_01010_, _23343_, _23046_);
  or (_01011_, _01010_, _01009_);
  and (_01012_, _01011_, _22938_);
  and (_01013_, _23635_, _23147_);
  and (_01014_, _23343_, _23173_);
  and (_01015_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_01016_, _01015_, _01014_);
  or (_01017_, _01016_, _01013_);
  or (_01018_, _01017_, _01012_);
  or (_01019_, _01018_, _01008_);
  or (_01020_, _01019_, _01001_);
  or (_01021_, _01020_, _00997_);
  and (_01022_, _01021_, _26799_);
  and (_01023_, _26801_, _26019_);
  not (_01024_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01025_, _00963_, _01024_);
  and (_01026_, _00963_, _01024_);
  nor (_01027_, _01026_, _01025_);
  not (_01028_, _01027_);
  and (_01029_, _01028_, _00045_);
  and (_01030_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_01031_, _01030_, _01029_);
  or (_01032_, _01031_, _01023_);
  nor (_01033_, _01032_, _01022_);
  nand (_01034_, _01033_, _26378_);
  or (_01035_, _01034_, _00990_);
  or (_01036_, _01035_, _00989_);
  nand (_01037_, _00975_, _01024_);
  or (_01038_, _00975_, _01024_);
  and (_01040_, _01038_, _01037_);
  or (_01041_, _01040_, _26378_);
  and (_01042_, _01041_, _22773_);
  and (_26861_[13], _01042_, _01036_);
  not (_01043_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01044_, _00624_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01045_, _01044_, _00983_);
  or (_01046_, _00982_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01047_, _01046_, _01045_);
  nand (_01048_, _01047_, _01043_);
  or (_01049_, _01047_, _01043_);
  and (_01050_, _01049_, _01048_);
  and (_01051_, _01050_, _00040_);
  and (_01052_, _00564_, _24643_);
  and (_01053_, _23518_, _23173_);
  and (_01054_, _23635_, _23128_);
  and (_01055_, _01002_, _23324_);
  and (_01056_, _23343_, _23060_);
  and (_01057_, _01056_, _00935_);
  nor (_01058_, _01057_, _01055_);
  nor (_01059_, _01058_, _23518_);
  and (_01060_, _01058_, _23518_);
  or (_01061_, _01060_, _01059_);
  and (_01062_, _01061_, _23067_);
  and (_01063_, _23511_, _23048_);
  not (_01064_, _01063_);
  and (_01065_, _23520_, _23046_);
  nor (_01066_, _01065_, _23316_);
  and (_01067_, _01066_, _01064_);
  or (_01068_, _01067_, _01062_);
  or (_01069_, _01068_, _01054_);
  and (_01070_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_01071_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01072_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _01043_);
  nor (_01073_, _01072_, _01071_);
  not (_01074_, _01073_);
  and (_01075_, _01074_, _00995_);
  nor (_01076_, _01074_, _00995_);
  nor (_01077_, _01076_, _01075_);
  and (_01078_, _01077_, _23597_);
  and (_01079_, _26754_, _26722_);
  not (_01080_, _01079_);
  and (_01081_, _01080_, _26755_);
  and (_01082_, _01081_, _26607_);
  or (_01083_, _01082_, _01078_);
  or (_01084_, _01083_, _01070_);
  or (_01085_, _01084_, _01069_);
  or (_01086_, _01085_, _01053_);
  and (_01087_, _01086_, _26799_);
  and (_01088_, _26801_, _26108_);
  not (_01089_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01090_, _01026_, _01089_);
  and (_01091_, _01026_, _01089_);
  nor (_01092_, _01091_, _01090_);
  not (_01093_, _01092_);
  and (_01094_, _01093_, _00045_);
  and (_01095_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01096_, _01095_, _01094_);
  or (_01098_, _01096_, _01088_);
  nor (_01099_, _01098_, _01087_);
  nand (_01100_, _01099_, _26378_);
  or (_01101_, _01100_, _01052_);
  or (_01102_, _01101_, _01051_);
  and (_01103_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01104_, _01103_, _00766_);
  and (_01105_, _01104_, _00974_);
  and (_01106_, _01105_, _00645_);
  and (_01108_, _01106_, _25591_);
  nor (_01109_, _01108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_01110_, _01108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01112_, _01110_, _01109_);
  or (_01113_, _01112_, _26378_);
  and (_01114_, _01113_, _22773_);
  and (_26861_[14], _01114_, _01102_);
  and (_01116_, _24537_, _00818_);
  nor (_01117_, _00693_, _24664_);
  and (_01118_, _01117_, _01116_);
  not (_01119_, _01118_);
  nor (_01120_, _24610_, _24586_);
  and (_01121_, _24632_, _24561_);
  and (_01122_, _01121_, _01120_);
  not (_01123_, _01122_);
  not (_01124_, _24610_);
  nor (_01125_, _24632_, _24586_);
  and (_01127_, _01125_, _01124_);
  and (_01128_, _01127_, _24561_);
  nor (_01129_, _01128_, _24610_);
  and (_01130_, _01129_, _01123_);
  nor (_01132_, _01130_, _01119_);
  not (_01133_, _01132_);
  and (_01135_, _00750_, _24518_);
  and (_01136_, _01135_, _01117_);
  and (_01137_, _01116_, _00693_);
  and (_01139_, _01137_, _24664_);
  nor (_01140_, _01139_, _01136_);
  nor (_01141_, _01140_, _01123_);
  not (_01142_, _01141_);
  and (_01143_, _24632_, _24586_);
  and (_01144_, _01143_, _01124_);
  and (_01145_, _01144_, _24561_);
  and (_01146_, _24537_, _24518_);
  and (_01148_, _01146_, _00693_);
  and (_01149_, _01148_, _01145_);
  not (_01151_, _01145_);
  and (_01152_, _01116_, _24495_);
  and (_01153_, _01152_, _24664_);
  nor (_01154_, _24537_, _24495_);
  and (_01155_, _01154_, _24518_);
  and (_01156_, _01155_, _24664_);
  nor (_01157_, _01156_, _01153_);
  nor (_01158_, _01157_, _01151_);
  nor (_01159_, _01158_, _01149_);
  and (_01160_, _01159_, _01142_);
  and (_01161_, _00750_, _24495_);
  and (_01162_, _01161_, _00818_);
  nor (_01163_, _24495_, _24664_);
  and (_01164_, _01163_, _01116_);
  nor (_01166_, _01164_, _01162_);
  nor (_01167_, _01166_, _01123_);
  and (_01168_, _24495_, _24664_);
  and (_01169_, _01168_, _01135_);
  or (_01170_, _01143_, _01125_);
  nor (_01171_, _24632_, _24561_);
  nor (_01172_, _01171_, _24610_);
  and (_01173_, _01172_, _01170_);
  and (_01174_, _01173_, _01169_);
  nor (_01175_, _01174_, _01167_);
  not (_01176_, _01128_);
  nor (_01177_, _01164_, _01153_);
  nor (_01178_, _01177_, _01176_);
  not (_01179_, _24561_);
  and (_01180_, _01144_, _01179_);
  and (_01181_, _01180_, _01146_);
  nor (_01183_, _01181_, _01178_);
  and (_01185_, _01183_, _01175_);
  and (_01186_, _01185_, _01160_);
  and (_01187_, _01186_, _01133_);
  and (_01188_, _00693_, _24664_);
  and (_01189_, _01146_, _01188_);
  and (_01191_, _01189_, _01122_);
  nor (_01192_, _01169_, _01155_);
  nor (_01193_, _01192_, _01123_);
  nor (_01194_, _01193_, _01191_);
  not (_01195_, _01194_);
  and (_01196_, _01170_, _01155_);
  nor (_01197_, _01196_, _24664_);
  not (_01198_, _01197_);
  not (_01199_, _24664_);
  not (_01200_, _24632_);
  and (_01201_, _01200_, _24586_);
  nor (_01202_, _01201_, _01199_);
  not (_01203_, _01202_);
  nor (_01204_, _01155_, _01137_);
  nor (_01205_, _01204_, _24610_);
  and (_01206_, _01205_, _01203_);
  and (_01207_, _01206_, _01198_);
  nor (_01208_, _01207_, _01195_);
  nor (_01209_, _24537_, _24518_);
  and (_01210_, _01209_, _01163_);
  and (_01211_, _01210_, _01180_);
  not (_01212_, _01211_);
  and (_01213_, _01180_, _01139_);
  and (_01215_, _01171_, _01120_);
  and (_01216_, _01215_, _01169_);
  nor (_01217_, _01216_, _01213_);
  and (_01218_, _01217_, _01212_);
  and (_01219_, _01218_, _01208_);
  not (_01220_, _01137_);
  and (_01221_, _01162_, _24664_);
  nor (_01222_, _01221_, _01156_);
  and (_01223_, _01222_, _01220_);
  nor (_01224_, _01223_, _01124_);
  not (_01225_, _01224_);
  not (_01226_, _01180_);
  and (_01227_, _01209_, _01117_);
  nor (_01228_, _01227_, _01153_);
  nor (_01229_, _01228_, _01226_);
  not (_01230_, _01229_);
  and (_01231_, _01116_, _01199_);
  and (_01232_, _01201_, _01124_);
  and (_01233_, _01232_, _01231_);
  and (_01234_, _24632_, _01179_);
  and (_01235_, _01234_, _01120_);
  nor (_01236_, _01235_, _01233_);
  and (_01237_, _01236_, _01230_);
  and (_01238_, _01237_, _01225_);
  and (_01239_, _01215_, _01136_);
  and (_01240_, _01153_, _01122_);
  nor (_01241_, _01240_, _01239_);
  not (_01242_, _01241_);
  nor (_01243_, _01227_, _01139_);
  and (_01244_, _01243_, _01222_);
  nor (_01245_, _01244_, _01176_);
  nor (_01246_, _01245_, _01242_);
  and (_01247_, _01246_, _01238_);
  and (_01248_, _01247_, _01219_);
  not (_01249_, _01173_);
  and (_01250_, _01154_, _00818_);
  and (_01251_, _01250_, _24664_);
  and (_01252_, _01251_, _01180_);
  nor (_01253_, _01252_, _01136_);
  nor (_01254_, _01253_, _01249_);
  not (_01255_, _01254_);
  nor (_01256_, _01188_, _01117_);
  and (_01258_, _01256_, _01146_);
  and (_01259_, _01258_, _01122_);
  and (_01260_, _01221_, _01180_);
  nor (_01261_, _01260_, _01259_);
  and (_01262_, _01146_, _24495_);
  and (_01264_, _01262_, _01128_);
  not (_01265_, _01264_);
  and (_01266_, _01145_, _01139_);
  nor (_01267_, _01156_, _01118_);
  nor (_01268_, _01267_, _01226_);
  nor (_01269_, _01268_, _01266_);
  and (_01270_, _01269_, _01265_);
  and (_01271_, _01270_, _01261_);
  and (_01272_, _01271_, _01255_);
  and (_01273_, _01272_, _01248_);
  and (_01274_, _01273_, _01187_);
  and (_01275_, _01163_, _01135_);
  and (_01276_, _01275_, _01215_);
  not (_01278_, _01276_);
  nor (_01279_, _01201_, _24610_);
  not (_01280_, _01279_);
  and (_01281_, _01280_, _01139_);
  nor (_01282_, _01281_, _01191_);
  and (_01283_, _01282_, _01278_);
  and (_01284_, _01241_, _01217_);
  and (_01285_, _01284_, _01283_);
  and (_01286_, _01285_, _01271_);
  not (_01287_, _01286_);
  nor (_01288_, _01287_, _01274_);
  not (_01289_, _01288_);
  and (_01290_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01291_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01292_, _01291_, _01290_);
  and (_01293_, _01292_, _01289_);
  nor (_01294_, _01292_, _01289_);
  nor (_01295_, _01294_, _01293_);
  or (_01296_, _01295_, _24817_);
  or (_01297_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_01298_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01299_, _01298_, _01297_);
  and (_01300_, _01299_, _01296_);
  and (_01301_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _22773_);
  and (_01302_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_26862_[0], _01302_, _01300_);
  and (_01303_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01304_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01305_, _01304_, _01303_);
  and (_01306_, _01305_, _01290_);
  nor (_01307_, _01305_, _01290_);
  nor (_01308_, _01307_, _01306_);
  not (_01309_, _01308_);
  nor (_01310_, _01309_, _01274_);
  and (_01311_, _01309_, _01274_);
  nor (_01312_, _01311_, _01310_);
  and (_01313_, _01312_, _01293_);
  nor (_01314_, _01312_, _01293_);
  nor (_01315_, _01314_, _01313_);
  or (_01316_, _01315_, _24817_);
  or (_01317_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01318_, _01317_, _01298_);
  and (_01319_, _01318_, _01316_);
  and (_01320_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_26862_[1], _01320_, _01319_);
  and (_01321_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01322_, _01313_, _01310_);
  not (_01323_, _01322_);
  nor (_01324_, _01306_, _01303_);
  and (_01325_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01326_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01327_, _01326_, _01325_);
  not (_01328_, _01327_);
  nor (_01330_, _01328_, _01324_);
  and (_01331_, _01328_, _01324_);
  nor (_01332_, _01331_, _01330_);
  and (_01333_, _01332_, _01323_);
  nor (_01335_, _01332_, _01323_);
  nor (_01336_, _01335_, _01333_);
  or (_01338_, _01336_, _24817_);
  or (_01339_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01340_, _01339_, _01298_);
  and (_01341_, _01340_, _01338_);
  or (_26862_[2], _01341_, _01321_);
  nor (_01342_, _01330_, _01325_);
  nor (_01343_, _01342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01344_, _01342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_01345_, _01344_, _01343_);
  and (_01346_, _01345_, _01333_);
  nor (_01347_, _01345_, _01333_);
  nor (_01348_, _01347_, _01346_);
  or (_01349_, _01348_, _24817_);
  or (_01350_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01351_, _01350_, _01298_);
  and (_01352_, _01351_, _01349_);
  and (_01353_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_26862_[3], _01353_, _01352_);
  not (_01355_, _01342_);
  nand (_01356_, _01355_, _00888_);
  and (_01357_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_01358_, _00888_, _01357_);
  or (_01359_, _01358_, _01343_);
  and (_01360_, _01359_, _01356_);
  and (_01361_, _01360_, _01346_);
  or (_01362_, _01360_, _01346_);
  nand (_01363_, _01362_, _24816_);
  nor (_01364_, _01363_, _01361_);
  nor (_01365_, _24816_, _22939_);
  or (_01366_, _01365_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01367_, _01366_, _01364_);
  not (_01368_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01369_, _01368_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01370_, _01369_, _22773_);
  and (_26862_[4], _01370_, _01367_);
  or (_01371_, _01368_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_01372_, _01371_, _22773_);
  nand (_01373_, _01342_, _00888_);
  and (_01374_, _01373_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_01375_, _01342_, _00889_);
  or (_01376_, _01375_, _01374_);
  or (_01378_, _01376_, _01361_);
  and (_01379_, _01376_, _01360_);
  and (_01380_, _01379_, _01346_);
  nor (_01381_, _01380_, _24817_);
  and (_01382_, _01381_, _01378_);
  nor (_01383_, _24816_, _23296_);
  or (_01384_, _01383_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01385_, _01384_, _01382_);
  and (_26862_[5], _01385_, _01372_);
  and (_01386_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_01387_, _01375_, _00886_);
  and (_01388_, _01342_, _00890_);
  or (_01389_, _01388_, _01387_);
  and (_01390_, _01389_, _01380_);
  nor (_01391_, _01389_, _01380_);
  nor (_01393_, _01391_, _01390_);
  or (_01394_, _01393_, _24817_);
  or (_01395_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01396_, _01395_, _01298_);
  and (_01397_, _01396_, _01394_);
  or (_26862_[6], _01397_, _01386_);
  and (_01399_, _01342_, _00891_);
  nor (_01400_, _01388_, _00885_);
  nor (_01401_, _01400_, _01399_);
  not (_01403_, _01401_);
  and (_01404_, _01403_, _01390_);
  nor (_01405_, _01403_, _01390_);
  nor (_01406_, _01405_, _01404_);
  or (_01407_, _01406_, _24817_);
  or (_01408_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01409_, _01408_, _01298_);
  and (_01410_, _01409_, _01407_);
  and (_01411_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_26862_[7], _01411_, _01410_);
  nor (_01412_, _01399_, _00884_);
  and (_01413_, _01342_, _00892_);
  or (_01414_, _01413_, _01412_);
  and (_01415_, _01414_, _01404_);
  nor (_01417_, _01414_, _01404_);
  nor (_01418_, _01417_, _01415_);
  or (_01419_, _01418_, _24817_);
  or (_01420_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01421_, _01420_, _01298_);
  and (_01422_, _01421_, _01419_);
  and (_01423_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_26862_[8], _01423_, _01422_);
  or (_01425_, _01413_, _00883_);
  nand (_01426_, _01413_, _00883_);
  and (_01427_, _01426_, _01425_);
  not (_01428_, _01427_);
  and (_01429_, _01428_, _01415_);
  nor (_01430_, _01428_, _01415_);
  nor (_01431_, _01430_, _01429_);
  or (_01432_, _01431_, _24817_);
  or (_01433_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_01434_, _01433_, _01298_);
  and (_01435_, _01434_, _01432_);
  and (_01436_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_26862_[9], _01436_, _01435_);
  and (_01437_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01438_, _00893_, _00882_);
  nor (_01439_, _01438_, _00894_);
  nand (_01440_, _01355_, _00893_);
  and (_01441_, _01440_, _01439_);
  and (_01442_, _01355_, _00894_);
  nor (_01443_, _01442_, _01441_);
  and (_01444_, _01443_, _01429_);
  nor (_01445_, _01443_, _01429_);
  nor (_01446_, _01445_, _01444_);
  or (_01447_, _01446_, _24817_);
  or (_01448_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01449_, _01448_, _01298_);
  and (_01450_, _01449_, _01447_);
  or (_26862_[10], _01450_, _01437_);
  nor (_01451_, _01442_, _00898_);
  and (_01452_, _01355_, _00896_);
  nor (_01453_, _01452_, _01451_);
  and (_01454_, _01453_, _01444_);
  nor (_01455_, _01453_, _01444_);
  nor (_01456_, _01455_, _01454_);
  or (_01457_, _01456_, _24817_);
  or (_01458_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01459_, _01458_, _01298_);
  and (_01460_, _01459_, _01457_);
  and (_01461_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_26862_[11], _01461_, _01460_);
  or (_01462_, _01452_, _00964_);
  and (_01463_, _01452_, _00961_);
  not (_01464_, _01463_);
  and (_01465_, _01464_, _01462_);
  and (_01466_, _01465_, _01454_);
  nor (_01467_, _01465_, _01454_);
  nor (_01468_, _01467_, _01466_);
  or (_01469_, _01468_, _24817_);
  or (_01470_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01471_, _01470_, _01298_);
  and (_01472_, _01471_, _01469_);
  and (_01473_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_26862_[12], _01473_, _01472_);
  and (_01474_, _01464_, _01027_);
  and (_01475_, _01355_, _01026_);
  nor (_01476_, _01475_, _01474_);
  and (_01477_, _01476_, _01466_);
  nor (_01478_, _01476_, _01466_);
  nor (_01479_, _01478_, _01477_);
  or (_01480_, _01479_, _24817_);
  or (_01481_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01482_, _01481_, _01298_);
  and (_01483_, _01482_, _01480_);
  and (_01484_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_26862_[13], _01484_, _01483_);
  and (_01485_, _01301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01486_, _01475_, _01093_);
  and (_01487_, _01355_, _01091_);
  nor (_01488_, _01487_, _01486_);
  or (_01489_, _01488_, _01477_);
  nand (_01490_, _01488_, _01477_);
  and (_01491_, _01490_, _01489_);
  or (_01492_, _01491_, _24817_);
  or (_01493_, _24816_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01494_, _01493_, _01298_);
  and (_01495_, _01494_, _01492_);
  or (_26862_[14], _01495_, _01485_);
  and (_01496_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_01497_, _25490_, _23751_);
  or (_22681_, _01497_, _01496_);
  nor (_01498_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_01500_, _01499_, _01498_);
  nor (_01501_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_01502_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_01503_, _01502_, _01501_);
  and (_01504_, _01503_, _01500_);
  and (_01505_, _01504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01506_, _01505_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_26866_[0], _01506_, _22773_);
  and (_01508_, _01504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01509_, _01508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_26866_[1], _01509_, _22773_);
  and (_01510_, _01504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_01511_, _01510_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_26866_[2], _01511_, _22773_);
  and (_01512_, _01504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_01513_, _01512_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_26866_[3], _01513_, _22773_);
  and (_01514_, _01504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01515_, _01514_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_26866_[4], _01515_, _22773_);
  and (_01516_, _01504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_01517_, _01516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_26866_[5], _01517_, _22773_);
  and (_01518_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22773_);
  and (_01520_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _22773_);
  and (_01522_, _01520_, _01504_);
  or (_26866_[6], _01522_, _01518_);
  nor (_01524_, _01288_, _24883_);
  nand (_01525_, _01524_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_01526_, _01524_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_01527_, _01526_, _01298_);
  and (_26867_[0], _01527_, _01525_);
  and (_01528_, _01289_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01529_, _01274_, _24472_);
  and (_01530_, _01274_, _24472_);
  nor (_01531_, _01530_, _01529_);
  and (_01532_, _01531_, _01528_);
  nor (_01533_, _01531_, _01528_);
  nor (_01534_, _01533_, _01532_);
  or (_01535_, _01534_, _24883_);
  or (_01536_, _23760_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01537_, _01536_, _01298_);
  and (_26867_[1], _01537_, _01535_);
  and (_01538_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_01539_, _25490_, _23693_);
  or (_22682_, _01539_, _01538_);
  and (_01541_, _25164_, _23930_);
  and (_01542_, _01541_, _24027_);
  not (_01543_, _01541_);
  and (_01544_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_22683_, _01544_, _01542_);
  and (_01545_, _01541_, _23920_);
  and (_01546_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_22684_, _01546_, _01545_);
  nor (_26858_[3], _26071_, rst);
  not (_01548_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_01550_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _01548_);
  and (_01551_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01552_, _01551_, _01550_);
  and (_26870_[0], _01552_, _22773_);
  and (_01553_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _01548_);
  and (_01554_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01555_, _01554_, _01553_);
  and (_26870_[1], _01555_, _22773_);
  and (_01556_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _01548_);
  and (_01557_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01558_, _01557_, _01556_);
  and (_26870_[2], _01558_, _22773_);
  and (_01559_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _01548_);
  and (_01560_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01562_, _01560_, _01559_);
  and (_26870_[3], _01562_, _22773_);
  and (_01563_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _01548_);
  and (_01564_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01565_, _01564_, _01563_);
  and (_26870_[4], _01565_, _22773_);
  and (_01566_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _01548_);
  and (_01567_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01568_, _01567_, _01566_);
  and (_26870_[5], _01568_, _22773_);
  and (_01569_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _01548_);
  and (_01570_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01571_, _01570_, _01569_);
  and (_26870_[6], _01571_, _22773_);
  not (_01572_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01573_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01574_, _01573_, _01572_);
  and (_01575_, _01573_, _01572_);
  nor (_01577_, _01575_, _01574_);
  and (_26873_[0], _01577_, _22773_);
  nor (_01578_, _01574_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01579_, _01574_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01580_, _01579_, _01578_);
  nor (_26873_[1], _01580_, rst);
  and (_01582_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01583_, _01582_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01584_, _01582_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01585_, _01584_, _01583_);
  or (_01586_, _01585_, _01573_);
  and (_26873_[2], _01586_, _22773_);
  and (_01587_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_01588_, _25524_, _25526_);
  or (_01589_, _01588_, _01587_);
  and (_26875_[0], _01589_, _22773_);
  and (_01590_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_01591_, _25524_, _25530_);
  or (_01592_, _01591_, _01590_);
  and (_26875_[1], _01592_, _22773_);
  and (_01594_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_01595_, _25524_, _25534_);
  or (_01597_, _01595_, _01594_);
  and (_26875_[2], _01597_, _22773_);
  and (_01599_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_01601_, _25524_, _25538_);
  or (_01602_, _01601_, _01599_);
  and (_26875_[3], _01602_, _22773_);
  and (_01604_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_01605_, _25524_, _25542_);
  or (_01606_, _01605_, _01604_);
  and (_26875_[4], _01606_, _22773_);
  and (_01607_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_01608_, _25524_, _25546_);
  or (_01609_, _01608_, _01607_);
  and (_26875_[5], _01609_, _22773_);
  and (_01610_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_01611_, _25524_, _25551_);
  or (_01612_, _01611_, _01610_);
  and (_26875_[6], _01612_, _22773_);
  and (_01613_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_01614_, _25524_, _25557_);
  or (_01615_, _01614_, _01613_);
  and (_26875_[7], _01615_, _22773_);
  and (_01616_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_01617_, _25524_, _25561_);
  or (_01618_, _01617_, _01616_);
  and (_26875_[8], _01618_, _22773_);
  and (_01619_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_01620_, _25524_, _25566_);
  or (_01621_, _01620_, _01619_);
  and (_26875_[9], _01621_, _22773_);
  and (_01622_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_01624_, _25524_, _25570_);
  or (_01625_, _01624_, _01622_);
  and (_26875_[10], _01625_, _22773_);
  and (_01626_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_01627_, _25524_, _25574_);
  or (_01628_, _01627_, _01626_);
  and (_26875_[11], _01628_, _22773_);
  and (_01629_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_01630_, _25524_, _25578_);
  or (_01631_, _01630_, _01629_);
  and (_26875_[12], _01631_, _22773_);
  and (_01632_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_01633_, _25524_, _25582_);
  or (_01634_, _01633_, _01632_);
  and (_26875_[13], _01634_, _22773_);
  and (_01635_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_01636_, _25524_, _25586_);
  or (_01637_, _01636_, _01635_);
  and (_26875_[14], _01637_, _22773_);
  or (_01638_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_01639_, _25591_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_01640_, _01639_, _22773_);
  and (_26875_[15], _01640_, _01638_);
  and (_01641_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01642_, _25524_, _25595_);
  or (_01643_, _01642_, _01641_);
  and (_26875_[16], _01643_, _22773_);
  and (_01644_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01645_, _25524_, _25600_);
  or (_01646_, _01645_, _01644_);
  and (_26875_[17], _01646_, _22773_);
  and (_01647_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01648_, _25524_, _25605_);
  or (_01650_, _01648_, _01647_);
  and (_26875_[18], _01650_, _22773_);
  and (_01651_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01652_, _25524_, _25609_);
  or (_01653_, _01652_, _01651_);
  and (_26875_[19], _01653_, _22773_);
  and (_01654_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01655_, _25524_, _25613_);
  or (_01656_, _01655_, _01654_);
  and (_26875_[20], _01656_, _22773_);
  and (_01657_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01658_, _25524_, _25618_);
  or (_01659_, _01658_, _01657_);
  and (_26875_[21], _01659_, _22773_);
  and (_01660_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01661_, _25524_, _25622_);
  or (_01662_, _01661_, _01660_);
  and (_26875_[22], _01662_, _22773_);
  or (_01663_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_01664_, _25591_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_01665_, _01664_, _22773_);
  and (_26875_[23], _01665_, _01663_);
  and (_01666_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01667_, _25524_, _25630_);
  or (_01668_, _01667_, _01666_);
  and (_26875_[24], _01668_, _22773_);
  and (_01669_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01670_, _25524_, _25634_);
  or (_01671_, _01670_, _01669_);
  and (_26875_[25], _01671_, _22773_);
  and (_01672_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01673_, _25524_, _25638_);
  or (_01674_, _01673_, _01672_);
  and (_26875_[26], _01674_, _22773_);
  and (_01675_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01676_, _25524_, _25642_);
  or (_01678_, _01676_, _01675_);
  and (_26875_[27], _01678_, _22773_);
  and (_01679_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01680_, _25524_, _25646_);
  or (_01681_, _01680_, _01679_);
  and (_26875_[28], _01681_, _22773_);
  and (_01682_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01683_, _25524_, _25650_);
  or (_01684_, _01683_, _01682_);
  and (_26875_[29], _01684_, _22773_);
  and (_01685_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01686_, _25524_, _25654_);
  or (_01687_, _01686_, _01685_);
  and (_26875_[30], _01687_, _22773_);
  and (_01688_, _24740_, _24027_);
  and (_01689_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_22685_, _01689_, _01688_);
  nand (_01691_, _24561_, _23759_);
  or (_01692_, _23759_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_01693_, _01692_, _22773_);
  and (_26835_[0], _01693_, _01691_);
  and (_01694_, _25503_, _24053_);
  and (_01695_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_26917_, _01695_, _01694_);
  and (_01697_, _23983_, _23925_);
  and (_01698_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_22686_, _01698_, _01697_);
  and (_01699_, _25482_, _23715_);
  and (_01700_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_27228_, _01700_, _01699_);
  and (_01701_, _23890_, _23719_);
  and (_01702_, _01701_, _24027_);
  not (_01703_, _01701_);
  and (_01704_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or (_22687_, _01704_, _01702_);
  and (_01705_, _24319_, _23983_);
  and (_01707_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_22688_, _01707_, _01705_);
  and (_01709_, _25175_, _24157_);
  and (_01711_, _01709_, _24053_);
  not (_01712_, _01709_);
  and (_01713_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_22689_, _01713_, _01711_);
  and (_01714_, _01541_, _23983_);
  and (_01715_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_22690_, _01715_, _01714_);
  nor (_01716_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_01717_, _01716_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not (_01718_, _01717_);
  or (_01719_, _01718_, _26798_);
  or (_01720_, _01717_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_01721_, _01720_, _22773_);
  and (_26879_[0], _01721_, _01719_);
  or (_01722_, _01718_, _00101_);
  or (_01723_, _01717_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_01724_, _01723_, _22773_);
  and (_26879_[1], _01724_, _01722_);
  or (_01725_, _01718_, _00183_);
  or (_01726_, _01717_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_01727_, _01726_, _22773_);
  and (_26879_[2], _01727_, _01725_);
  or (_01728_, _01718_, _00277_);
  or (_01729_, _01717_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_01730_, _01729_, _22773_);
  and (_26879_[3], _01730_, _01728_);
  and (_26831_[3], _24610_, _22773_);
  and (_01731_, _24027_, _23892_);
  and (_01732_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or (_27224_, _01732_, _01731_);
  and (_01733_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_01734_, _25490_, _23715_);
  or (_22691_, _01734_, _01733_);
  and (_01735_, _24758_, _24332_);
  and (_01736_, _01735_, _24373_);
  nand (_01737_, _01736_, _23681_);
  and (_01738_, _25320_, _24406_);
  not (_01739_, _01738_);
  or (_01740_, _01736_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_01741_, _01740_, _01739_);
  and (_01742_, _01741_, _01737_);
  nor (_01743_, _01739_, _24017_);
  or (_01744_, _01743_, _01742_);
  and (_22692_, _01744_, _22773_);
  and (_01745_, _24097_, _23706_);
  and (_01746_, _01745_, _23900_);
  not (_01747_, _01745_);
  and (_01748_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or (_22693_, _01748_, _01746_);
  nor (_01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_01750_, _01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _22773_);
  and (_01752_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_22694_, _01752_, _01750_);
  and (_01753_, _01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_01754_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_22695_, _01754_, _01753_);
  and (_01755_, _01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_01756_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_22696_, _01756_, _01755_);
  and (_01757_, _23983_, _23939_);
  and (_01758_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or (_22697_, _01758_, _01757_);
  and (_01759_, _24274_, _23909_);
  and (_01760_, _01759_, _24053_);
  not (_01761_, _01759_);
  and (_01762_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  or (_22698_, _01762_, _01760_);
  and (_01764_, _01541_, _23751_);
  and (_01765_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_26899_, _01765_, _01764_);
  and (_01766_, _01541_, _24053_);
  and (_01767_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_22699_, _01767_, _01766_);
  and (_01768_, _24235_, _24084_);
  not (_01769_, _01768_);
  and (_01770_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_01771_, _01768_, _23920_);
  or (_26998_, _01771_, _01770_);
  and (_22700_, _01518_, _24855_);
  and (_01772_, _24855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_01773_, _01772_, _24920_);
  and (_22701_, _01773_, _22773_);
  or (_01774_, _25075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01775_, _25074_, _24851_);
  and (_01776_, _01775_, _01774_);
  not (_01777_, _24851_);
  or (_01778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_01779_, _01778_, _01777_);
  or (_01780_, _01779_, _01776_);
  and (_01781_, _01780_, _24844_);
  and (_01783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _24859_);
  and (_01784_, _24851_, _24837_);
  or (_01785_, _01784_, _24843_);
  and (_01786_, _01785_, _01783_);
  nor (_01787_, _01786_, _24854_);
  nand (_01788_, _01787_, _24879_);
  or (_01789_, _01788_, _01781_);
  or (_01790_, _25057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01791_, _01790_, _25061_);
  not (_01792_, _24869_);
  and (_01793_, _01778_, _01792_);
  or (_01794_, _01793_, _01791_);
  and (_01795_, _01794_, _24866_);
  and (_01796_, _24875_, _24869_);
  or (_01797_, _01796_, _24865_);
  and (_01798_, _01797_, _01783_);
  or (_01799_, _01798_, _24879_);
  or (_01800_, _01799_, _01795_);
  and (_01801_, _01800_, _01789_);
  or (_01802_, _01801_, _24855_);
  or (_01803_, _24920_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01804_, _01803_, _22773_);
  and (_22702_, _01804_, _01802_);
  or (_01805_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _24859_);
  or (_01806_, _01805_, _24869_);
  and (_01807_, _01806_, _24866_);
  or (_01808_, _24925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01809_, _01808_, _24924_);
  or (_01810_, _01809_, _01792_);
  and (_01811_, _01810_, _01807_);
  and (_01812_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_01813_, _01812_, _01797_);
  or (_01814_, _01813_, _24879_);
  or (_01815_, _01814_, _01811_);
  or (_01816_, _24950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01817_, _24949_, _24851_);
  and (_01818_, _01817_, _01816_);
  and (_01819_, _01805_, _01777_);
  or (_01820_, _01819_, _01818_);
  and (_01821_, _01820_, _24844_);
  and (_01822_, _01812_, _01785_);
  nor (_01823_, _01822_, _24854_);
  nand (_01824_, _01823_, _24879_);
  or (_01825_, _01824_, _01821_);
  and (_01826_, _01825_, _01815_);
  or (_01827_, _01826_, _24855_);
  or (_01829_, _24920_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01830_, _01829_, _22773_);
  and (_22703_, _01830_, _01827_);
  and (_01831_, _24411_, _23208_);
  or (_01832_, _01831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_01833_, _01832_, _24417_);
  nand (_01834_, _01831_, _23681_);
  and (_01835_, _01834_, _01833_);
  nor (_01836_, _24417_, _23357_);
  or (_01837_, _01836_, _01835_);
  and (_22704_, _01837_, _22773_);
  and (_01838_, _24431_, _24333_);
  not (_01839_, _24333_);
  or (_01840_, _24425_, _01839_);
  or (_01841_, _01840_, _24337_);
  and (_01842_, _01841_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01843_, _01842_, _24344_);
  or (_01844_, _01843_, _01838_);
  or (_01846_, _24347_, _23205_);
  and (_01847_, _01846_, _22773_);
  and (_22705_, _01847_, _01844_);
  and (_01848_, _01541_, _23715_);
  and (_01849_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_22707_, _01849_, _01848_);
  and (_01851_, _01541_, _23693_);
  and (_01852_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_22708_, _01852_, _01851_);
  and (_01854_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_01855_, _01768_, _23983_);
  or (_27000_, _01855_, _01854_);
  and (_01856_, _23450_, _22823_);
  and (_01857_, _01856_, _22927_);
  and (_01858_, _01857_, _25673_);
  and (_01859_, _01858_, _23247_);
  not (_01860_, _01858_);
  and (_01861_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_27318_, _01861_, _01859_);
  and (_01862_, _01858_, _23744_);
  and (_01863_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_27317_, _01863_, _01862_);
  and (_01864_, _01858_, _24788_);
  and (_01865_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_22709_, _01865_, _01864_);
  and (_01866_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_01867_, _01768_, _23751_);
  or (_22710_, _01867_, _01866_);
  and (_01868_, _01858_, _23920_);
  and (_01869_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_22711_, _01869_, _01868_);
  and (_01870_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_01871_, _01768_, _24053_);
  or (_22712_, _01871_, _01870_);
  and (_01872_, _01858_, _23900_);
  and (_01873_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_22713_, _01873_, _01872_);
  and (_01874_, _01858_, _23413_);
  and (_01875_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_22714_, _01875_, _01874_);
  and (_01876_, _25164_, _24108_);
  and (_01877_, _01876_, _23693_);
  not (_01878_, _01876_);
  and (_01879_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_22715_, _01879_, _01877_);
  and (_01880_, _01876_, _23900_);
  and (_01881_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_22716_, _01881_, _01880_);
  and (_01882_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_01883_, _01768_, _23715_);
  or (_22717_, _01883_, _01882_);
  and (_01885_, _24677_, _24648_);
  and (_01886_, _23760_, _22773_);
  nand (_01887_, _01886_, _01885_);
  nand (_01888_, _01886_, _24696_);
  or (_01889_, _01888_, _26241_);
  and (_26833_[1], _01889_, _01887_);
  and (_01890_, _24268_, _23983_);
  and (_01891_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or (_22719_, _01891_, _01890_);
  and (_01892_, _23988_, _23983_);
  and (_01893_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_22720_, _01893_, _01892_);
  not (_01894_, _23759_);
  or (_01895_, _24610_, _01894_);
  or (_01896_, _23759_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_01897_, _01896_, _22773_);
  and (_26835_[3], _01897_, _01895_);
  nand (_01898_, _24495_, _23759_);
  or (_01900_, _23759_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_01901_, _01900_, _22773_);
  and (_26835_[5], _01901_, _01898_);
  and (_01902_, _01876_, _23715_);
  and (_01903_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_22721_, _01903_, _01902_);
  and (_01904_, _24027_, _23988_);
  and (_01905_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_22722_, _01905_, _01904_);
  and (_01906_, _01745_, _23920_);
  and (_01907_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or (_22723_, _01907_, _01906_);
  and (_01908_, _24157_, _23719_);
  and (_01909_, _01908_, _23693_);
  not (_01910_, _01908_);
  and (_01911_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or (_22724_, _01911_, _01909_);
  and (_01913_, _01908_, _23715_);
  and (_01914_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or (_22725_, _01914_, _01913_);
  and (_01915_, _25482_, _23900_);
  and (_01916_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_27229_, _01916_, _01915_);
  and (_01917_, _23983_, _23910_);
  and (_01918_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_27110_, _01918_, _01917_);
  and (_01919_, _25428_, _23920_);
  and (_01920_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_22726_, _01920_, _01919_);
  and (_01921_, _01908_, _23900_);
  and (_01922_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or (_22727_, _01922_, _01921_);
  and (_01923_, _01701_, _23715_);
  and (_01924_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or (_22728_, _01924_, _01923_);
  and (_01925_, _23925_, _23693_);
  and (_01926_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_22729_, _01926_, _01925_);
  and (_01927_, _25164_, _24145_);
  and (_01928_, _01927_, _23983_);
  not (_01929_, _01927_);
  and (_01931_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_22730_, _01931_, _01928_);
  and (_01932_, _24123_, _23719_);
  and (_01933_, _01932_, _24053_);
  not (_01934_, _01932_);
  and (_01935_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_22731_, _01935_, _01933_);
  and (_01936_, _24388_, _24068_);
  and (_01937_, _01936_, _24027_);
  not (_01938_, _01936_);
  and (_01939_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_22732_, _01939_, _01937_);
  and (_01940_, _25169_, _23751_);
  and (_01941_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_22734_, _01941_, _01940_);
  and (_01942_, _01876_, _23983_);
  and (_01944_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_27303_, _01944_, _01942_);
  and (_01945_, _01876_, _24027_);
  and (_01946_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_27302_, _01946_, _01945_);
  and (_01947_, _01876_, _23920_);
  and (_01948_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_22735_, _01948_, _01947_);
  and (_01949_, _23988_, _23900_);
  and (_01951_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_22736_, _01951_, _01949_);
  and (_01952_, _23905_, _23453_);
  and (_01953_, _01952_, _23693_);
  not (_01954_, _01952_);
  and (_01955_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or (_22737_, _01955_, _01953_);
  and (_01957_, _25364_, _24027_);
  and (_01958_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or (_22738_, _01958_, _01957_);
  and (_01959_, _24343_, _22857_);
  or (_01960_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_01961_, _01960_, _22773_);
  not (_01962_, _01959_);
  or (_01963_, _01962_, _23247_);
  and (_22739_, _01963_, _01961_);
  or (_01964_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_01965_, _01964_, _22773_);
  or (_01966_, _01962_, _23413_);
  and (_22740_, _01966_, _01965_);
  not (_01967_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_01969_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_01970_, _25320_, _22920_);
  and (_01971_, _01970_, _01969_);
  and (_01972_, _01971_, _01967_);
  and (_01974_, _01972_, _26145_);
  nor (_01975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_01976_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_01977_, _01976_, _01975_);
  not (_01978_, _01975_);
  and (_01979_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_01980_, _01979_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_01981_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_01982_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_01983_, _01982_, _01981_);
  and (_01984_, _01983_, _01980_);
  nor (_01986_, _01984_, _01977_);
  not (_01987_, _01986_);
  and (_01988_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_01990_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_01991_, _01990_, _01988_);
  nor (_01992_, _01991_, _01970_);
  and (_01994_, _01978_, _01970_);
  not (_01995_, _01994_);
  nor (_01996_, _01995_, _24017_);
  or (_01997_, _01996_, _01992_);
  or (_01998_, _01997_, _01974_);
  and (_22741_, _01998_, _22773_);
  nand (_01999_, _01994_, _23976_);
  and (_02000_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_02001_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_02003_, _02001_, _02000_);
  or (_02004_, _02003_, _01970_);
  and (_02005_, _02004_, _22773_);
  and (_22742_, _02005_, _01999_);
  and (_02006_, _01972_, _23744_);
  and (_02007_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_02008_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02009_, _02008_, _02007_);
  nor (_02010_, _02009_, _01970_);
  and (_02011_, _01994_, _24788_);
  or (_02012_, _02011_, _02010_);
  or (_02013_, _02012_, _02006_);
  and (_22743_, _02013_, _22773_);
  and (_02014_, _01972_, _23247_);
  and (_02015_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_02016_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_02017_, _02016_, _02015_);
  nor (_02018_, _02017_, _01970_);
  and (_02019_, _01994_, _23744_);
  or (_02020_, _02019_, _02018_);
  or (_02021_, _02020_, _02014_);
  and (_22744_, _02021_, _22773_);
  not (_02022_, _24184_);
  nor (_02023_, _02022_, _23681_);
  not (_02024_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_02025_, _24184_, _02024_);
  nand (_02026_, _02025_, _01735_);
  or (_02027_, _02026_, _02023_);
  nor (_02028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_02029_, _02028_, _01978_);
  and (_02030_, _02029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_02031_, _02029_, _02024_);
  or (_02032_, _02031_, _02030_);
  or (_02033_, _02032_, _01735_);
  and (_02034_, _02033_, _02027_);
  or (_02035_, _02034_, _01738_);
  or (_02036_, _01739_, _23247_);
  and (_02037_, _02036_, _22773_);
  and (_22745_, _02037_, _02035_);
  and (_02038_, _01735_, _23208_);
  nand (_02039_, _02038_, _23681_);
  or (_02040_, _02038_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_02041_, _02040_, _01739_);
  and (_02043_, _02041_, _02039_);
  nor (_02044_, _01739_, _23357_);
  or (_02045_, _02044_, _02043_);
  and (_22746_, _02045_, _22773_);
  or (_02046_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_02047_, _02046_, _22773_);
  nand (_02048_, _01959_, _23357_);
  and (_22747_, _02048_, _02047_);
  and (_02049_, _01962_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_02050_, _01959_, _24788_);
  or (_02051_, _02050_, _02049_);
  and (_22748_, _02051_, _22773_);
  and (_02052_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_02053_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_02054_, _02053_, _02052_);
  nor (_02055_, _02054_, _01970_);
  or (_02056_, _01969_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_02058_, _02056_, _01994_);
  or (_02059_, _02058_, _02055_);
  and (_22749_, _02059_, _22773_);
  and (_02060_, _01972_, _25813_);
  and (_02062_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02063_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_02064_, _02063_, _02062_);
  nor (_02066_, _02064_, _01970_);
  and (_02067_, _01994_, _23205_);
  or (_02068_, _02067_, _02066_);
  or (_02069_, _02068_, _02060_);
  and (_22750_, _02069_, _22773_);
  and (_02070_, _01975_, _01970_);
  and (_02071_, _02070_, _23413_);
  and (_02072_, _01994_, _23247_);
  and (_02073_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_02074_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02075_, _02074_, _02073_);
  nor (_02076_, _02075_, _01970_);
  or (_02077_, _02076_, _02072_);
  or (_02079_, _02077_, _02071_);
  and (_22751_, _02079_, _22773_);
  and (_02080_, _24405_, _23708_);
  not (_02081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02082_, _24405_, _02081_);
  nand (_02083_, _02082_, _01735_);
  or (_02084_, _02083_, _02080_);
  not (_02085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_02086_, _02085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_02087_, _02086_, _01975_);
  and (_02088_, _02087_, _02028_);
  or (_02089_, _02088_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02090_, _02089_, _01735_);
  and (_02091_, _02090_, _02084_);
  or (_02092_, _02091_, _01738_);
  nand (_02093_, _01738_, _24047_);
  and (_02094_, _02093_, _22773_);
  and (_22752_, _02094_, _02092_);
  and (_02096_, _01735_, _23250_);
  nand (_02097_, _02096_, _23681_);
  or (_02098_, _02096_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_02099_, _02098_, _01739_);
  and (_02100_, _02099_, _02097_);
  and (_02101_, _01738_, _23413_);
  or (_02103_, _02101_, _02100_);
  and (_22753_, _02103_, _22773_);
  or (_02104_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_02105_, _02104_, _22773_);
  nand (_02106_, _01959_, _24017_);
  and (_22754_, _02106_, _02105_);
  or (_02109_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_02110_, _02109_, _22773_);
  or (_02111_, _01962_, _23744_);
  and (_22755_, _02111_, _02110_);
  and (_02112_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_02113_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_02114_, _02113_, _02112_);
  nor (_02115_, _02114_, _01970_);
  nor (_02116_, _01995_, _23357_);
  and (_02117_, _02070_, _25833_);
  or (_02118_, _02117_, _02116_);
  or (_02119_, _02118_, _02115_);
  and (_22756_, _02119_, _22773_);
  and (_02120_, _02070_, _23205_);
  and (_02121_, _01994_, _23413_);
  and (_02122_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02123_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_02124_, _02123_, _02122_);
  nor (_02125_, _02124_, _01970_);
  or (_02126_, _02125_, _02121_);
  or (_02127_, _02126_, _02120_);
  and (_22757_, _02127_, _22773_);
  or (_02128_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_02129_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_02130_, _02129_, _01984_);
  and (_02132_, _02130_, _02128_);
  nor (_02133_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor (_02134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02135_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02136_, _02135_, _02134_);
  and (_02137_, _02136_, _02133_);
  nor (_02138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02139_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02140_, _02139_, _02138_);
  and (_02141_, _02140_, _01977_);
  and (_02142_, _02141_, _02137_);
  and (_02143_, _02142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_02144_, _02143_, _02132_);
  nor (_02145_, _02144_, _01970_);
  and (_02146_, _02070_, _24788_);
  or (_02147_, _02146_, _02145_);
  and (_22758_, _02147_, _22773_);
  or (_02148_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_02149_, _02148_, _01735_);
  and (_02150_, _23708_, _22895_);
  not (_02151_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_02152_, _22895_, _02151_);
  nand (_02153_, _02152_, _01735_);
  or (_02154_, _02153_, _02150_);
  and (_02155_, _02154_, _02149_);
  or (_02156_, _02155_, _01738_);
  or (_02157_, _01739_, _23744_);
  and (_02158_, _02157_, _22773_);
  and (_22759_, _02158_, _02156_);
  and (_02159_, _24432_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02160_, _02159_, _24431_);
  and (_02161_, _02160_, _01735_);
  not (_02162_, _01735_);
  or (_02163_, _02162_, _24426_);
  and (_02164_, _02163_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02165_, _02164_, _01738_);
  or (_02166_, _02165_, _02161_);
  or (_02167_, _01739_, _23205_);
  and (_02168_, _02167_, _22773_);
  and (_22760_, _02168_, _02166_);
  and (_02170_, _24084_, _23890_);
  not (_02171_, _02170_);
  and (_02172_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and (_02173_, _02170_, _23900_);
  or (_22761_, _02173_, _02172_);
  or (_02174_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_02175_, _02174_, _22773_);
  or (_02176_, _01962_, _23205_);
  and (_22762_, _02176_, _02175_);
  not (_02177_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_02178_, _01975_, _02177_);
  and (_02179_, _02178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_02181_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_02182_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _02181_);
  not (_02183_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02184_, _02183_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_02185_, _02184_, _02182_);
  and (_02186_, _02185_, _02179_);
  and (_02187_, _02177_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02188_, _01975_, _02081_);
  and (_02189_, _02188_, _02187_);
  and (_02190_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02191_, _02190_, _01978_);
  nor (_02192_, _02191_, _02189_);
  nor (_02193_, _02192_, _02179_);
  or (_02194_, _02193_, _02186_);
  and (_02195_, _01975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02196_, _02195_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_02197_, _02196_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_02198_, _02197_, _02194_);
  nor (_02199_, _02196_, _02186_);
  or (_02200_, _02199_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02201_, _02200_, _01751_);
  and (_02202_, _02201_, _02198_);
  or (_22763_, _02202_, _01750_);
  and (_02203_, _25164_, _24157_);
  and (_02204_, _02203_, _24027_);
  not (_02205_, _02203_);
  and (_02206_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_27287_, _02206_, _02204_);
  not (_02207_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_02208_, _02199_);
  nor (_02209_, _02208_, _02193_);
  nor (_02210_, _02209_, _02207_);
  or (_02211_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_02212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _02207_);
  or (_02213_, _02212_, _02199_);
  and (_02214_, _02213_, _22773_);
  and (_22764_, _02214_, _02211_);
  and (_02215_, _02203_, _23920_);
  and (_02216_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_27286_, _02216_, _02215_);
  and (_02217_, _01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_02218_, _02191_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  not (_02219_, _02179_);
  nor (_02220_, _02185_, _02219_);
  and (_02221_, _02220_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor (_02222_, _02179_, _02189_);
  or (_02223_, _02222_, _02221_);
  and (_02224_, _02223_, _02218_);
  not (_02225_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_02226_, _02199_, _02225_);
  or (_02227_, _02226_, _02224_);
  nand (_02228_, _02196_, _02225_);
  and (_02229_, _02228_, _01751_);
  and (_02230_, _02229_, _02227_);
  or (_22765_, _02230_, _02217_);
  and (_02231_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and (_02232_, _02170_, _24027_);
  or (_22766_, _02232_, _02231_);
  and (_02233_, _01876_, _24053_);
  and (_02234_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_22767_, _02234_, _02233_);
  and (_02235_, _23983_, _23892_);
  and (_02236_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_22768_, _02236_, _02235_);
  or (_02237_, _24586_, _01894_);
  or (_02238_, _23759_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_02239_, _02238_, _22773_);
  and (_26835_[2], _02239_, _02237_);
  and (_02240_, _02203_, _24053_);
  and (_02241_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_22769_, _02241_, _02240_);
  and (_02242_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  and (_02243_, _02170_, _23751_);
  or (_22770_, _02243_, _02242_);
  nor (_26868_[4], _00372_, rst);
  and (_02244_, _24145_, _23891_);
  and (_02245_, _02244_, _23751_);
  not (_02246_, _02244_);
  and (_02247_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or (_27244_, _02247_, _02245_);
  and (_02248_, _24061_, _23719_);
  and (_02249_, _02248_, _23983_);
  not (_02250_, _02248_);
  and (_02251_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or (_22771_, _02251_, _02249_);
  and (_02252_, _25169_, _24027_);
  and (_02253_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_22772_, _02253_, _02252_);
  and (_02254_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_02255_, _02170_, _24053_);
  or (_22777_, _02255_, _02254_);
  not (_02256_, _02209_);
  or (_02257_, _02256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_02258_, _02199_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02259_, _02258_, _01751_);
  and (_02260_, _02259_, _02257_);
  or (_22788_, _02260_, _01755_);
  and (_26831_[2], _24586_, _22773_);
  and (_02261_, _02185_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_02262_, _02261_, _02192_);
  or (_02263_, _02262_, _02209_);
  and (_02264_, _02263_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02265_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _02207_);
  nand (_02266_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_02267_, _02266_, _02199_);
  or (_02268_, _02267_, _02265_);
  or (_02269_, _02268_, _02264_);
  and (_22830_, _02269_, _22773_);
  nor (_02270_, _02191_, _02179_);
  or (_02271_, _02270_, _02207_);
  or (_02272_, _02271_, _02183_);
  and (_02273_, _02179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02274_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_02275_, _02274_, _22773_);
  and (_22833_, _02275_, _02272_);
  nor (_26868_[5], _00463_, rst);
  nor (_26868_[0], _00028_, rst);
  nand (_02276_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22773_);
  nor (_02277_, _02276_, _02210_);
  or (_02278_, _02262_, _02208_);
  and (_02279_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_02280_, _02279_, _02278_);
  or (_22843_, _02280_, _02277_);
  and (_02281_, _02271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_02282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_02283_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_02284_, _02283_, _02282_);
  and (_02285_, _02284_, _02273_);
  or (_02286_, _02285_, _02281_);
  and (_22847_, _02286_, _22773_);
  and (_02287_, _02203_, _23751_);
  and (_02288_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_27284_, _02288_, _02287_);
  or (_02289_, _01980_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_02290_, _01980_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_02291_, _02290_, rst);
  nand (_02292_, _02291_, _02289_);
  nor (_22893_, _02292_, _01970_);
  and (_02293_, _02282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02295_, _02293_, _02181_);
  and (_02296_, _02273_, _02295_);
  or (_02297_, _02296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not (_02298_, rxd_i);
  nand (_02300_, _02296_, _02298_);
  and (_02301_, _02300_, _22773_);
  and (_22909_, _02301_, _02297_);
  or (_02302_, _02290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_02303_, _02290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02304_, _02303_, rst);
  nand (_02305_, _02304_, _02302_);
  nor (_22916_, _02305_, _01970_);
  nor (_02306_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_02307_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_02309_, _02307_, _02306_);
  nand (_02310_, _02309_, _22773_);
  nor (_22919_, _02310_, _01970_);
  and (_02311_, _02203_, _23715_);
  and (_02312_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_22921_, _02312_, _02311_);
  and (_02313_, _23920_, _23707_);
  and (_02314_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_22925_, _02314_, _02313_);
  or (_02315_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_02316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _02207_);
  or (_02317_, _02316_, _02199_);
  and (_02318_, _02317_, _22773_);
  and (_22929_, _02318_, _02315_);
  and (_02319_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and (_02320_, _02170_, _23693_);
  or (_22934_, _02320_, _02319_);
  and (_02321_, _02203_, _23693_);
  and (_02322_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_22936_, _02322_, _02321_);
  nor (_26831_[1], _24632_, rst);
  nand (_02323_, _24537_, _23759_);
  or (_02324_, _23759_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_02325_, _02324_, _22773_);
  and (_26835_[6], _02325_, _02323_);
  and (_02326_, _24068_, _23987_);
  and (_02327_, _02326_, _23900_);
  not (_02328_, _02326_);
  and (_02329_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or (_27253_, _02329_, _02327_);
  and (_02330_, _02271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_02331_, _02293_, _02219_);
  or (_02332_, _02331_, _02330_);
  and (_02333_, _02282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02334_, _02333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02335_, _02334_, _22773_);
  and (_22985_, _02335_, _02332_);
  and (_02336_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_23001_, _02336_, _02217_);
  and (_02337_, _23719_, _23444_);
  and (_02338_, _02337_, _24053_);
  not (_02339_, _02337_);
  and (_02340_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_23018_, _02340_, _02338_);
  and (_02341_, _01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02343_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_23022_, _02343_, _02341_);
  and (_02344_, _25164_, _24123_);
  and (_02345_, _02344_, _23751_);
  not (_02346_, _02344_);
  and (_02347_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_23027_, _02347_, _02345_);
  and (_02348_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02349_, _02348_, _02265_);
  and (_23031_, _02349_, _22773_);
  and (_02350_, _25175_, _24061_);
  and (_02351_, _02350_, _23693_);
  not (_02352_, _02350_);
  and (_02353_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_23042_, _02353_, _02351_);
  nor (_26831_[0], _24561_, rst);
  and (_02354_, _02344_, _24053_);
  and (_02355_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_23049_, _02355_, _02354_);
  and (_02356_, _01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02357_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_23052_, _02357_, _02356_);
  or (_02358_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _02207_);
  or (_02360_, _02359_, _02199_);
  and (_02361_, _02360_, _22773_);
  and (_23066_, _02361_, _02358_);
  and (_02362_, _24097_, _24084_);
  not (_02363_, _02362_);
  and (_02364_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and (_02365_, _02362_, _23920_);
  or (_23072_, _02365_, _02364_);
  or (_02366_, _02256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_02367_, _02199_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02368_, _02367_, _01751_);
  and (_02369_, _02368_, _02366_);
  or (_23075_, _02369_, _01753_);
  or (_02370_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02371_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _02207_);
  or (_02372_, _02371_, _02199_);
  and (_02373_, _02372_, _22773_);
  and (_23078_, _02373_, _02370_);
  or (_02375_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02376_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _02207_);
  or (_02377_, _02376_, _02199_);
  and (_02378_, _02377_, _22773_);
  and (_23081_, _02378_, _02375_);
  and (_02379_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and (_02380_, _02362_, _23900_);
  or (_23113_, _02380_, _02379_);
  nor (_26858_[0], _26340_, rst);
  and (_02381_, _02344_, _23693_);
  and (_02382_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_23141_, _02382_, _02381_);
  and (_02383_, _02344_, _23900_);
  and (_02384_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_27262_, _02384_, _02383_);
  and (_02385_, _02344_, _23715_);
  and (_02386_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_23203_, _02386_, _02385_);
  and (_02387_, _25440_, _23983_);
  and (_02388_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or (_27208_, _02388_, _02387_);
  and (_02390_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and (_02391_, _02362_, _24027_);
  or (_23320_, _02391_, _02390_);
  and (_02392_, _25164_, _24235_);
  and (_02393_, _02392_, _23751_);
  not (_02394_, _02392_);
  and (_02395_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_23329_, _02395_, _02393_);
  and (_02396_, _02392_, _23715_);
  and (_02397_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_23334_, _02397_, _02396_);
  and (_02399_, _02392_, _23693_);
  and (_02400_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_23339_, _02400_, _02399_);
  and (_02401_, _02248_, _24027_);
  and (_02402_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or (_23358_, _02402_, _02401_);
  and (_02403_, _24235_, _23719_);
  and (_02404_, _02403_, _23920_);
  not (_02405_, _02403_);
  and (_02406_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_23369_, _02406_, _02404_);
  and (_02407_, _01709_, _23693_);
  and (_02408_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_23382_, _02408_, _02407_);
  and (_02409_, _24084_, _24068_);
  not (_02410_, _02409_);
  and (_02411_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_02412_, _02409_, _23983_);
  or (_26991_, _02412_, _02411_);
  and (_02413_, _02392_, _24027_);
  and (_02414_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_23410_, _02414_, _02413_);
  and (_02415_, _02392_, _23920_);
  and (_02416_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_27238_, _02416_, _02415_);
  and (_02417_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_02418_, _02409_, _24027_);
  or (_23430_, _02418_, _02417_);
  and (_02419_, _02392_, _23900_);
  and (_02420_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_27237_, _02420_, _02419_);
  and (_02421_, _24268_, _23715_);
  and (_02422_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or (_23438_, _02422_, _02421_);
  and (_02423_, _24123_, _23453_);
  and (_02424_, _02423_, _23900_);
  not (_02425_, _02423_);
  and (_02426_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or (_23457_, _02426_, _02424_);
  and (_02427_, _25164_, _23890_);
  and (_02428_, _02427_, _23920_);
  not (_02429_, _02427_);
  and (_02430_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_23473_, _02430_, _02428_);
  and (_02431_, _02427_, _23900_);
  and (_02432_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_23477_, _02432_, _02431_);
  and (_02434_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  and (_02435_, _02362_, _23693_);
  or (_23486_, _02435_, _02434_);
  and (_02436_, _24268_, _23693_);
  and (_02437_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or (_23491_, _02437_, _02436_);
  and (_02438_, _25954_, _22857_);
  nand (_02439_, _02438_, _23681_);
  or (_02440_, _02438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02441_, _02440_, _24330_);
  and (_02443_, _02441_, _02439_);
  or (_02444_, _25237_, _23744_);
  or (_02445_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02446_, _02445_, _22915_);
  and (_02447_, _02446_, _02444_);
  not (_02448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_02450_, _22914_, _02448_);
  or (_02451_, _02450_, rst);
  or (_02452_, _02451_, _02447_);
  or (_23500_, _02452_, _02443_);
  and (_02453_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and (_02454_, _02362_, _23751_);
  or (_26993_, _02454_, _02453_);
  and (_02455_, _24097_, _23891_);
  and (_02456_, _02455_, _24027_);
  not (_02457_, _02455_);
  and (_02458_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or (_23517_, _02458_, _02456_);
  and (_02460_, _24164_, _23983_);
  and (_02461_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_27100_, _02461_, _02460_);
  and (_02462_, _25440_, _24027_);
  and (_02463_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or (_23556_, _02463_, _02462_);
  and (_02464_, _24061_, _23909_);
  and (_02465_, _02464_, _23751_);
  not (_02466_, _02464_);
  and (_02467_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  or (_27101_, _02467_, _02465_);
  and (_02468_, _02427_, _23983_);
  and (_02469_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_23574_, _02469_, _02468_);
  and (_02470_, _02427_, _24027_);
  and (_02471_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_23592_, _02471_, _02470_);
  and (_02472_, _23907_, _22823_);
  and (_02473_, _02472_, _23251_);
  nand (_02474_, _02473_, _23357_);
  not (_02475_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_02476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_02477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_02478_, _02477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_02479_, _02478_, _02476_);
  not (_02480_, _02479_);
  and (_02481_, _02472_, _24185_);
  nor (_02482_, _02481_, _02480_);
  nor (_02483_, _02482_, _02475_);
  and (_02484_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_02485_, _02484_, _02483_);
  or (_02486_, _02485_, _02473_);
  and (_02487_, _02486_, _22773_);
  and (_23609_, _02487_, _02474_);
  and (_02488_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_02489_, _02409_, _23693_);
  or (_23619_, _02489_, _02488_);
  and (_02491_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_02492_, _02409_, _23900_);
  or (_23646_, _02492_, _02491_);
  and (_02493_, _01701_, _23900_);
  and (_02494_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or (_23674_, _02494_, _02493_);
  and (_02495_, _02427_, _23693_);
  and (_02496_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_27220_, _02496_, _02495_);
  and (_02497_, _02427_, _23751_);
  and (_02498_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_23684_, _02498_, _02497_);
  and (_02499_, _24084_, _23700_);
  not (_02500_, _02499_);
  and (_02501_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_02502_, _02499_, _23983_);
  or (_26988_, _02502_, _02501_);
  nor (_26868_[3], _00296_, rst);
  nor (_26868_[6], _00507_, rst);
  and (_02503_, _25164_, _24097_);
  and (_02504_, _02503_, _23693_);
  not (_02505_, _02503_);
  and (_02506_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_23720_, _02506_, _02504_);
  and (_02507_, _02464_, _23693_);
  and (_02508_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  or (_23762_, _02508_, _02507_);
  and (_02509_, _24108_, _23719_);
  and (_02510_, _02509_, _23920_);
  not (_02512_, _02509_);
  and (_02513_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_23773_, _02513_, _02510_);
  and (_02514_, _02464_, _23920_);
  and (_02515_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or (_23807_, _02515_, _02514_);
  and (_02516_, _25316_, _24184_);
  nand (_02517_, _02516_, _23681_);
  or (_02518_, _02516_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02519_, _02518_, _24330_);
  and (_02520_, _02519_, _02517_);
  not (_02521_, _25321_);
  or (_02522_, _02521_, _23247_);
  or (_02523_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02524_, _02523_, _22915_);
  and (_02525_, _02524_, _02522_);
  and (_02526_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_02527_, _02526_, rst);
  or (_02528_, _02527_, _02525_);
  or (_23815_, _02528_, _02520_);
  and (_02529_, _02464_, _24027_);
  and (_02530_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  or (_23826_, _02530_, _02529_);
  and (_02531_, _23930_, _23909_);
  and (_02532_, _02531_, _24053_);
  not (_02533_, _02531_);
  and (_02534_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  or (_23829_, _02534_, _02532_);
  and (_02535_, _02244_, _23920_);
  and (_02536_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or (_23834_, _02536_, _02535_);
  and (_02538_, _02244_, _23900_);
  and (_02539_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or (_23838_, _02539_, _02538_);
  nor (_02540_, _26245_, _25850_);
  nor (_02541_, _02540_, _25848_);
  nor (_02542_, _25901_, _25884_);
  nor (_02543_, _26221_, _25920_);
  and (_02544_, _02543_, _25900_);
  and (_02545_, _02544_, _02542_);
  and (_02546_, _02545_, _25883_);
  nor (_02547_, _02546_, _24647_);
  nor (_02548_, _02547_, _02541_);
  nor (_26883_, _02548_, rst);
  and (_02549_, _01856_, _25235_);
  and (_02550_, _02549_, _25673_);
  nand (_02551_, _02550_, _23976_);
  or (_02552_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02553_, _02552_, _22773_);
  and (_26845_[7], _02553_, _02551_);
  and (_02554_, _01856_, _25954_);
  not (_02555_, _02554_);
  nor (_02556_, _02555_, _23976_);
  and (_02557_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_02558_, _02557_, _25674_);
  or (_02559_, _02558_, _02556_);
  or (_02560_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02561_, _02560_, _22773_);
  and (_26846_[7], _02561_, _02559_);
  and (_02562_, _24405_, _22926_);
  and (_02564_, _01856_, _02562_);
  and (_02565_, _02564_, _25673_);
  not (_02566_, _02565_);
  nor (_02567_, _02566_, _23976_);
  and (_02568_, _02566_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_02569_, _02568_, _02567_);
  and (_26847_[7], _02569_, _22773_);
  and (_02570_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_02571_, _01860_, _23976_);
  or (_02572_, _02571_, _02570_);
  and (_26848_[7], _02572_, _22773_);
  and (_02573_, _25319_, _23450_);
  and (_02574_, _02573_, _25235_);
  and (_02575_, _02574_, _26145_);
  nor (_02576_, _25674_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_02577_, _02574_, _25673_);
  nor (_02578_, _02577_, _02576_);
  or (_02579_, _02578_, _02575_);
  or (_02580_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_02581_, _02580_, _22773_);
  and (_26849_[7], _02581_, _02579_);
  and (_02582_, _02573_, _25954_);
  and (_02583_, _02582_, _25673_);
  not (_02584_, _02583_);
  and (_02585_, _02584_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_02586_, _02584_, _23976_);
  or (_02587_, _02586_, _02585_);
  and (_26850_[7], _02587_, _22773_);
  or (_02588_, _02582_, _02574_);
  or (_02589_, _02588_, _01857_);
  nor (_02590_, _02554_, _02549_);
  not (_02591_, _02590_);
  or (_02592_, _02564_, _01857_);
  or (_02593_, _02574_, _02592_);
  nor (_02594_, _02593_, _02591_);
  not (_02595_, _02582_);
  and (_02596_, _02595_, _02594_);
  and (_02597_, _02573_, _02562_);
  not (_02598_, _02597_);
  and (_02599_, _02598_, _02596_);
  nand (_02601_, _02590_, _25673_);
  or (_02602_, _02601_, _02564_);
  or (_02603_, _02602_, _02599_);
  or (_02604_, _02603_, _02589_);
  and (_02605_, _02604_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_02606_, _02597_, _25673_);
  and (_02607_, _02606_, _26145_);
  or (_02608_, _02607_, _02605_);
  and (_26851_[7], _02608_, _22773_);
  and (_02609_, _02573_, _22927_);
  and (_02610_, _02609_, _25673_);
  not (_02611_, _02610_);
  nor (_02612_, _02611_, _23976_);
  and (_02613_, _02611_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_02614_, _02613_, _02612_);
  and (_26852_[7], _02614_, _22773_);
  and (_02615_, _02455_, _23920_);
  and (_02616_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or (_23857_, _02616_, _02615_);
  and (_02617_, _02503_, _23751_);
  and (_02618_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_23908_, _02618_, _02617_);
  and (_02619_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_02620_, _02499_, _24027_);
  or (_26987_, _02620_, _02619_);
  and (_02621_, _02503_, _24053_);
  and (_02622_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_23916_, _02622_, _02621_);
  nand (_02623_, _24186_, _23976_);
  and (_02624_, _24192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_02625_, _24975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_02626_, _25010_, _24984_);
  nor (_02627_, _02626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nor (_02628_, _02627_, _25012_);
  and (_02629_, _25001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02630_, _02629_, _25012_);
  or (_02631_, _02630_, _02628_);
  and (_02632_, _02631_, _24976_);
  nor (_02633_, _02632_, _02625_);
  nor (_02634_, _02633_, _24192_);
  or (_02636_, _02634_, _24186_);
  or (_02637_, _02636_, _02624_);
  and (_02638_, _02637_, _22773_);
  and (_23931_, _02638_, _02623_);
  and (_02639_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_02640_, _02409_, _24053_);
  or (_23947_, _02640_, _02639_);
  and (_02641_, _02503_, _23920_);
  and (_02642_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_23956_, _02642_, _02641_);
  and (_02643_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_02644_, _02409_, _23751_);
  or (_23962_, _02644_, _02643_);
  and (_02646_, _02503_, _23900_);
  and (_02647_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_24001_, _02647_, _02646_);
  and (_02648_, _02503_, _23715_);
  and (_02649_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_24007_, _02649_, _02648_);
  and (_02650_, _25164_, _24068_);
  and (_02651_, _02650_, _23920_);
  not (_02652_, _02650_);
  and (_02653_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_24070_, _02653_, _02651_);
  and (_02654_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_02655_, _02499_, _23693_);
  or (_24073_, _02655_, _02654_);
  and (_02656_, _02650_, _23900_);
  and (_02657_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_24075_, _02657_, _02656_);
  and (_02658_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_02659_, _02499_, _23900_);
  or (_24125_, _02659_, _02658_);
  and (_02660_, _02650_, _23983_);
  and (_02661_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_27178_, _02661_, _02660_);
  nor (_26868_[2], _00202_, rst);
  and (_02662_, _24084_, _23938_);
  not (_02663_, _02662_);
  and (_02664_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and (_02666_, _02662_, _23983_);
  or (_24187_, _02666_, _02664_);
  and (_02667_, _02650_, _24053_);
  and (_02668_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_24208_, _02668_, _02667_);
  and (_02669_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_02670_, _02499_, _24053_);
  or (_24256_, _02670_, _02669_);
  and (_02671_, _25159_, _24027_);
  and (_02672_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or (_24260_, _02672_, _02671_);
  and (_02674_, _02650_, _23751_);
  and (_02675_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_24291_, _02675_, _02674_);
  and (_02676_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and (_02677_, _24275_, _23751_);
  or (_24306_, _02677_, _02676_);
  and (_02679_, _25159_, _23920_);
  and (_02680_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or (_24311_, _02680_, _02679_);
  and (_02681_, _25164_, _23700_);
  and (_02682_, _02681_, _23715_);
  not (_02683_, _02681_);
  and (_02684_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_24327_, _02684_, _02682_);
  and (_02685_, _02681_, _23900_);
  and (_02686_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_24334_, _02686_, _02685_);
  nor (_26868_[1], _00120_, rst);
  and (_02687_, _24084_, _23905_);
  not (_02688_, _02687_);
  and (_02689_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_02691_, _02687_, _23983_);
  or (_24409_, _02691_, _02689_);
  and (_02693_, _02681_, _24027_);
  and (_02694_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_27062_, _02694_, _02693_);
  and (_02695_, _24098_, _23983_);
  and (_02696_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or (_24430_, _02696_, _02695_);
  nand (_02697_, _02550_, _24017_);
  or (_02699_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_24465_, _02699_, _02697_);
  nand (_02700_, _02550_, _23357_);
  or (_02701_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_24491_, _02701_, _02700_);
  not (_02702_, _02550_);
  or (_02704_, _02702_, _23205_);
  or (_02705_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_24493_, _02705_, _02704_);
  or (_02707_, _02702_, _23413_);
  or (_02708_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_24496_, _02708_, _02707_);
  and (_02709_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_02710_, _02687_, _23693_);
  or (_24499_, _02710_, _02709_);
  or (_02711_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_24547_, _02711_, _02551_);
  and (_02712_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_02714_, _02687_, _23900_);
  or (_24552_, _02714_, _02712_);
  and (_02715_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_02716_, _02687_, _23715_);
  or (_24558_, _02716_, _02715_);
  and (_02717_, _23907_, _23702_);
  and (_02718_, _02717_, _23924_);
  not (_02719_, _02718_);
  and (_02720_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  and (_02721_, _02718_, _24053_);
  or (_27161_, _02721_, _02720_);
  and (_02722_, _02717_, _24145_);
  not (_02723_, _02722_);
  and (_02724_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_02725_, _02722_, _23715_);
  or (_27160_, _02725_, _02724_);
  and (_02726_, _02717_, _24274_);
  not (_02727_, _02726_);
  and (_02728_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_02730_, _02726_, _24027_);
  or (_24584_, _02730_, _02728_);
  and (_02731_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_02732_, _02726_, _23751_);
  or (_24587_, _02732_, _02731_);
  and (_02733_, _25316_, _23250_);
  nand (_02734_, _02733_, _23681_);
  or (_02735_, _02733_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02736_, _02735_, _24330_);
  and (_02737_, _02736_, _02734_);
  or (_02738_, _02521_, _23413_);
  or (_02739_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02740_, _02739_, _22915_);
  and (_02741_, _02740_, _02738_);
  not (_02742_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_02744_, _22914_, _02742_);
  or (_02745_, _02744_, rst);
  or (_02746_, _02745_, _02741_);
  or (_24593_, _02746_, _02737_);
  and (_02748_, _02717_, _23444_);
  not (_02749_, _02748_);
  and (_02750_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  and (_02751_, _02748_, _23693_);
  or (_24600_, _02751_, _02750_);
  and (_02752_, _24084_, _23444_);
  not (_02753_, _02752_);
  and (_02754_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_02755_, _02752_, _23983_);
  or (_24607_, _02755_, _02754_);
  and (_02756_, _02717_, _24108_);
  not (_02758_, _02756_);
  and (_02759_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  and (_02760_, _02756_, _23715_);
  or (_24614_, _02760_, _02759_);
  or (_02761_, _02702_, _23744_);
  or (_02762_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_26885_, _02762_, _02761_);
  and (_02763_, _02717_, _24157_);
  not (_02764_, _02763_);
  and (_02765_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_02766_, _02763_, _23920_);
  or (_27151_, _02766_, _02765_);
  nand (_02767_, _02550_, _24047_);
  or (_02768_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_24645_, _02768_, _02767_);
  and (_02769_, _02717_, _23890_);
  not (_02771_, _02769_);
  and (_02772_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_02773_, _02769_, _23900_);
  or (_27144_, _02773_, _02772_);
  and (_02775_, _02717_, _24097_);
  not (_02776_, _02775_);
  and (_02777_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_02778_, _02775_, _23751_);
  or (_24656_, _02778_, _02777_);
  and (_02779_, _25175_, _24145_);
  and (_02780_, _02779_, _23693_);
  not (_02782_, _02779_);
  and (_02783_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_24692_, _02783_, _02780_);
  and (_02785_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_02786_, _02687_, _24053_);
  or (_24695_, _02786_, _02785_);
  and (_02789_, _25175_, _24274_);
  and (_02790_, _02789_, _23900_);
  not (_02791_, _02789_);
  and (_02792_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_24701_, _02792_, _02790_);
  and (_02794_, _25175_, _23905_);
  and (_02795_, _02794_, _24053_);
  not (_02796_, _02794_);
  and (_02797_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or (_24713_, _02797_, _02795_);
  and (_02798_, _25175_, _23930_);
  and (_02799_, _02798_, _23751_);
  not (_02800_, _02798_);
  and (_02801_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_24734_, _02801_, _02799_);
  and (_02802_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  and (_02803_, _24795_, _23983_);
  or (_24739_, _02803_, _02802_);
  and (_02805_, _25316_, _24190_);
  nand (_02807_, _02805_, _23681_);
  or (_02809_, _02805_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02810_, _02809_, _24330_);
  and (_02811_, _02810_, _02807_);
  or (_02813_, _02521_, _23205_);
  or (_02814_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02815_, _02814_, _22915_);
  and (_02816_, _02815_, _02813_);
  not (_02817_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_02818_, _22914_, _02817_);
  or (_02820_, _02818_, rst);
  or (_02821_, _02820_, _02816_);
  or (_24744_, _02821_, _02811_);
  and (_02822_, _02423_, _23715_);
  and (_02823_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or (_27201_, _02823_, _02822_);
  and (_02825_, _01709_, _23715_);
  and (_02826_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_24760_, _02826_, _02825_);
  and (_02827_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_02828_, _02752_, _24053_);
  or (_24766_, _02828_, _02827_);
  and (_02829_, _25175_, _24123_);
  and (_02831_, _02829_, _23693_);
  not (_02832_, _02829_);
  and (_02833_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or (_24771_, _02833_, _02831_);
  and (_02835_, _25176_, _23983_);
  and (_02836_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or (_24776_, _02836_, _02835_);
  and (_02838_, _02717_, _24068_);
  not (_02839_, _02838_);
  and (_02840_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  and (_02841_, _02838_, _23715_);
  or (_24780_, _02841_, _02840_);
  and (_02842_, _02717_, _23700_);
  not (_02843_, _02842_);
  and (_02844_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  and (_02845_, _02842_, _23920_);
  or (_24783_, _02845_, _02844_);
  and (_02846_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  and (_02847_, _02842_, _23751_);
  or (_24786_, _02847_, _02846_);
  and (_02848_, _02717_, _23938_);
  not (_02849_, _02848_);
  and (_02850_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_02851_, _02848_, _24053_);
  or (_24792_, _02851_, _02850_);
  and (_02853_, _25175_, _23924_);
  and (_02855_, _02853_, _24027_);
  not (_02856_, _02853_);
  and (_02857_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or (_27134_, _02857_, _02855_);
  and (_02858_, _25316_, _23208_);
  nand (_02860_, _02858_, _23681_);
  or (_02861_, _02858_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02862_, _02861_, _24330_);
  and (_02863_, _02862_, _02860_);
  nand (_02864_, _25321_, _23357_);
  or (_02865_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02866_, _02865_, _22915_);
  and (_02867_, _02866_, _02864_);
  not (_02869_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_02870_, _22914_, _02869_);
  or (_02871_, _02870_, rst);
  or (_02872_, _02871_, _02867_);
  or (_24800_, _02872_, _02863_);
  and (_02873_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and (_02874_, _24795_, _23900_);
  or (_27012_, _02874_, _02873_);
  or (_02876_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_02877_, _02876_, _22773_);
  and (_26845_[0], _02877_, _02767_);
  or (_02879_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_02880_, _02879_, _22773_);
  and (_26845_[1], _02880_, _02761_);
  or (_02882_, _02702_, _23247_);
  or (_02883_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_02884_, _02883_, _22773_);
  and (_26845_[2], _02884_, _02882_);
  or (_02885_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_02886_, _02885_, _22773_);
  and (_26845_[3], _02886_, _02707_);
  or (_02888_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_02889_, _02888_, _22773_);
  and (_26845_[4], _02889_, _02704_);
  or (_02891_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_02892_, _02891_, _22773_);
  and (_26845_[5], _02892_, _02700_);
  or (_02893_, _02550_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02894_, _02893_, _22773_);
  and (_26845_[6], _02894_, _02697_);
  and (_02895_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_02896_, _02554_, _24788_);
  or (_02897_, _02896_, _25674_);
  or (_02898_, _02897_, _02895_);
  or (_02899_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_02900_, _02899_, _22773_);
  and (_26846_[0], _02900_, _02898_);
  and (_02901_, _02554_, _23744_);
  and (_02902_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_02903_, _02902_, _25674_);
  or (_02904_, _02903_, _02901_);
  or (_02905_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_02906_, _02905_, _22773_);
  and (_26846_[1], _02906_, _02904_);
  and (_02907_, _02554_, _23247_);
  and (_02908_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_02909_, _02908_, _25674_);
  or (_02910_, _02909_, _02907_);
  or (_02911_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_02912_, _02911_, _22773_);
  and (_26846_[2], _02912_, _02910_);
  and (_02913_, _02554_, _23413_);
  and (_02914_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_02916_, _02914_, _25674_);
  or (_02917_, _02916_, _02913_);
  or (_02918_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_02919_, _02918_, _22773_);
  and (_26846_[3], _02919_, _02917_);
  and (_02920_, _02554_, _23205_);
  and (_02921_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_02922_, _02921_, _25674_);
  or (_02923_, _02922_, _02920_);
  or (_02924_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_02925_, _02924_, _22773_);
  and (_26846_[4], _02925_, _02923_);
  nor (_02926_, _02555_, _23357_);
  and (_02927_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_02928_, _02927_, _25674_);
  or (_02929_, _02928_, _02926_);
  or (_02930_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_02931_, _02930_, _22773_);
  and (_26846_[5], _02931_, _02929_);
  nor (_02932_, _02555_, _24017_);
  and (_02933_, _02555_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_02934_, _02933_, _25674_);
  or (_02935_, _02934_, _02932_);
  or (_02936_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_02937_, _02936_, _22773_);
  and (_26846_[6], _02937_, _02935_);
  nand (_02938_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_02939_, _02938_, _02590_);
  nor (_02940_, _02564_, _02591_);
  or (_02941_, _02940_, _25674_);
  and (_02942_, _02941_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_02943_, _02565_, _24788_);
  or (_02944_, _02943_, _02942_);
  or (_02945_, _02944_, _02939_);
  and (_26847_[0], _02945_, _22773_);
  and (_02947_, _02565_, _23744_);
  and (_02949_, _02566_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_02950_, _02949_, _02947_);
  and (_26847_[1], _02950_, _22773_);
  and (_02951_, _02566_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_02952_, _02565_, _23247_);
  or (_02953_, _02952_, _02951_);
  and (_26847_[2], _02953_, _22773_);
  and (_02954_, _02565_, _23413_);
  and (_02956_, _02566_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_02957_, _02956_, _02954_);
  and (_26847_[3], _02957_, _22773_);
  and (_02958_, _02565_, _23205_);
  and (_02959_, _02566_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_02960_, _02959_, _02958_);
  and (_26847_[4], _02960_, _22773_);
  nor (_02962_, _02566_, _23357_);
  and (_02963_, _02566_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_02964_, _02963_, _02962_);
  and (_26847_[5], _02964_, _22773_);
  nor (_02966_, _02566_, _24017_);
  and (_02967_, _02566_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_02968_, _02967_, _02966_);
  and (_26847_[6], _02968_, _22773_);
  and (_02970_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_02971_, _02970_, _01864_);
  and (_26848_[0], _02971_, _22773_);
  and (_02973_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_02974_, _02973_, _01862_);
  and (_26848_[1], _02974_, _22773_);
  and (_02975_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_02976_, _02975_, _01859_);
  and (_26848_[2], _02976_, _22773_);
  and (_02977_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_02978_, _02977_, _01874_);
  and (_26848_[3], _02978_, _22773_);
  and (_02980_, _01858_, _23205_);
  and (_02981_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_02982_, _02981_, _02980_);
  and (_26848_[4], _02982_, _22773_);
  nor (_02983_, _01860_, _23357_);
  and (_02984_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_02985_, _02984_, _02983_);
  and (_26848_[5], _02985_, _22773_);
  nor (_02986_, _01860_, _24017_);
  and (_02988_, _01860_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_02989_, _02988_, _02986_);
  and (_26848_[6], _02989_, _22773_);
  or (_02991_, _02594_, _25674_);
  and (_02992_, _02991_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_02994_, _02592_, _02591_);
  nand (_02995_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_02996_, _02995_, _02994_);
  and (_02997_, _02577_, _24788_);
  or (_02998_, _02997_, _02996_);
  or (_02999_, _02998_, _02992_);
  and (_26849_[0], _02999_, _22773_);
  or (_03000_, _02991_, _02549_);
  and (_03001_, _03000_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or (_03002_, _02592_, _02554_);
  and (_03003_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_03004_, _03003_, _03002_);
  and (_03005_, _02577_, _23744_);
  or (_03006_, _03005_, _03004_);
  or (_03007_, _03006_, _03001_);
  and (_26849_[1], _03007_, _22773_);
  and (_03008_, _02577_, _23247_);
  and (_03009_, _03000_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_03010_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_03011_, _03010_, _03002_);
  or (_03012_, _03011_, _03009_);
  or (_03013_, _03012_, _03008_);
  and (_26849_[2], _03013_, _22773_);
  and (_03014_, _02577_, _23413_);
  and (_03015_, _03000_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03016_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03017_, _03016_, _03002_);
  or (_03018_, _03017_, _03015_);
  or (_03019_, _03018_, _03014_);
  and (_26849_[3], _03019_, _22773_);
  and (_03020_, _02577_, _23205_);
  and (_03021_, _03000_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03022_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03023_, _03022_, _03002_);
  or (_03024_, _03023_, _03021_);
  or (_03025_, _03024_, _03020_);
  and (_26849_[4], _03025_, _22773_);
  and (_03026_, _02577_, _25813_);
  and (_03027_, _03000_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_03028_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_03029_, _03028_, _03002_);
  or (_03030_, _03029_, _03027_);
  or (_03031_, _03030_, _03026_);
  and (_26849_[5], _03031_, _22773_);
  and (_03032_, _02577_, _25833_);
  not (_03033_, _02994_);
  or (_03034_, _02991_, _03033_);
  and (_03035_, _03034_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_03036_, _03035_, _03032_);
  and (_26849_[6], _03036_, _22773_);
  and (_03037_, _02593_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_03038_, _03037_, _25673_);
  or (_03039_, _02601_, _02596_);
  and (_03040_, _03039_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_03042_, _02583_, _24788_);
  or (_03043_, _03042_, _03040_);
  or (_03044_, _03043_, _03038_);
  and (_26850_[0], _03044_, _22773_);
  and (_03046_, _03039_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_03047_, _02583_, _23744_);
  and (_03048_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_03049_, _03048_, _02593_);
  or (_03050_, _03049_, _03047_);
  or (_03051_, _03050_, _03046_);
  and (_26850_[1], _03051_, _22773_);
  and (_03052_, _02584_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_03053_, _02583_, _23247_);
  or (_03054_, _03053_, _03052_);
  and (_26850_[2], _03054_, _22773_);
  and (_03055_, _02583_, _23413_);
  and (_03056_, _03039_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_03057_, _02593_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_03058_, _03057_, _25673_);
  or (_03059_, _03058_, _03056_);
  or (_03060_, _03059_, _03055_);
  and (_26850_[3], _03060_, _22773_);
  and (_03061_, _02584_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_03062_, _02583_, _23205_);
  or (_03063_, _03062_, _03061_);
  and (_26850_[4], _03063_, _22773_);
  and (_03064_, _02584_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_03065_, _02584_, _23357_);
  or (_03066_, _03065_, _03064_);
  and (_26850_[5], _03066_, _22773_);
  and (_03067_, _02584_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_03068_, _02584_, _24017_);
  or (_03069_, _03068_, _03067_);
  and (_26850_[6], _03069_, _22773_);
  and (_03070_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_03071_, _03070_, _02589_);
  and (_03072_, _02603_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_03073_, _02606_, _24788_);
  or (_03074_, _03073_, _03072_);
  or (_03075_, _03074_, _03071_);
  and (_26851_[0], _03075_, _22773_);
  and (_03076_, _02603_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_03077_, _02606_, _23744_);
  and (_03078_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_03079_, _03078_, _02589_);
  or (_03080_, _03079_, _03077_);
  or (_03082_, _03080_, _03076_);
  and (_26851_[1], _03082_, _22773_);
  and (_03083_, _02603_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_03084_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_03085_, _03084_, _02589_);
  and (_03086_, _02606_, _23247_);
  or (_03087_, _03086_, _03085_);
  or (_03088_, _03087_, _03083_);
  and (_26851_[2], _03088_, _22773_);
  and (_03089_, _02603_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_03090_, _02606_, _23413_);
  and (_03091_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_03092_, _03091_, _02589_);
  or (_03093_, _03092_, _03090_);
  or (_03094_, _03093_, _03089_);
  and (_26851_[3], _03094_, _22773_);
  and (_03095_, _02603_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_03096_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_03097_, _03096_, _02589_);
  and (_03098_, _02606_, _23205_);
  or (_03099_, _03098_, _03097_);
  or (_03100_, _03099_, _03095_);
  and (_26851_[4], _03100_, _22773_);
  and (_03101_, _02606_, _25813_);
  and (_03102_, _02603_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_03103_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_03104_, _03103_, _02589_);
  or (_03105_, _03104_, _03102_);
  or (_03106_, _03105_, _03101_);
  and (_26851_[5], _03106_, _22773_);
  and (_03107_, _02606_, _25833_);
  and (_03108_, _02589_, _25673_);
  or (_03109_, _03108_, _02603_);
  and (_03110_, _03109_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_03111_, _03110_, _03107_);
  and (_26851_[6], _03111_, _22773_);
  and (_03112_, _02609_, _24788_);
  and (_03113_, _02611_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_03114_, _03113_, _03112_);
  or (_03115_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03116_, _03115_, _22773_);
  and (_26852_[0], _03116_, _03114_);
  not (_03117_, _02609_);
  and (_03118_, _03117_, _02599_);
  or (_03119_, _02601_, _02592_);
  or (_03120_, _03119_, _03118_);
  and (_03121_, _03120_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_03122_, _02610_, _23744_);
  or (_03123_, _02597_, _02588_);
  and (_03124_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_03125_, _03124_, _03123_);
  or (_03126_, _03125_, _03122_);
  or (_03127_, _03126_, _03121_);
  and (_26852_[1], _03127_, _22773_);
  and (_03128_, _02611_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_03130_, _02610_, _23247_);
  or (_03131_, _03130_, _03128_);
  and (_26852_[2], _03131_, _22773_);
  and (_03132_, _03120_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_03133_, _02610_, _23413_);
  and (_03134_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_03135_, _03134_, _03123_);
  or (_03136_, _03135_, _03133_);
  or (_03137_, _03136_, _03132_);
  and (_26852_[3], _03137_, _22773_);
  and (_03138_, _03120_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_03139_, _02610_, _23205_);
  and (_03140_, _25673_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_03141_, _03140_, _03123_);
  or (_03142_, _03141_, _03139_);
  or (_03143_, _03142_, _03138_);
  and (_26852_[4], _03143_, _22773_);
  and (_03145_, _02611_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_03146_, _02611_, _23357_);
  or (_03147_, _03146_, _03145_);
  and (_26852_[5], _03147_, _22773_);
  and (_03148_, _02611_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_03149_, _02611_, _24017_);
  or (_03150_, _03149_, _03148_);
  and (_26852_[6], _03150_, _22773_);
  and (_03151_, _02244_, _23715_);
  and (_03152_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or (_25070_, _03152_, _03151_);
  and (_03153_, _02455_, _23900_);
  and (_03154_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or (_25073_, _03154_, _03153_);
  and (_03155_, _25176_, _23920_);
  and (_03156_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or (_25130_, _03156_, _03155_);
  and (_03157_, _02717_, _23905_);
  not (_03158_, _03157_);
  and (_03159_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  and (_03160_, _03157_, _23751_);
  or (_25286_, _03160_, _03159_);
  and (_03161_, _02717_, _23930_);
  not (_03162_, _03161_);
  and (_03163_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_03164_, _03161_, _23715_);
  or (_25296_, _03164_, _03163_);
  and (_03165_, _02717_, _24123_);
  not (_03166_, _03165_);
  and (_03167_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  and (_03168_, _03165_, _23983_);
  or (_27148_, _03168_, _03167_);
  and (_03169_, _02717_, _24235_);
  not (_03170_, _03169_);
  and (_03171_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and (_03172_, _03169_, _23751_);
  or (_27146_, _03172_, _03171_);
  and (_03173_, _24901_, _23751_);
  and (_03174_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_27043_, _03174_, _03173_);
  and (_03175_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_03176_, _02775_, _23983_);
  or (_25366_, _03176_, _03175_);
  and (_03178_, _02853_, _23751_);
  and (_03179_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or (_25371_, _03179_, _03178_);
  and (_03180_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and (_03181_, _24795_, _24027_);
  or (_25377_, _03181_, _03180_);
  and (_03182_, _02798_, _24027_);
  and (_03183_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_25391_, _03183_, _03182_);
  not (_03184_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03185_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_03186_, _03185_, _03184_);
  and (_03188_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _22773_);
  and (_27322_, _03188_, _03186_);
  nor (_03189_, _03186_, rst);
  nand (_03190_, _03185_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03191_, _03185_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03192_, _03191_, _03190_);
  and (_27323_[3], _03192_, _03189_);
  not (_03194_, _26041_);
  nor (_03195_, _26112_, _03194_);
  not (_03196_, _26153_);
  nor (_03197_, _03196_, _26013_);
  and (_03198_, _03197_, _26076_);
  and (_03199_, _03198_, _03195_);
  not (_03201_, _26271_);
  and (_03202_, _00352_, _03201_);
  nor (_03203_, _24190_, _23055_);
  or (_03204_, _03203_, _24431_);
  and (_03205_, _26275_, _26272_);
  and (_03206_, _03205_, _03204_);
  and (_03207_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03208_, _03207_, _26264_);
  or (_03209_, _03208_, _03206_);
  or (_03210_, _03209_, _03202_);
  or (_03211_, _00958_, _26265_);
  and (_03212_, _03211_, _03210_);
  and (_03213_, _00443_, _03201_);
  nand (_03214_, _23681_, _23208_);
  or (_03215_, _23208_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03216_, _03215_, _03205_);
  and (_03217_, _03216_, _03214_);
  and (_03218_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03219_, _03218_, _26264_);
  or (_03220_, _03219_, _03217_);
  or (_03221_, _03220_, _03213_);
  or (_03222_, _01021_, _26265_);
  and (_03223_, _03222_, _03221_);
  or (_03224_, _03223_, _03212_);
  nand (_03225_, _03223_, _03212_);
  nand (_03226_, _03225_, _03224_);
  nand (_03227_, _00564_, _03201_);
  not (_03228_, _03205_);
  not (_03229_, _24373_);
  nor (_03230_, _03229_, _23681_);
  nor (_03231_, _24373_, _23514_);
  nor (_03232_, _03231_, _03230_);
  nor (_03233_, _03232_, _03228_);
  and (_03234_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03235_, _03234_, _26264_);
  nor (_03236_, _03235_, _03233_);
  nand (_03237_, _03236_, _03227_);
  or (_03238_, _01086_, _26265_);
  and (_03239_, _03238_, _03237_);
  nand (_03240_, _00619_, _03201_);
  not (_03241_, _24341_);
  nor (_03242_, _03241_, _23681_);
  nor (_03243_, _24341_, _23482_);
  nor (_03244_, _03243_, _03242_);
  nor (_03246_, _03244_, _03228_);
  and (_03247_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03249_, _03247_, _26264_);
  nor (_03250_, _03249_, _03246_);
  nand (_03251_, _03250_, _03240_);
  and (_03252_, _23487_, _23173_);
  and (_03253_, _23635_, _23152_);
  nor (_03255_, _01065_, _24002_);
  not (_03256_, _03255_);
  nor (_03258_, _03256_, _01058_);
  and (_03259_, _03258_, _23485_);
  nor (_03260_, _03258_, _23485_);
  or (_03261_, _03260_, _03259_);
  and (_03262_, _03261_, _23067_);
  and (_03263_, _23487_, _23046_);
  nor (_03265_, _03263_, _23658_);
  nor (_03267_, _03265_, _23316_);
  or (_03268_, _03267_, _03262_);
  or (_03270_, _03268_, _03253_);
  and (_03271_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_03273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_03274_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_03275_, _03274_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_03276_, _03275_, _03273_);
  nor (_03277_, _03276_, _01076_);
  and (_03278_, _03276_, _01076_);
  or (_03279_, _03278_, _23598_);
  or (_03280_, _03279_, _03277_);
  and (_03282_, _26756_, _26716_);
  not (_03283_, _03282_);
  and (_03285_, _03283_, _26757_);
  and (_03287_, _03285_, _26607_);
  not (_03288_, _03287_);
  nand (_03289_, _03288_, _03280_);
  or (_03290_, _03289_, _03271_);
  or (_03292_, _03290_, _03270_);
  or (_03293_, _03292_, _03252_);
  or (_03294_, _03293_, _26265_);
  and (_03295_, _03294_, _03251_);
  or (_03296_, _03295_, _03239_);
  nand (_03297_, _03295_, _03239_);
  and (_03298_, _03297_, _03296_);
  nand (_03299_, _03298_, _03226_);
  or (_03300_, _03298_, _03226_);
  nand (_03301_, _03300_, _03299_);
  nand (_03302_, _26798_, _03201_);
  nor (_03303_, _24405_, _23551_);
  nor (_03305_, _03303_, _02080_);
  nor (_03306_, _03305_, _03228_);
  and (_03307_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03309_, _03307_, _26264_);
  nor (_03310_, _03309_, _03306_);
  nand (_03311_, _03310_, _03302_);
  or (_03312_, _00691_, _26265_);
  and (_03313_, _03312_, _03311_);
  nand (_03314_, _00101_, _03201_);
  nor (_03315_, _22895_, _23542_);
  nor (_03316_, _03315_, _02150_);
  nor (_03318_, _03316_, _03228_);
  and (_03319_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03321_, _03319_, _26264_);
  nor (_03322_, _03321_, _03318_);
  nand (_03323_, _03322_, _03314_);
  and (_03324_, _00747_, _26264_);
  not (_03325_, _03324_);
  and (_03326_, _03325_, _03323_);
  or (_03327_, _03326_, _03313_);
  nand (_03329_, _03326_, _03313_);
  nand (_03330_, _03329_, _03327_);
  nand (_03331_, _00183_, _03201_);
  nor (_03332_, _24184_, _23214_);
  nor (_03333_, _03332_, _02023_);
  nor (_03334_, _03333_, _03228_);
  and (_03335_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03336_, _03335_, _26264_);
  nor (_03337_, _03336_, _03334_);
  nand (_03338_, _03337_, _03331_);
  and (_03339_, _00815_, _26264_);
  not (_03340_, _03339_);
  and (_03341_, _03340_, _03338_);
  nand (_03342_, _00277_, _03201_);
  nor (_03343_, _23250_, _23385_);
  nor (_03344_, _03343_, _24323_);
  nor (_03345_, _03344_, _03228_);
  and (_03346_, _26277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_03347_, _03346_, _26264_);
  not (_03349_, _03347_);
  nor (_03350_, _03349_, _03345_);
  nand (_03351_, _03350_, _03342_);
  and (_03352_, _00878_, _26264_);
  not (_03353_, _03352_);
  nand (_03354_, _03353_, _03351_);
  nand (_03355_, _03354_, _03341_);
  or (_03356_, _03354_, _03341_);
  and (_03357_, _03356_, _03355_);
  nand (_03358_, _03357_, _03330_);
  or (_03359_, _03357_, _03330_);
  nand (_03360_, _03359_, _03358_);
  nand (_03361_, _03360_, _03301_);
  or (_03362_, _03360_, _03301_);
  and (_03363_, _03362_, _03361_);
  nand (_03364_, _03363_, _26365_);
  and (_03365_, _26345_, _26312_);
  or (_03366_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03367_, _03366_, _03365_);
  and (_03368_, _03367_, _03364_);
  not (_03369_, _26365_);
  not (_03370_, _26345_);
  and (_03371_, _03370_, _26312_);
  and (_03373_, _03371_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_03374_, _03370_, _26312_);
  and (_03375_, _03374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_03376_, _03375_, _03373_);
  and (_03377_, _03376_, _03369_);
  nor (_03378_, _26345_, _26312_);
  and (_03379_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  not (_03380_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_03382_, _26365_, _03380_);
  or (_03383_, _03382_, _03379_);
  and (_03384_, _03383_, _03378_);
  and (_03385_, _03371_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03386_, _03374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03387_, _03386_, _03385_);
  and (_03388_, _03387_, _26365_);
  or (_03389_, _03388_, _03384_);
  or (_03390_, _03389_, _03377_);
  or (_03391_, _03390_, _03368_);
  and (_03392_, _03391_, _03199_);
  not (_03393_, _26076_);
  and (_03394_, _26153_, _26013_);
  and (_03395_, _03394_, _03195_);
  and (_03396_, _03395_, _03393_);
  and (_03397_, _03374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_03398_, _03365_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_03399_, _03398_, _03397_);
  and (_03400_, _03399_, _03369_);
  and (_03401_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_03402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_03403_, _26365_, _03402_);
  or (_03404_, _03403_, _03401_);
  and (_03405_, _03404_, _03371_);
  and (_03406_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03407_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_03408_, _03407_, _03406_);
  and (_03410_, _03408_, _03378_);
  or (_03411_, _03410_, _03405_);
  and (_03413_, _03374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_03414_, _03365_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_03415_, _03414_, _03413_);
  and (_03416_, _03415_, _26365_);
  or (_03417_, _03416_, _03411_);
  or (_03418_, _03417_, _03400_);
  and (_03419_, _03418_, _03396_);
  nand (_03420_, _26153_, _26112_);
  or (_03421_, _03420_, _26076_);
  not (_03422_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_03423_, _03198_, _03422_);
  and (_03424_, _03423_, _03421_);
  not (_03425_, _03195_);
  and (_03426_, _03394_, _26076_);
  and (_03427_, _03426_, _03425_);
  nor (_03428_, _03427_, _03396_);
  and (_03429_, _03428_, _03424_);
  nor (_03430_, _26112_, _26041_);
  and (_03431_, _03430_, _03426_);
  and (_03432_, _03378_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03433_, _03371_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03435_, _03433_, _03432_);
  and (_03436_, _03435_, _03369_);
  and (_03438_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_03440_, _26365_, _23055_);
  or (_03441_, _03440_, _03438_);
  and (_03442_, _03441_, _03365_);
  nor (_03443_, _26365_, _23514_);
  and (_03444_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03445_, _03444_, _03443_);
  and (_03446_, _03445_, _03374_);
  or (_03447_, _03446_, _03442_);
  and (_03448_, _03378_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03449_, _03371_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03450_, _03449_, _03448_);
  and (_03451_, _03450_, _26365_);
  or (_03452_, _03451_, _03447_);
  or (_03453_, _03452_, _03436_);
  and (_03454_, _03453_, _03431_);
  or (_03455_, _03454_, _03429_);
  or (_03456_, _03455_, _03419_);
  and (_03458_, _26374_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_03459_, _26112_, _26041_);
  and (_03460_, _03197_, _03393_);
  and (_03461_, _03460_, _03459_);
  and (_03462_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_03463_, _26365_, _01969_);
  or (_03465_, _03463_, _03462_);
  and (_03466_, _03465_, _03378_);
  nor (_03467_, _26365_, _01967_);
  and (_03468_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03469_, _03468_, _03467_);
  and (_03471_, _03469_, _03374_);
  or (_03473_, _03471_, _03466_);
  and (_03474_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  not (_03476_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_03477_, _26365_, _03476_);
  or (_03478_, _03477_, _03474_);
  and (_03479_, _03478_, _03365_);
  and (_03481_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_03482_, _26365_, _02085_);
  or (_03483_, _03482_, _03481_);
  and (_03484_, _03483_, _03371_);
  or (_03485_, _03484_, _03479_);
  or (_03486_, _03485_, _03473_);
  and (_03487_, _03486_, _03461_);
  and (_03488_, _26112_, _03194_);
  and (_03489_, _03488_, _03460_);
  and (_03490_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_03491_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03492_, _03491_, _03490_);
  and (_03493_, _03492_, _03378_);
  and (_03494_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03495_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03496_, _03495_, _03494_);
  and (_03497_, _03496_, _03374_);
  or (_03498_, _03497_, _03493_);
  and (_03499_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_03500_, _26365_, _24825_);
  or (_03501_, _03500_, _03499_);
  and (_03502_, _03501_, _03365_);
  and (_03503_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_03504_, _26365_, _24830_);
  or (_03506_, _03504_, _03503_);
  and (_03507_, _03506_, _03371_);
  or (_03508_, _03507_, _03502_);
  or (_03509_, _03508_, _03498_);
  and (_03510_, _03509_, _03489_);
  and (_03511_, _03430_, _03198_);
  and (_03512_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_03513_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_03514_, _26365_, _03513_);
  or (_03515_, _03514_, _03512_);
  and (_03516_, _03515_, _03378_);
  not (_03517_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_03518_, _26365_, _03517_);
  and (_03520_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03521_, _03520_, _03518_);
  and (_03522_, _03521_, _03374_);
  or (_03523_, _03522_, _03516_);
  and (_03524_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_03525_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_03526_, _26365_, _03525_);
  or (_03527_, _03526_, _03524_);
  and (_03528_, _03527_, _03365_);
  and (_03529_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_03530_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_03531_, _26365_, _03530_);
  or (_03532_, _03531_, _03529_);
  and (_03533_, _03532_, _03371_);
  or (_03534_, _03533_, _03528_);
  or (_03535_, _03534_, _03523_);
  and (_03537_, _03535_, _03511_);
  or (_03538_, _03537_, _03510_);
  or (_03539_, _03538_, _03487_);
  or (_03540_, _03539_, _03458_);
  or (_03541_, _03540_, _03456_);
  and (_03543_, _03394_, _03393_);
  and (_03544_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_03546_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_03547_, _03546_, _03544_);
  and (_03548_, _03547_, _03365_);
  or (_03549_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03550_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03551_, _03550_, _03378_);
  and (_03552_, _03551_, _03549_);
  or (_03554_, _03552_, _03548_);
  and (_03555_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_03556_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03557_, _03556_, _03555_);
  and (_03558_, _03557_, _03371_);
  or (_03559_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03560_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03561_, _03560_, _03374_);
  and (_03562_, _03561_, _03559_);
  or (_03563_, _03562_, _03558_);
  or (_03564_, _03563_, _03554_);
  and (_03565_, _03564_, _03459_);
  and (_03566_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03567_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03568_, _03567_, _03566_);
  and (_03569_, _03568_, _03378_);
  or (_03570_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_03571_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_03572_, _03571_, _03365_);
  and (_03573_, _03572_, _03570_);
  or (_03574_, _03573_, _03569_);
  and (_03576_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03578_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03580_, _03578_, _03576_);
  and (_03582_, _03580_, _03374_);
  or (_03583_, _26365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_03584_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03585_, _03584_, _03371_);
  and (_03586_, _03585_, _03583_);
  or (_03587_, _03586_, _03582_);
  or (_03588_, _03587_, _03574_);
  and (_03589_, _03588_, _03488_);
  or (_03590_, _03589_, _03565_);
  and (_03592_, _03590_, _03543_);
  not (_03593_, _25903_);
  and (_03594_, _26228_, _24704_);
  nor (_03595_, _03594_, _03593_);
  and (_03596_, _25924_, _24681_);
  and (_03597_, _24704_, _24690_);
  nor (_03598_, _03597_, _03596_);
  nor (_03599_, _26232_, _25931_);
  and (_03600_, _03599_, _03598_);
  nor (_03601_, _24522_, _24503_);
  and (_03602_, _03601_, _24615_);
  or (_03603_, _03602_, _25913_);
  nor (_03604_, _03603_, _25899_);
  and (_03605_, _24690_, _24670_);
  and (_03606_, _03605_, _24680_);
  or (_03607_, _25905_, _24725_);
  nor (_03608_, _03607_, _03606_);
  and (_03609_, _03608_, _03604_);
  and (_03610_, _03609_, _03600_);
  and (_03611_, _03610_, _03595_);
  and (_03612_, _03611_, _25896_);
  nor (_03613_, _03612_, _24647_);
  nor (_03614_, _03613_, p3_in[4]);
  not (_03615_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03616_, _03613_, _03615_);
  nor (_03617_, _03616_, _03614_);
  and (_03618_, _03617_, _03369_);
  nor (_03619_, _03613_, p3_in[0]);
  not (_03620_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_03621_, _03613_, _03620_);
  nor (_03622_, _03621_, _03619_);
  and (_03623_, _03622_, _26365_);
  or (_03624_, _03623_, _03618_);
  and (_03625_, _03624_, _03365_);
  nor (_03626_, _03613_, p3_in[3]);
  not (_03627_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03628_, _03613_, _03627_);
  nor (_03629_, _03628_, _03626_);
  or (_03630_, _03629_, _03369_);
  or (_03631_, _03613_, p3_in[7]);
  not (_03632_, _03613_);
  or (_03633_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03634_, _03633_, _03631_);
  or (_03635_, _03634_, _26365_);
  and (_03636_, _03635_, _03378_);
  and (_03637_, _03636_, _03630_);
  or (_03638_, _03637_, _03625_);
  nor (_03639_, _03613_, p3_in[5]);
  not (_03640_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03641_, _03613_, _03640_);
  nor (_03642_, _03641_, _03639_);
  and (_03643_, _03642_, _03369_);
  nor (_03644_, _03613_, p3_in[1]);
  not (_03645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03646_, _03613_, _03645_);
  nor (_03647_, _03646_, _03644_);
  and (_03648_, _03647_, _26365_);
  or (_03649_, _03648_, _03643_);
  and (_03650_, _03649_, _03371_);
  or (_03651_, _03613_, p3_in[2]);
  or (_03652_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03653_, _03652_, _03651_);
  or (_03654_, _03653_, _03369_);
  or (_03655_, _03613_, p3_in[6]);
  or (_03656_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03657_, _03656_, _03655_);
  or (_03658_, _03657_, _26365_);
  and (_03659_, _03658_, _03374_);
  and (_03660_, _03659_, _03654_);
  or (_03661_, _03660_, _03650_);
  or (_03662_, _03661_, _03638_);
  and (_03664_, _03662_, _03198_);
  nor (_03665_, _03613_, p2_in[4]);
  not (_03666_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03667_, _03613_, _03666_);
  nor (_03668_, _03667_, _03665_);
  and (_03669_, _03668_, _03369_);
  nor (_03670_, _03613_, p2_in[0]);
  not (_03671_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_03672_, _03613_, _03671_);
  nor (_03673_, _03672_, _03670_);
  and (_03674_, _03673_, _26365_);
  or (_03675_, _03674_, _03669_);
  and (_03676_, _03675_, _03365_);
  nor (_03677_, _03613_, p2_in[3]);
  not (_03679_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03680_, _03613_, _03679_);
  nor (_03681_, _03680_, _03677_);
  or (_03682_, _03681_, _03369_);
  or (_03683_, _03613_, p2_in[7]);
  or (_03684_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03685_, _03684_, _03683_);
  or (_03686_, _03685_, _26365_);
  and (_03687_, _03686_, _03378_);
  and (_03688_, _03687_, _03682_);
  or (_03689_, _03688_, _03676_);
  nor (_03690_, _03613_, p2_in[5]);
  not (_03692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03694_, _03613_, _03692_);
  nor (_03695_, _03694_, _03690_);
  and (_03696_, _03695_, _03369_);
  nor (_03697_, _03613_, p2_in[1]);
  not (_03698_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03699_, _03613_, _03698_);
  nor (_03700_, _03699_, _03697_);
  and (_03701_, _03700_, _26365_);
  or (_03702_, _03701_, _03696_);
  and (_03703_, _03702_, _03371_);
  or (_03704_, _03613_, p2_in[2]);
  or (_03705_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03706_, _03705_, _03704_);
  or (_03707_, _03706_, _03369_);
  or (_03708_, _03613_, p2_in[6]);
  or (_03709_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03710_, _03709_, _03708_);
  or (_03711_, _03710_, _26365_);
  and (_03712_, _03711_, _03374_);
  and (_03713_, _03712_, _03707_);
  or (_03714_, _03713_, _03703_);
  or (_03715_, _03714_, _03689_);
  and (_03716_, _03715_, _03426_);
  or (_03717_, _03716_, _03664_);
  and (_03718_, _03717_, _03488_);
  nor (_03719_, _03613_, p1_in[4]);
  and (_03720_, _03613_, _02817_);
  nor (_03721_, _03720_, _03719_);
  and (_03723_, _03721_, _03369_);
  nor (_03724_, _03613_, p1_in[0]);
  and (_03725_, _03613_, _25328_);
  nor (_03727_, _03725_, _03724_);
  and (_03728_, _03727_, _26365_);
  or (_03730_, _03728_, _03723_);
  and (_03731_, _03730_, _03365_);
  nor (_03732_, _03613_, p1_in[3]);
  and (_03733_, _03613_, _02742_);
  nor (_03734_, _03733_, _03732_);
  or (_03735_, _03734_, _03369_);
  or (_03736_, _03613_, p1_in[7]);
  or (_03737_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03738_, _03737_, _03736_);
  or (_03739_, _03738_, _26365_);
  and (_03740_, _03739_, _03378_);
  and (_03741_, _03740_, _03735_);
  or (_03742_, _03741_, _03731_);
  nor (_03743_, _03613_, p1_in[5]);
  and (_03745_, _03613_, _02869_);
  nor (_03746_, _03745_, _03743_);
  and (_03747_, _03746_, _03369_);
  nor (_03748_, _03613_, p1_in[1]);
  not (_03749_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03750_, _03613_, _03749_);
  nor (_03751_, _03750_, _03748_);
  and (_03752_, _03751_, _26365_);
  or (_03753_, _03752_, _03747_);
  and (_03754_, _03753_, _03371_);
  or (_03755_, _03613_, p1_in[2]);
  or (_03756_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03757_, _03756_, _03755_);
  or (_03758_, _03757_, _03369_);
  or (_03759_, _03613_, p1_in[6]);
  or (_03760_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03761_, _03760_, _03759_);
  or (_03762_, _03761_, _26365_);
  and (_03763_, _03762_, _03374_);
  and (_03764_, _03763_, _03758_);
  or (_03765_, _03764_, _03754_);
  or (_03766_, _03765_, _03742_);
  and (_03767_, _03766_, _03198_);
  nor (_03768_, _03613_, p0_in[4]);
  and (_03769_, _03613_, _25287_);
  nor (_03770_, _03769_, _03768_);
  and (_03771_, _03770_, _03369_);
  nor (_03772_, _03613_, p0_in[0]);
  not (_03773_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_03774_, _03613_, _03773_);
  nor (_03775_, _03774_, _03772_);
  and (_03776_, _03775_, _26365_);
  or (_03777_, _03776_, _03771_);
  and (_03778_, _03777_, _03365_);
  nor (_03779_, _03613_, p0_in[3]);
  and (_03780_, _03613_, _25242_);
  nor (_03781_, _03780_, _03779_);
  or (_03782_, _03781_, _03369_);
  or (_03783_, _03613_, p0_in[7]);
  or (_03784_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03785_, _03784_, _03783_);
  or (_03786_, _03785_, _26365_);
  and (_03787_, _03786_, _03378_);
  and (_03788_, _03787_, _03782_);
  or (_03789_, _03788_, _03778_);
  nor (_03790_, _03613_, p0_in[5]);
  and (_03791_, _03613_, _25270_);
  nor (_03792_, _03791_, _03790_);
  and (_03793_, _03792_, _03369_);
  nor (_03794_, _03613_, p0_in[1]);
  and (_03795_, _03613_, _02448_);
  nor (_03796_, _03795_, _03794_);
  and (_03797_, _03796_, _26365_);
  or (_03798_, _03797_, _03793_);
  and (_03800_, _03798_, _03371_);
  or (_03801_, _03613_, p0_in[2]);
  or (_03802_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03803_, _03802_, _03801_);
  or (_03804_, _03803_, _03369_);
  or (_03805_, _03613_, p0_in[6]);
  or (_03806_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03807_, _03806_, _03805_);
  or (_03808_, _03807_, _26365_);
  and (_03809_, _03808_, _03374_);
  and (_03810_, _03809_, _03804_);
  or (_03811_, _03810_, _03800_);
  or (_03812_, _03811_, _03789_);
  and (_03813_, _03812_, _03426_);
  or (_03814_, _03813_, _03767_);
  and (_03815_, _03814_, _03459_);
  or (_03816_, _03815_, _03718_);
  or (_03817_, _03816_, _03592_);
  or (_03818_, _03817_, _03541_);
  or (_03819_, _03818_, _03392_);
  and (_03820_, _03431_, _26268_);
  nor (_03821_, _03820_, _26163_);
  nand (_03823_, _03458_, _23681_);
  and (_03824_, _03823_, _03821_);
  and (_03825_, _03824_, _03819_);
  and (_03826_, _03365_, _23205_);
  and (_03827_, _03374_, _25833_);
  or (_03828_, _03827_, _03826_);
  and (_03829_, _03828_, _03369_);
  nor (_03830_, _26365_, _23976_);
  and (_03831_, _26365_, _23413_);
  or (_03832_, _03831_, _03830_);
  and (_03834_, _03832_, _03378_);
  nor (_03835_, _26365_, _23357_);
  and (_03836_, _26365_, _23744_);
  or (_03837_, _03836_, _03835_);
  and (_03838_, _03837_, _03371_);
  or (_03839_, _03838_, _03834_);
  and (_03840_, _03365_, _24788_);
  and (_03841_, _03374_, _23247_);
  or (_03842_, _03841_, _03840_);
  and (_03843_, _03842_, _26365_);
  or (_03844_, _03843_, _03839_);
  nor (_03845_, _03844_, _03829_);
  nor (_03846_, _03845_, _03821_);
  or (_03847_, _03846_, _03825_);
  and (_27324_, _03847_, _22773_);
  and (_03848_, _26365_, _26076_);
  and (_03849_, _03848_, _03365_);
  nor (_03851_, _03196_, _26112_);
  and (_03852_, _03194_, _26013_);
  and (_03853_, _03852_, _03851_);
  and (_03854_, _03853_, _03849_);
  and (_03855_, _03854_, _26264_);
  and (_03856_, _26267_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_03857_, _03459_, _03394_);
  and (_03858_, _03848_, _03378_);
  and (_03859_, _03858_, _03857_);
  and (_03860_, _03859_, _03856_);
  nor (_03861_, _03194_, _26013_);
  and (_03862_, _03861_, _03849_);
  and (_03864_, _03862_, _03851_);
  and (_03865_, _03864_, _26284_);
  or (_03867_, _03865_, _03860_);
  nor (_03869_, _03867_, _03855_);
  nor (_03870_, _03869_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_03871_, _03870_);
  and (_03872_, _26374_, _22855_);
  and (_03873_, _03872_, _22910_);
  not (_03874_, _03873_);
  and (_03875_, _03854_, _26268_);
  and (_03877_, _03378_, _03369_);
  not (_03878_, _03877_);
  and (_03879_, _26160_, _24331_);
  and (_03880_, _03879_, _03878_);
  nor (_03881_, _03880_, _03875_);
  and (_03882_, _03881_, _03874_);
  nand (_03883_, _03882_, _03871_);
  and (_03884_, _03848_, _03374_);
  and (_03885_, _03884_, _03857_);
  and (_03886_, _03885_, _03856_);
  nor (_03887_, _03886_, rst);
  and (_27325_, _03887_, _03883_);
  and (_03888_, _26365_, _03393_);
  and (_03890_, _03888_, _03365_);
  and (_03891_, _03890_, _03395_);
  and (_03892_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_03893_, _26365_, _26076_);
  and (_03894_, _03893_, _03365_);
  and (_03895_, _03894_, _03395_);
  and (_03896_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_03897_, _03896_, _03892_);
  and (_03898_, _03893_, _03371_);
  and (_03900_, _03898_, _03395_);
  and (_03902_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_03903_, _03888_, _03374_);
  and (_03904_, _03903_, _03395_);
  and (_03905_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_03906_, _03905_, _03902_);
  or (_03907_, _03906_, _03897_);
  and (_03908_, _03890_, _03857_);
  and (_03909_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03911_, _03888_, _03378_);
  and (_03912_, _03911_, _03395_);
  and (_03913_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_03914_, _03913_, _03909_);
  and (_03916_, _03488_, _03394_);
  and (_03917_, _03890_, _03916_);
  and (_03918_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03919_, _03877_, _26076_);
  and (_03920_, _03488_, _03197_);
  and (_03921_, _03920_, _03919_);
  and (_03922_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03923_, _03922_, _03918_);
  or (_03924_, _03923_, _03914_);
  or (_03925_, _03924_, _03907_);
  and (_03926_, _03911_, _03857_);
  and (_03927_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_03928_, _03888_, _03371_);
  and (_03929_, _03928_, _03857_);
  and (_03930_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_03931_, _03930_, _03927_);
  and (_03933_, _03898_, _03857_);
  and (_03934_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_03935_, _03903_, _03857_);
  and (_03936_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_03938_, _03936_, _03934_);
  or (_03939_, _03938_, _03931_);
  and (_03940_, _03459_, _03197_);
  and (_03941_, _03940_, _03928_);
  and (_03942_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03943_, _03940_, _03890_);
  and (_03944_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03945_, _03944_, _03942_);
  and (_03946_, _03919_, _03857_);
  and (_03948_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_03949_, _03894_, _03857_);
  and (_03950_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_03951_, _03950_, _03948_);
  or (_03952_, _03951_, _03945_);
  or (_03953_, _03952_, _03939_);
  or (_03954_, _03953_, _03925_);
  and (_03955_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_03956_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03957_, _03956_, _03955_);
  and (_03958_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_03959_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_03960_, _03959_, _03958_);
  and (_03961_, _03849_, _03197_);
  and (_03962_, _03961_, _03430_);
  and (_03963_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03964_, _03848_, _03371_);
  and (_03967_, _03964_, _03857_);
  and (_03968_, _03967_, _26125_);
  or (_03970_, _03968_, _03963_);
  or (_03971_, _03970_, _03960_);
  and (_03973_, _03916_, _03849_);
  and (_03974_, _03973_, _03685_);
  and (_03975_, _03920_, _03849_);
  and (_03976_, _03975_, _03634_);
  or (_03977_, _03976_, _03974_);
  and (_03978_, _03849_, _03857_);
  and (_03979_, _03978_, _03785_);
  and (_03980_, _03940_, _03849_);
  and (_03982_, _03980_, _03738_);
  or (_03983_, _03982_, _03979_);
  or (_03985_, _03983_, _03977_);
  or (_03986_, _03985_, _03971_);
  or (_03987_, _03986_, _03957_);
  nor (_03988_, _03987_, _03954_);
  or (_03989_, _03988_, _03883_);
  not (_03990_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor (_03992_, _03895_, _03891_);
  nor (_03993_, _03904_, _03900_);
  and (_03994_, _03993_, _03992_);
  nor (_03996_, _03912_, _03908_);
  nor (_03997_, _03921_, _03917_);
  and (_03998_, _03997_, _03996_);
  and (_03999_, _03998_, _03994_);
  nor (_04000_, _03929_, _03926_);
  nor (_04001_, _03935_, _03933_);
  and (_04002_, _04001_, _04000_);
  nor (_04004_, _03943_, _03941_);
  nor (_04006_, _03949_, _03946_);
  and (_04007_, _04006_, _04004_);
  and (_04008_, _04007_, _04002_);
  and (_04010_, _04008_, _03999_);
  nor (_04012_, _03864_, _03854_);
  nor (_04014_, _03885_, _03859_);
  nor (_04015_, _03967_, _03962_);
  and (_04016_, _04015_, _04014_);
  nor (_04017_, _03975_, _03973_);
  nor (_04018_, _03980_, _03978_);
  and (_04019_, _04018_, _04017_);
  and (_04020_, _04019_, _04016_);
  and (_04021_, _04020_, _04012_);
  and (_04022_, _04021_, _04010_);
  nor (_04023_, _04022_, _03870_);
  and (_04024_, _04023_, _03882_);
  or (_04025_, _04024_, _03990_);
  and (_04027_, _04025_, _03989_);
  nor (_04029_, _04027_, _03886_);
  and (_04030_, _03886_, _00619_);
  or (_04032_, _04030_, _04029_);
  and (_27326_[7], _04032_, _22773_);
  and (_04033_, _25175_, _24108_);
  and (_04035_, _04033_, _24027_);
  not (_04036_, _04033_);
  and (_04038_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or (_25498_, _04038_, _04035_);
  and (_04039_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and (_04040_, _24795_, _23920_);
  or (_27013_, _04040_, _04039_);
  and (_04041_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  and (_04042_, _02718_, _23751_);
  or (_25549_, _04042_, _04041_);
  and (_04044_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  and (_04045_, _02756_, _23900_);
  or (_25553_, _04045_, _04044_);
  and (_04046_, _24098_, _24027_);
  and (_04047_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or (_25555_, _04047_, _04046_);
  and (_04049_, _02403_, _23751_);
  and (_04050_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_25563_, _04050_, _04049_);
  and (_04051_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_04052_, _02752_, _23715_);
  or (_25588_, _04052_, _04051_);
  and (_04053_, _01709_, _23900_);
  and (_04054_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_25598_, _04054_, _04053_);
  and (_04056_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_04057_, _02752_, _23693_);
  or (_25602_, _04057_, _04056_);
  and (_04058_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and (_04059_, _02838_, _23900_);
  or (_25616_, _04059_, _04058_);
  and (_04060_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_04061_, _02848_, _24027_);
  or (_25629_, _04061_, _04060_);
  and (_04062_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_04063_, _02752_, _23920_);
  or (_27015_, _04063_, _04062_);
  and (_04064_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_04065_, _02752_, _23900_);
  or (_27014_, _04065_, _04064_);
  and (_04066_, _02853_, _23693_);
  and (_04067_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or (_27132_, _04067_, _04066_);
  and (_04069_, _02350_, _23920_);
  and (_04070_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_25669_, _04070_, _04069_);
  and (_04071_, _02403_, _23693_);
  and (_04072_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_25675_, _04072_, _04071_);
  and (_04073_, _24237_, _24061_);
  and (_04074_, _04073_, _24053_);
  not (_04075_, _04073_);
  and (_04076_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_25679_, _04076_, _04074_);
  and (_04077_, _24237_, _24108_);
  and (_04078_, _04077_, _23983_);
  not (_04080_, _04077_);
  and (_04081_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_25699_, _04081_, _04078_);
  and (_04082_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  and (_04083_, _02718_, _23693_);
  or (_25722_, _04083_, _04082_);
  and (_04085_, _02244_, _24053_);
  and (_04087_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or (_25724_, _04087_, _04085_);
  and (_04089_, _23925_, _23751_);
  and (_04090_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_27246_, _04090_, _04089_);
  and (_04091_, _24157_, _23909_);
  and (_04092_, _04091_, _23900_);
  not (_04093_, _04091_);
  and (_04094_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  or (_25760_, _04094_, _04092_);
  and (_04095_, _24123_, _23909_);
  and (_04096_, _04095_, _23920_);
  not (_04097_, _04095_);
  and (_04098_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_27098_, _04098_, _04096_);
  and (_04100_, _04091_, _23751_);
  and (_04102_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  or (_25770_, _04102_, _04100_);
  and (_04104_, _04091_, _23715_);
  and (_04105_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  or (_25772_, _04105_, _04104_);
  and (_04106_, _04073_, _23715_);
  and (_04107_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_25783_, _04107_, _04106_);
  and (_04109_, _04073_, _23693_);
  and (_04110_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_25788_, _04110_, _04109_);
  and (_04111_, _04073_, _23751_);
  and (_04113_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_25793_, _04113_, _04111_);
  and (_04114_, _04077_, _24053_);
  and (_04116_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_25819_, _04116_, _04114_);
  and (_04117_, _04077_, _23751_);
  and (_04118_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or (_25834_, _04118_, _04117_);
  and (_04120_, _23892_, _23751_);
  and (_04121_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or (_25839_, _04121_, _04120_);
  and (_04123_, _04077_, _23715_);
  and (_04124_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or (_27063_, _04124_, _04123_);
  and (_04125_, _04077_, _23920_);
  and (_04127_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_25927_, _04127_, _04125_);
  and (_04128_, _24053_, _23707_);
  and (_04130_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_25935_, _04130_, _04128_);
  and (_04133_, _24053_, _23892_);
  and (_04134_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or (_27222_, _04134_, _04133_);
  and (_04135_, _04077_, _23900_);
  and (_04136_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or (_25950_, _04136_, _04135_);
  and (_04137_, _24901_, _23693_);
  and (_04138_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_26000_, _04138_, _04137_);
  and (_04141_, _24237_, _23444_);
  and (_04142_, _04141_, _23920_);
  not (_04143_, _04141_);
  and (_04144_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_26011_, _04144_, _04142_);
  and (_04146_, _04091_, _24027_);
  and (_04147_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  or (_26015_, _04147_, _04146_);
  and (_04149_, _04091_, _23983_);
  and (_04150_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  or (_26020_, _04150_, _04149_);
  and (_04151_, _24027_, _23454_);
  and (_04152_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or (_26029_, _04152_, _04151_);
  and (_04154_, _24164_, _23920_);
  and (_04155_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_26085_, _04155_, _04154_);
  and (_04156_, _24164_, _23693_);
  and (_04158_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_26115_, _04158_, _04156_);
  and (_04159_, _24164_, _23715_);
  and (_04160_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_27099_, _04160_, _04159_);
  and (_04162_, _04091_, _23920_);
  and (_04163_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  or (_26141_, _04163_, _04162_);
  and (_04164_, _04141_, _24053_);
  and (_04165_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or (_27068_, _04165_, _04164_);
  and (_04166_, _23925_, _23900_);
  and (_04167_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_26159_, _04167_, _04166_);
  not (_04169_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_04170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_04171_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_04172_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_04173_, _04172_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_04174_, _04173_, _04171_);
  and (_04175_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01967_);
  or (_04176_, _04175_, _04174_);
  nor (_04177_, _04176_, _04170_);
  nand (_04178_, _04177_, _04169_);
  nor (_04179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_04180_, _04179_, _04177_);
  nand (_04182_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_04183_, _04182_, _04180_);
  and (_04185_, _04183_, _22773_);
  and (_26162_, _04185_, _04178_);
  nand (_04186_, _24632_, _23759_);
  or (_04187_, _23759_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_04188_, _04187_, _22773_);
  and (_26835_[1], _04188_, _04186_);
  not (_04189_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and (_04190_, _01979_, _04189_);
  and (_04191_, _02140_, _01983_);
  and (_04192_, _04191_, _04190_);
  and (_04194_, _04192_, _02137_);
  not (_04195_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or (_04196_, _02142_, _04195_);
  nor (_04197_, _04196_, _04194_);
  or (_04198_, _04197_, _01970_);
  and (_26181_, _04198_, _22773_);
  and (_26184_, _04180_, _22773_);
  and (_04200_, _24237_, _23930_);
  and (_04201_, _04200_, _23983_);
  not (_04202_, _04200_);
  and (_04203_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_26194_, _04203_, _04201_);
  and (_04204_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or (_04205_, _04204_, _01970_);
  nor (_04206_, _01971_, rst);
  and (_26203_, _04206_, _04205_);
  and (_04207_, \oc8051_top_1.oc8051_sfr1.wait_data , _22773_);
  and (_04208_, _04207_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_04209_, _25905_, _25892_);
  and (_04210_, _26228_, _24678_);
  or (_04211_, _04210_, _03594_);
  and (_04213_, _26228_, _24715_);
  and (_04214_, _26228_, _24543_);
  or (_04215_, _04214_, _04213_);
  or (_04216_, _04215_, _04211_);
  or (_04218_, _04216_, _04209_);
  and (_04219_, _04218_, _24566_);
  nor (_04220_, _24671_, _24503_);
  and (_04222_, _25924_, _04220_);
  or (_04223_, _04222_, _24691_);
  or (_04224_, _04223_, _03596_);
  or (_04225_, _04224_, _03606_);
  and (_04227_, _01885_, _24670_);
  and (_04228_, _25856_, _24697_);
  or (_04229_, _04228_, _25916_);
  or (_04230_, _04229_, _04227_);
  and (_04231_, _24721_, _24678_);
  and (_04232_, _25856_, _24699_);
  or (_04233_, _04232_, _25891_);
  or (_04234_, _04233_, _04231_);
  nand (_04235_, _25856_, _24712_);
  nand (_04236_, _26239_, _04235_);
  or (_04237_, _04236_, _04234_);
  or (_04238_, _04237_, _04230_);
  or (_04240_, _04238_, _04225_);
  or (_04242_, _04240_, _04219_);
  and (_04243_, _04242_, _01886_);
  or (_26838_[0], _04243_, _04208_);
  or (_04244_, _02307_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_04246_, _02307_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_04247_, _04246_, _04244_);
  nand (_04249_, _04247_, _22773_);
  nor (_26206_, _04249_, _01970_);
  not (_04250_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_04251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_04252_, _04173_, _03402_);
  or (_04253_, _04252_, _04175_);
  nor (_04254_, _04253_, _04251_);
  nand (_04255_, _04254_, _04250_);
  nor (_04256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_04258_, _04256_, _04254_);
  nand (_04259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_04260_, _04259_, _04258_);
  and (_04261_, _04260_, _22773_);
  and (_26218_, _04261_, _04255_);
  and (_26220_, _04258_, _22773_);
  and (_04262_, _23983_, _23454_);
  and (_04263_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or (_27211_, _04263_, _04262_);
  and (_04264_, _04141_, _23715_);
  and (_04265_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or (_26233_, _04265_, _04264_);
  not (_04266_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_04267_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _03476_);
  not (_04268_, _04267_);
  nor (_04269_, _01975_, _02207_);
  and (_04270_, _04269_, _04268_);
  and (_04271_, _04270_, _02219_);
  nor (_04272_, _04271_, _04266_);
  and (_04273_, _04271_, rxd_i);
  or (_04274_, _04273_, rst);
  or (_26235_, _04274_, _04272_);
  or (_04275_, _02199_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_04277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_04278_, _04277_, _01975_);
  or (_04280_, _04278_, _02179_);
  nand (_04281_, _04280_, _04275_);
  nand (_26237_, _04281_, _01751_);
  and (_04282_, _04141_, _23693_);
  and (_04283_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or (_26248_, _04283_, _04282_);
  and (_04284_, _04141_, _23751_);
  and (_04285_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or (_26251_, _04285_, _04284_);
  and (_04286_, _04200_, _23751_);
  and (_04287_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_26280_, _04287_, _04286_);
  and (_04288_, _04200_, _24053_);
  and (_04289_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_27064_, _04289_, _04288_);
  and (_04291_, _04073_, _23983_);
  and (_04292_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_26299_, _04292_, _04291_);
  and (_04293_, _04200_, _23715_);
  and (_04295_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_26316_, _04295_, _04293_);
  and (_04296_, _04200_, _23920_);
  and (_04298_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_27067_, _04298_, _04296_);
  and (_04300_, _04200_, _23900_);
  and (_04301_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_27066_, _04301_, _04300_);
  nor (_27323_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_04303_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_04304_, _03185_, rst);
  and (_27323_[1], _04304_, _04303_);
  nor (_04305_, _03185_, _03184_);
  or (_04306_, _04305_, _03186_);
  and (_04308_, _03190_, _22773_);
  and (_27323_[2], _04308_, _04306_);
  nand (_04310_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_04311_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_04312_, _04311_, _04310_);
  nand (_04313_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_04315_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_04316_, _04315_, _04313_);
  and (_04317_, _04316_, _04312_);
  nand (_04318_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_04319_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_04320_, _04319_, _04318_);
  nand (_04321_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_04322_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_04323_, _04322_, _04321_);
  and (_04324_, _04323_, _04320_);
  and (_04325_, _04324_, _04317_);
  nand (_04326_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_04327_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_04328_, _04327_, _04326_);
  nand (_04329_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_04330_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_04332_, _04330_, _04329_);
  and (_04333_, _04332_, _04328_);
  nand (_04334_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_04335_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_04336_, _04335_, _04334_);
  nand (_04337_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_04338_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_04339_, _04338_, _04337_);
  and (_04340_, _04339_, _04336_);
  and (_04341_, _04340_, _04333_);
  and (_04342_, _04341_, _04325_);
  nand (_04343_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand (_04344_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_04345_, _04344_, _04343_);
  nand (_04346_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_04347_, _03967_, _26325_);
  and (_04348_, _04347_, _04346_);
  and (_04349_, _04348_, _04345_);
  nand (_04350_, _03973_, _03673_);
  nand (_04351_, _03975_, _03622_);
  and (_04352_, _04351_, _04350_);
  nand (_04353_, _03980_, _03727_);
  nand (_04354_, _03978_, _03775_);
  and (_04355_, _04354_, _04353_);
  and (_04356_, _04355_, _04352_);
  and (_04358_, _04356_, _04349_);
  not (_04359_, _03864_);
  or (_04360_, _04359_, _03363_);
  nand (_04361_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_04362_, _04361_, _04360_);
  and (_04363_, _04362_, _04358_);
  and (_04364_, _04363_, _04342_);
  nor (_04365_, _04364_, _03883_);
  not (_04366_, _03886_);
  not (_04367_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_04368_, _04024_, _04367_);
  nand (_04369_, _04368_, _04366_);
  or (_04370_, _04369_, _04365_);
  or (_04371_, _04366_, _26798_);
  and (_04372_, _04371_, _22773_);
  and (_27326_[0], _04372_, _04370_);
  not (_04373_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_04374_, _04024_, _04373_);
  nand (_04375_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_04376_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_04377_, _04376_, _04375_);
  nand (_04378_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_04379_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_04380_, _04379_, _04378_);
  and (_04381_, _04380_, _04377_);
  nand (_04382_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_04383_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_04384_, _04383_, _04382_);
  nand (_04385_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nand (_04386_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04387_, _04386_, _04385_);
  and (_04388_, _04387_, _04384_);
  and (_04389_, _04388_, _04381_);
  nand (_04390_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_04391_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_04392_, _04391_, _04390_);
  nand (_04393_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_04394_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_04395_, _04394_, _04393_);
  and (_04396_, _04395_, _04392_);
  nand (_04397_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  nand (_04398_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_04399_, _04398_, _04397_);
  nand (_04400_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_04401_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_04402_, _04401_, _04400_);
  and (_04403_, _04402_, _04399_);
  and (_04404_, _04403_, _04396_);
  and (_04405_, _04404_, _04389_);
  nand (_04406_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand (_04407_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_04408_, _04407_, _04406_);
  nand (_04409_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand (_04410_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_04411_, _04410_, _04409_);
  nand (_04412_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_04413_, _03967_, _26303_);
  and (_04414_, _04413_, _04412_);
  and (_04415_, _04414_, _04411_);
  nand (_04416_, _03973_, _03700_);
  nand (_04417_, _03975_, _03647_);
  and (_04418_, _04417_, _04416_);
  nand (_04419_, _03978_, _03796_);
  nand (_04420_, _03980_, _03751_);
  and (_04421_, _04420_, _04419_);
  and (_04422_, _04421_, _04418_);
  and (_04423_, _04422_, _04415_);
  and (_04424_, _04423_, _04408_);
  and (_04425_, _04424_, _04405_);
  or (_04426_, _04425_, _03883_);
  and (_04427_, _04426_, _04374_);
  nand (_04428_, _04427_, _04366_);
  or (_04429_, _04366_, _00101_);
  and (_04430_, _04429_, _22773_);
  and (_27326_[1], _04430_, _04428_);
  and (_04431_, _03886_, _00183_);
  not (_04432_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or (_04433_, _04024_, _04432_);
  and (_04434_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_04435_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_04436_, _04435_, _04434_);
  and (_04437_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_04438_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_04439_, _04438_, _04437_);
  or (_04440_, _04439_, _04436_);
  and (_04441_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_04442_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_04443_, _04442_, _04441_);
  and (_04444_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_04445_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_04446_, _04445_, _04444_);
  or (_04447_, _04446_, _04443_);
  or (_04448_, _04447_, _04440_);
  and (_04449_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_04450_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_04451_, _04450_, _04449_);
  and (_04452_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_04453_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_04454_, _04453_, _04452_);
  or (_04455_, _04454_, _04451_);
  and (_04456_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04457_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_04458_, _04457_, _04456_);
  and (_04459_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_04460_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_04461_, _04460_, _04459_);
  or (_04462_, _04461_, _04458_);
  or (_04463_, _04462_, _04455_);
  or (_04464_, _04463_, _04448_);
  and (_04465_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_04466_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_04467_, _04466_, _04465_);
  and (_04468_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_04469_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_04470_, _04469_, _04468_);
  and (_04471_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_04472_, _03967_, _26359_);
  or (_04473_, _04472_, _04471_);
  or (_04474_, _04473_, _04470_);
  and (_04475_, _03973_, _03706_);
  and (_04476_, _03975_, _03653_);
  or (_04477_, _04476_, _04475_);
  and (_04478_, _03978_, _03803_);
  and (_04479_, _03980_, _03757_);
  or (_04480_, _04479_, _04478_);
  or (_04481_, _04480_, _04477_);
  or (_04482_, _04481_, _04474_);
  or (_04483_, _04482_, _04467_);
  nor (_04484_, _04483_, _04464_);
  or (_04485_, _04484_, _03883_);
  and (_04486_, _04485_, _04433_);
  nor (_04487_, _04486_, _03886_);
  or (_04488_, _04487_, _04431_);
  and (_27326_[2], _04488_, _22773_);
  not (_04489_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_04490_, _04024_, _04489_);
  nand (_04491_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand (_04492_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_04493_, _04492_, _04491_);
  nand (_04494_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand (_04495_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_04496_, _04495_, _04494_);
  and (_04497_, _04496_, _04493_);
  nand (_04498_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nand (_04499_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_04500_, _04499_, _04498_);
  nand (_04501_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand (_04502_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_04503_, _04502_, _04501_);
  and (_04504_, _04503_, _04500_);
  and (_04505_, _04504_, _04497_);
  nand (_04506_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_04507_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_04508_, _04507_, _04506_);
  nand (_04509_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_04510_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_04511_, _04510_, _04509_);
  and (_04512_, _04511_, _04508_);
  nand (_04513_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand (_04514_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_04515_, _04514_, _04513_);
  nand (_04516_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  nand (_04517_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_04518_, _04517_, _04516_);
  and (_04519_, _04518_, _04515_);
  and (_04520_, _04519_, _04512_);
  and (_04521_, _04520_, _04505_);
  nand (_04523_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_04524_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_04525_, _04524_, _04523_);
  nand (_04526_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand (_04527_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_04528_, _04527_, _04526_);
  nand (_04529_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_04530_, _03967_, _26054_);
  and (_04532_, _04530_, _04529_);
  and (_04533_, _04532_, _04528_);
  nand (_04534_, _03973_, _03681_);
  nand (_04535_, _03975_, _03629_);
  and (_04536_, _04535_, _04534_);
  nand (_04537_, _03978_, _03781_);
  nand (_04538_, _03980_, _03734_);
  and (_04539_, _04538_, _04537_);
  and (_04541_, _04539_, _04536_);
  and (_04542_, _04541_, _04533_);
  and (_04543_, _04542_, _04525_);
  and (_04544_, _04543_, _04521_);
  or (_04545_, _04544_, _03883_);
  and (_04546_, _04545_, _04490_);
  nand (_04547_, _04546_, _04366_);
  or (_04548_, _04366_, _00277_);
  and (_04549_, _04548_, _22773_);
  and (_27326_[3], _04549_, _04547_);
  not (_04550_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_04551_, _04024_, _04550_);
  nand (_04553_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand (_04554_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_04555_, _04554_, _04553_);
  nand (_04556_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand (_04557_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_04558_, _04557_, _04556_);
  and (_04560_, _04558_, _04555_);
  nand (_04561_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand (_04563_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_04564_, _04563_, _04561_);
  nand (_04565_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_04566_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_04568_, _04566_, _04565_);
  and (_04569_, _04568_, _04564_);
  and (_04570_, _04569_, _04560_);
  nand (_04571_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_04572_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_04573_, _04572_, _04571_);
  nand (_04574_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_04576_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_04577_, _04576_, _04574_);
  and (_04578_, _04577_, _04573_);
  nand (_04579_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand (_04581_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_04582_, _04581_, _04579_);
  nand (_04583_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  nand (_04585_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_04586_, _04585_, _04583_);
  and (_04587_, _04586_, _04582_);
  and (_04588_, _04587_, _04578_);
  and (_04589_, _04588_, _04570_);
  nand (_04590_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand (_04591_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_04592_, _04591_, _04590_);
  nand (_04593_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_04594_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_04595_, _04594_, _04593_);
  nand (_04596_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_04598_, _25982_);
  nand (_04599_, _03967_, _04598_);
  and (_04600_, _04599_, _04596_);
  and (_04601_, _04600_, _04595_);
  nand (_04602_, _03973_, _03668_);
  nand (_04604_, _03975_, _03617_);
  and (_04605_, _04604_, _04602_);
  nand (_04606_, _03980_, _03721_);
  nand (_04607_, _03978_, _03770_);
  and (_04608_, _04607_, _04606_);
  and (_04609_, _04608_, _04605_);
  and (_04610_, _04609_, _04601_);
  and (_04611_, _04610_, _04592_);
  and (_04612_, _04611_, _04589_);
  or (_04614_, _04612_, _03883_);
  and (_04615_, _04614_, _04551_);
  nand (_04616_, _04615_, _04366_);
  or (_04617_, _04366_, _00352_);
  and (_04618_, _04617_, _22773_);
  and (_27326_[4], _04618_, _04616_);
  not (_04619_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor (_04621_, _04024_, _04619_);
  nand (_04622_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand (_04623_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04624_, _04623_, _04622_);
  nand (_04625_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  nand (_04627_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04628_, _04627_, _04625_);
  and (_04629_, _04628_, _04624_);
  nand (_04630_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand (_04631_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04632_, _04631_, _04630_);
  nand (_04634_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand (_04635_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_04636_, _04635_, _04634_);
  and (_04637_, _04636_, _04632_);
  and (_04639_, _04637_, _04629_);
  nand (_04640_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand (_04641_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_04642_, _04641_, _04640_);
  nand (_04643_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand (_04644_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_04645_, _04644_, _04643_);
  and (_04646_, _04645_, _04642_);
  nand (_04647_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nand (_04648_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_04649_, _04648_, _04647_);
  nand (_04650_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  nand (_04651_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_04652_, _04651_, _04650_);
  and (_04653_, _04652_, _04649_);
  and (_04654_, _04653_, _04646_);
  and (_04655_, _04654_, _04639_);
  nand (_04656_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_04657_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_04658_, _04657_, _04656_);
  and (_04660_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_04661_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_04662_, _04661_, _04660_);
  nand (_04663_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_04665_, _26035_);
  nand (_04666_, _03967_, _04665_);
  and (_04667_, _04666_, _04663_);
  and (_04668_, _04667_, _04662_);
  nand (_04669_, _03973_, _03695_);
  nand (_04670_, _03975_, _03642_);
  and (_04671_, _04670_, _04669_);
  nand (_04672_, _03980_, _03746_);
  nand (_04673_, _03978_, _03792_);
  and (_04674_, _04673_, _04672_);
  and (_04676_, _04674_, _04671_);
  and (_04677_, _04676_, _04668_);
  and (_04678_, _04677_, _04658_);
  and (_04680_, _04678_, _04655_);
  nor (_04681_, _04680_, _03883_);
  or (_04682_, _04681_, _03886_);
  or (_04683_, _04682_, _04621_);
  or (_04684_, _04366_, _00443_);
  and (_04686_, _04684_, _22773_);
  and (_27326_[5], _04686_, _04683_);
  and (_04688_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_04689_, _03895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_04691_, _04689_, _04688_);
  and (_04692_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_04694_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_04695_, _04694_, _04692_);
  or (_04697_, _04695_, _04691_);
  and (_04698_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_04699_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_04700_, _04699_, _04698_);
  and (_04702_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_04704_, _03917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_04705_, _04704_, _04702_);
  or (_04707_, _04705_, _04700_);
  or (_04708_, _04707_, _04697_);
  and (_04709_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_04710_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or (_04711_, _04710_, _04709_);
  and (_04712_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_04714_, _03935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_04715_, _04714_, _04712_);
  or (_04717_, _04715_, _04711_);
  and (_04718_, _03943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_04719_, _03941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_04721_, _04719_, _04718_);
  and (_04722_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_04724_, _03946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_04725_, _04724_, _04722_);
  or (_04727_, _04725_, _04721_);
  or (_04728_, _04727_, _04717_);
  or (_04730_, _04728_, _04708_);
  and (_04731_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_04733_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_04734_, _04733_, _04731_);
  and (_04735_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_04736_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_04738_, _04736_, _04735_);
  and (_04740_, _03962_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_04741_, _26091_);
  and (_04742_, _03967_, _04741_);
  or (_04744_, _04742_, _04740_);
  or (_04745_, _04744_, _04738_);
  and (_04746_, _03973_, _03710_);
  and (_04747_, _03975_, _03657_);
  or (_04748_, _04747_, _04746_);
  and (_04749_, _03980_, _03761_);
  and (_04750_, _03978_, _03807_);
  or (_04751_, _04750_, _04749_);
  or (_04752_, _04751_, _04748_);
  or (_04753_, _04752_, _04745_);
  or (_04754_, _04753_, _04734_);
  or (_04755_, _04754_, _04730_);
  and (_04756_, _04755_, _03871_);
  not (_04757_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor (_04758_, _04023_, _04757_);
  nor (_04759_, _04758_, _04756_);
  nand (_04760_, _04759_, _03882_);
  or (_04761_, _03882_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_04762_, _04761_, _04760_);
  or (_04763_, _04762_, _03886_);
  or (_04765_, _04366_, _00564_);
  and (_04766_, _04765_, _22773_);
  and (_27326_[6], _04766_, _04763_);
  and (_04767_, _24123_, _23706_);
  and (_04768_, _04767_, _23693_);
  not (_04769_, _04767_);
  and (_04770_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_00033_, _04770_, _04768_);
  and (_04771_, _23987_, _23700_);
  and (_04772_, _04771_, _23920_);
  not (_04773_, _04771_);
  and (_04774_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or (_00105_, _04774_, _04772_);
  and (_04775_, _25428_, _23715_);
  and (_04777_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_00125_, _04777_, _04775_);
  and (_04778_, _01927_, _24027_);
  and (_04779_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_00142_, _04779_, _04778_);
  and (_04782_, _04771_, _24027_);
  and (_04783_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or (_00164_, _04783_, _04782_);
  and (_04786_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_04787_, _02848_, _23920_);
  or (_00375_, _04787_, _04786_);
  and (_04788_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_04790_, _02848_, _23715_);
  or (_00379_, _04790_, _04788_);
  and (_04792_, _24543_, _24669_);
  and (_04793_, _24721_, _04792_);
  nor (_04794_, _04793_, _25850_);
  nor (_04795_, _04794_, _26810_);
  and (_04796_, _24721_, _24712_);
  nor (_04797_, _04796_, _25901_);
  not (_04799_, _25897_);
  and (_04800_, _24722_, _24639_);
  not (_04801_, _04800_);
  and (_04802_, _24721_, _24674_);
  nor (_04803_, _04802_, _25879_);
  and (_04805_, _04803_, _04801_);
  and (_04806_, _04805_, _04799_);
  not (_04807_, _25920_);
  and (_04808_, _04794_, _04807_);
  nor (_04809_, _24676_, _24669_);
  and (_04811_, _24542_, _04809_);
  and (_04812_, _24721_, _04811_);
  not (_04813_, _04812_);
  and (_04814_, _04813_, _25878_);
  and (_04815_, _04814_, _04808_);
  and (_04816_, _04815_, _04806_);
  and (_04817_, _04816_, _04797_);
  nor (_04818_, _04817_, _24647_);
  nor (_04819_, _04818_, _04795_);
  not (_04820_, _04819_);
  or (_04821_, _04820_, _26345_);
  or (_04822_, _04819_, _26153_);
  or (_04823_, _04822_, _26076_);
  nand (_04824_, _04823_, _04821_);
  and (_04825_, _04824_, _23422_);
  nor (_04826_, _04824_, _23422_);
  nor (_04827_, _04826_, _04825_);
  or (_04828_, _04820_, _26312_);
  or (_04830_, _04822_, _26013_);
  and (_04832_, _04830_, _04828_);
  and (_04833_, _04832_, _23429_);
  nor (_04834_, _04832_, _23429_);
  or (_04835_, _04834_, _04833_);
  and (_04836_, _04835_, _04827_);
  not (_04837_, _23445_);
  nor (_04838_, _02548_, _26153_);
  nor (_04839_, _04838_, _03194_);
  and (_04840_, _04839_, _04837_);
  not (_04841_, _04840_);
  not (_04842_, _23703_);
  nor (_04843_, _04838_, _26112_);
  nor (_04844_, _04843_, _04842_);
  and (_04845_, _04843_, _04842_);
  nor (_04846_, _04845_, _04844_);
  and (_04847_, _04846_, _04841_);
  not (_04848_, _26156_);
  nor (_04849_, _04838_, _26013_);
  nor (_04850_, _04849_, _23448_);
  nor (_04851_, _04839_, _04837_);
  nor (_04852_, _04851_, _04850_);
  and (_04853_, _04852_, _04848_);
  and (_04854_, _04853_, _04847_);
  and (_04856_, _04854_, _04836_);
  nor (_04857_, _04838_, _03393_);
  and (_04858_, _04838_, _26112_);
  nor (_04859_, _04858_, _04857_);
  and (_04860_, _04859_, _23436_);
  nor (_04861_, _04859_, _23436_);
  or (_04863_, _04861_, _04860_);
  not (_04864_, _04863_);
  not (_04865_, _23442_);
  nor (_04866_, _04820_, _26365_);
  nor (_04867_, _04822_, _26041_);
  nor (_04868_, _04867_, _04866_);
  nor (_04869_, _04868_, _04865_);
  and (_04870_, _04868_, _04865_);
  nor (_04871_, _04870_, _04869_);
  and (_04872_, _04871_, _04864_);
  and (_04873_, _04849_, _23448_);
  nor (_04874_, _04873_, _23424_);
  and (_04875_, _04874_, _04872_);
  and (_04876_, _04875_, _04856_);
  and (_26881_, _04876_, _22773_);
  nor (_26882_[7], _23982_, rst);
  nor (_26884_[2], _26365_, rst);
  and (_04877_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  and (_04879_, _02842_, _24027_);
  or (_00418_, _04879_, _04877_);
  and (_04880_, _01932_, _23693_);
  and (_04881_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_00421_, _04881_, _04880_);
  and (_04883_, _02853_, _23983_);
  and (_04884_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or (_27135_, _04884_, _04883_);
  and (_04886_, _04073_, _24027_);
  and (_04887_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_00437_, _04887_, _04886_);
  and (_04888_, _04073_, _23920_);
  and (_04889_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_00445_, _04889_, _04888_);
  and (_04890_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_04891_, _02848_, _23983_);
  or (_00490_, _04891_, _04890_);
  and (_04892_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and (_04893_, _02662_, _24027_);
  or (_00510_, _04893_, _04892_);
  and (_04895_, _02455_, _23983_);
  and (_04896_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or (_00516_, _04896_, _04895_);
  and (_04899_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  and (_04900_, _02842_, _23693_);
  or (_00520_, _04900_, _04899_);
  and (_04901_, _24237_, _24123_);
  and (_04902_, _04901_, _24027_);
  not (_04904_, _04901_);
  and (_04905_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or (_00525_, _04905_, _04902_);
  and (_04906_, _04901_, _23920_);
  and (_04908_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_00537_, _04908_, _04906_);
  and (_26882_[0], _24052_, _22773_);
  and (_26882_[1], _23750_, _22773_);
  and (_26882_[2], _23692_, _22773_);
  and (_26882_[3], _23714_, _22773_);
  and (_26882_[4], _23899_, _22773_);
  and (_26882_[5], _23919_, _22773_);
  nor (_26882_[6], _24026_, rst);
  nor (_26884_[0], _26345_, rst);
  nor (_26884_[1], _26312_, rst);
  and (_04911_, _02326_, _24027_);
  and (_04912_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or (_00629_, _04912_, _04911_);
  and (_04913_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  and (_04914_, _02842_, _23983_);
  or (_27139_, _04914_, _04913_);
  and (_04915_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_04916_, _04915_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_04917_, _04915_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_04918_, _04917_, _04916_);
  and (_00732_, _04918_, _22773_);
  and (_04919_, _24696_, _24669_);
  and (_04920_, _04919_, _25856_);
  and (_04921_, _24699_, _24615_);
  or (_04922_, _04921_, _04920_);
  and (_04923_, _25856_, _24682_);
  and (_04924_, _24697_, _24615_);
  or (_04925_, _04924_, _04923_);
  or (_04926_, _04925_, _04922_);
  or (_04927_, _04213_, _04210_);
  or (_04928_, _04228_, _04214_);
  or (_04929_, _04928_, _04927_);
  or (_04931_, _04929_, _04926_);
  and (_04932_, _25930_, _25856_);
  and (_04934_, _25856_, _25849_);
  and (_04935_, _25856_, _24722_);
  or (_04937_, _04935_, _04934_);
  or (_04938_, _04937_, _04932_);
  or (_04939_, _04938_, _04234_);
  or (_04940_, _04939_, _04931_);
  and (_04941_, _26231_, _24698_);
  and (_04942_, _24543_, _24615_);
  or (_04943_, _04942_, _04941_);
  and (_04944_, _24543_, _24690_);
  and (_04945_, _26231_, _24677_);
  or (_04947_, _04945_, _04944_);
  or (_04948_, _04947_, _04943_);
  and (_04949_, _24542_, _24648_);
  or (_04950_, _04949_, _24702_);
  or (_04952_, _04950_, _04948_);
  or (_04953_, _03597_, _25926_);
  or (_04954_, _03596_, _03594_);
  or (_04955_, _04954_, _04953_);
  or (_04957_, _24716_, _24693_);
  or (_04959_, _04957_, _24675_);
  or (_04960_, _04959_, _04955_);
  or (_04961_, _04960_, _04952_);
  or (_04962_, _04961_, _04940_);
  and (_04963_, _04962_, _23760_);
  and (_04964_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_04965_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_04966_, _25848_, _04965_);
  not (_04967_, _24697_);
  not (_04968_, _24616_);
  or (_04969_, _25886_, _04968_);
  nor (_04970_, _04969_, _04967_);
  nor (_04971_, _04970_, _01885_);
  not (_04973_, _04971_);
  and (_04975_, _04973_, _04966_);
  or (_04977_, _04975_, _04964_);
  or (_04979_, _04977_, _04963_);
  and (_26837_[0], _04979_, _22773_);
  not (_04981_, word_in[7]);
  nor (_04982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04983_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01548_);
  nor (_04985_, _04983_, _04982_);
  not (_04986_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_04988_, _00319_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04989_, _01548_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_04991_, _04989_, _04988_);
  and (_04992_, _04991_, _04986_);
  nor (_04993_, _04991_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_04994_, _04993_, _04992_);
  not (_04995_, _04994_);
  nor (_04996_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04998_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01548_);
  nor (_04999_, _04998_, _04996_);
  not (_05001_, _04999_);
  nor (_05002_, _00224_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_05003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01548_);
  nor (_05005_, _05003_, _05002_);
  and (_05006_, _05005_, _05001_);
  nand (_05007_, _05006_, _04995_);
  and (_05008_, _05007_, _04985_);
  nor (_05009_, _05005_, _05001_);
  not (_05010_, _05009_);
  not (_05011_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_05012_, _04991_, _05011_);
  and (_05013_, _04991_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05014_, _05013_, _05012_);
  nor (_05015_, _05014_, _05010_);
  and (_05016_, _05005_, _04999_);
  not (_05017_, _05016_);
  not (_05018_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_05019_, _04991_, _05018_);
  and (_05020_, _04991_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_05021_, _05020_, _05019_);
  nor (_05022_, _05021_, _05017_);
  nor (_05023_, _05022_, _05015_);
  not (_05024_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05025_, _04991_, _05024_);
  nor (_05026_, _04991_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_05027_, _05005_, _04999_);
  not (_05028_, _05027_);
  or (_05029_, _05028_, _05026_);
  or (_05030_, _05029_, _05025_);
  and (_05031_, _05030_, _05023_);
  and (_05032_, _05031_, _05008_);
  not (_05033_, _04985_);
  not (_05035_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_05036_, _04991_, _05035_);
  and (_05037_, _04991_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05038_, _05037_, _05036_);
  nor (_05039_, _05038_, _05005_);
  not (_05040_, _05005_);
  not (_05041_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05042_, _04991_, _05041_);
  nor (_05043_, _04991_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_05044_, _05043_, _05042_);
  nor (_05045_, _05044_, _05040_);
  nor (_05046_, _05045_, _05039_);
  nor (_05047_, _05046_, _04999_);
  nor (_05048_, _04991_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_05049_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05050_, _04991_, _05049_);
  or (_05051_, _05050_, _05048_);
  nor (_05052_, _05051_, _05017_);
  and (_05053_, _04991_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_05054_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05055_, _04991_, _05054_);
  nor (_05056_, _05055_, _05053_);
  nor (_05057_, _05056_, _05010_);
  nor (_05058_, _05057_, _05052_);
  not (_05059_, _05058_);
  nor (_05061_, _05059_, _05047_);
  and (_05062_, _05061_, _05033_);
  nor (_05063_, _05062_, _05032_);
  nor (_05064_, _05063_, _04981_);
  not (_05065_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_05067_, _04985_, _05065_);
  or (_05068_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_05069_, _05068_, _05067_);
  and (_05070_, _05069_, _05027_);
  or (_05071_, _05070_, _04991_);
  not (_05072_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_05073_, _04985_, _05072_);
  or (_05074_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_05075_, _05074_, _05073_);
  and (_05076_, _05075_, _05016_);
  not (_05077_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_05079_, _04985_, _05077_);
  or (_05080_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_05081_, _05080_, _05079_);
  and (_05082_, _05081_, _05006_);
  not (_05083_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_05084_, _04985_, _05083_);
  or (_05085_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_05086_, _05085_, _05084_);
  and (_05087_, _05086_, _05009_);
  or (_05088_, _05087_, _05082_);
  or (_05089_, _05088_, _05076_);
  or (_05090_, _05089_, _05071_);
  not (_05091_, _04991_);
  not (_05092_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_05093_, _04985_, _05092_);
  or (_05094_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05096_, _05094_, _05093_);
  and (_05097_, _05096_, _05027_);
  or (_05098_, _05097_, _05091_);
  not (_05099_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_05100_, _04985_, _05099_);
  or (_05101_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_05102_, _05101_, _05100_);
  and (_05103_, _05102_, _05006_);
  not (_05104_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_05105_, _04985_, _05104_);
  or (_05107_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_05108_, _05107_, _05105_);
  and (_05109_, _05108_, _05016_);
  or (_05110_, _05109_, _05103_);
  not (_05111_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_05112_, _04985_, _05111_);
  or (_05113_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_05114_, _05113_, _05112_);
  and (_05115_, _05114_, _05009_);
  or (_05116_, _05115_, _05110_);
  or (_05117_, _05116_, _05098_);
  and (_05118_, _05117_, _05090_);
  and (_05119_, _05118_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _05119_, _05064_);
  nor (_05120_, _04999_, _04985_);
  not (_05122_, _05120_);
  and (_05123_, _04999_, _04985_);
  and (_05124_, _05123_, _05005_);
  nor (_05125_, _05123_, _05005_);
  nor (_05126_, _05125_, _05124_);
  not (_05127_, _05126_);
  nor (_05128_, _05127_, _04994_);
  nor (_05129_, _05124_, _05091_);
  nor (_05130_, _05040_, _04991_);
  and (_05131_, _05130_, _05123_);
  nor (_05132_, _05131_, _05129_);
  nor (_05133_, _05132_, _05126_);
  and (_05134_, _05133_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05135_, _05132_, _05127_);
  and (_05136_, _05135_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05137_, _05136_, _05134_);
  nor (_05138_, _05137_, _05128_);
  nor (_05139_, _05138_, _05122_);
  not (_05140_, _05139_);
  and (_05141_, _05124_, _04991_);
  nand (_05142_, _05141_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_05143_, _05123_);
  nor (_05144_, _05127_, _05044_);
  and (_05145_, _05133_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05146_, _05145_, _05144_);
  or (_05148_, _05146_, _05143_);
  and (_05149_, _05148_, _05142_);
  and (_05150_, _05149_, _05140_);
  and (_05151_, _05001_, _04985_);
  not (_05153_, _05151_);
  nor (_05154_, _05127_, _05051_);
  and (_05155_, _05135_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_05156_, _05133_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05157_, _05156_, _05155_);
  nor (_05159_, _05157_, _05154_);
  nor (_05160_, _05159_, _05153_);
  and (_05161_, _04999_, _05033_);
  not (_05162_, _05161_);
  nor (_05163_, _05127_, _05021_);
  and (_05164_, _05135_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05165_, _05133_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05166_, _05165_, _05164_);
  nor (_05167_, _05166_, _05163_);
  nor (_05168_, _05167_, _05162_);
  nor (_05169_, _05168_, _05160_);
  and (_05170_, _05169_, _05150_);
  or (_05172_, _05120_, _05123_);
  not (_05173_, _05172_);
  not (_05174_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_05176_, _04985_, _05174_);
  or (_05177_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_05178_, _05177_, _05176_);
  and (_05179_, _05178_, _05173_);
  not (_05180_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_05181_, _04985_, _05180_);
  or (_05182_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_05183_, _05182_, _05181_);
  and (_05184_, _05183_, _05172_);
  or (_05185_, _05184_, _05179_);
  and (_05186_, _05185_, _05135_);
  not (_05187_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_05188_, _04985_, _05187_);
  or (_05189_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_05190_, _05189_, _05188_);
  and (_05191_, _05190_, _05173_);
  not (_05193_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_05194_, _04985_, _05193_);
  or (_05196_, _04985_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_05197_, _05196_, _05194_);
  and (_05198_, _05197_, _05172_);
  or (_05199_, _05198_, _05191_);
  and (_05201_, _05199_, _05133_);
  and (_05202_, _05126_, _05091_);
  not (_05204_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_05205_, _04985_, _05204_);
  or (_05206_, _04985_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_05207_, _05206_, _05205_);
  and (_05208_, _05207_, _05173_);
  not (_05209_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_05210_, _04985_, _05209_);
  or (_05212_, _04985_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_05213_, _05212_, _05210_);
  and (_05214_, _05213_, _05172_);
  or (_05215_, _05214_, _05208_);
  and (_05217_, _05215_, _05202_);
  and (_05218_, _05126_, _04991_);
  not (_05219_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_05220_, _04985_, _05219_);
  or (_05221_, _04985_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_05222_, _05221_, _05220_);
  and (_05223_, _05222_, _05173_);
  not (_05224_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_05225_, _04985_, _05224_);
  or (_05226_, _04985_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_05227_, _05226_, _05225_);
  and (_05228_, _05227_, _05172_);
  or (_05229_, _05228_, _05223_);
  and (_05230_, _05229_, _05218_);
  or (_05232_, _05230_, _05217_);
  or (_05233_, _05232_, _05201_);
  nor (_05234_, _05233_, _05186_);
  nor (_05235_, _05234_, _05170_);
  and (_05236_, _05170_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _05236_, _05235_);
  nor (_05238_, _05027_, _05016_);
  nor (_05239_, _05016_, _04991_);
  and (_05240_, _05016_, _04991_);
  nor (_05241_, _05240_, _05239_);
  nor (_05242_, _05241_, _05238_);
  and (_05243_, _05242_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_05245_, _05238_);
  and (_05246_, _05241_, _05245_);
  and (_05247_, _05246_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05248_, _05245_, _05051_);
  or (_05249_, _05248_, _05247_);
  nor (_05250_, _05249_, _05243_);
  nor (_05251_, _05250_, _05122_);
  not (_05252_, _05251_);
  nor (_05253_, _05245_, _05044_);
  and (_05254_, _05242_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05255_, _05246_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05257_, _05255_, _05254_);
  or (_05258_, _05257_, _05253_);
  nand (_05260_, _05258_, _05161_);
  and (_05261_, _05260_, _05252_);
  nor (_05262_, _05245_, _04994_);
  and (_05263_, _05246_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05264_, _05242_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05265_, _05264_, _05263_);
  nor (_05266_, _05265_, _05262_);
  nor (_05267_, _05266_, _05143_);
  nor (_05269_, _05245_, _05021_);
  and (_05270_, _05246_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05271_, _05242_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05273_, _05271_, _05270_);
  nor (_05274_, _05273_, _05269_);
  nor (_05275_, _05274_, _05153_);
  nor (_05276_, _05275_, _05267_);
  and (_05278_, _05276_, _05261_);
  and (_05280_, _05108_, _05006_);
  and (_05281_, _05096_, _05091_);
  or (_05282_, _05281_, _05280_);
  and (_05283_, _05102_, _05009_);
  and (_05285_, _05114_, _05027_);
  or (_05286_, _05285_, _05283_);
  or (_05287_, _05286_, _05282_);
  and (_05288_, _05287_, _05241_);
  not (_05289_, _05241_);
  and (_05291_, _05081_, _05009_);
  and (_05293_, _05086_, _05027_);
  or (_05294_, _05293_, _05291_);
  and (_05295_, _05075_, _05006_);
  and (_05296_, _05069_, _05016_);
  or (_05298_, _05296_, _05295_);
  or (_05300_, _05298_, _05294_);
  and (_05301_, _05300_, _05289_);
  nor (_05303_, _05301_, _05288_);
  nor (_05304_, _05303_, _05278_);
  and (_05306_, _05278_, word_in[23]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _05306_, _05304_);
  nor (_05307_, _05122_, _05005_);
  not (_05308_, _05307_);
  nand (_05309_, _05122_, _05005_);
  and (_05310_, _05309_, _05308_);
  not (_05311_, _05310_);
  nor (_05312_, _05051_, _05311_);
  nor (_05313_, _05309_, _04991_);
  and (_05314_, _05309_, _04991_);
  nor (_05316_, _05314_, _05313_);
  nor (_05317_, _05316_, _05310_);
  and (_05318_, _05317_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05319_, _05318_, _05312_);
  nor (_05320_, _05319_, _05143_);
  not (_05321_, _05320_);
  and (_05322_, _05141_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05323_, _05044_, _05311_);
  and (_05324_, _05316_, _05311_);
  and (_05325_, _05324_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05326_, _05317_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05327_, _05326_, _05325_);
  nor (_05328_, _05327_, _05323_);
  nor (_05329_, _05328_, _05153_);
  nor (_05330_, _05329_, _05322_);
  and (_05332_, _05330_, _05321_);
  nor (_05334_, _05311_, _04994_);
  and (_05335_, _05324_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05336_, _05317_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_05337_, _05336_, _05335_);
  nor (_05338_, _05337_, _05334_);
  nor (_05339_, _05338_, _05162_);
  nor (_05340_, _05311_, _05021_);
  and (_05341_, _05317_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05343_, _05341_, _05340_);
  nor (_05344_, _05343_, _05122_);
  and (_05345_, _05307_, _05012_);
  or (_05346_, _05345_, _05344_);
  nor (_05347_, _05346_, _05339_);
  and (_05349_, _05347_, _05332_);
  and (_05350_, _05183_, _05173_);
  and (_05351_, _05178_, _05172_);
  or (_05352_, _05351_, _05350_);
  and (_05354_, _05352_, _05324_);
  and (_05355_, _05197_, _05173_);
  and (_05356_, _05190_, _05172_);
  or (_05357_, _05356_, _05355_);
  and (_05358_, _05357_, _05317_);
  and (_05359_, _05310_, _05091_);
  and (_05361_, _05213_, _05173_);
  and (_05362_, _05207_, _05172_);
  or (_05363_, _05362_, _05361_);
  and (_05364_, _05363_, _05359_);
  and (_05365_, _05227_, _05173_);
  and (_05367_, _05222_, _05172_);
  or (_05368_, _05367_, _05365_);
  and (_05369_, _05314_, _05308_);
  and (_05371_, _05369_, _05368_);
  or (_05372_, _05371_, _05364_);
  or (_05374_, _05372_, _05358_);
  nor (_05375_, _05374_, _05354_);
  nor (_05376_, _05375_, _05349_);
  and (_05377_, _05349_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _05377_, _05376_);
  and (_05380_, _04901_, _23900_);
  and (_05381_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or (_00779_, _05381_, _05380_);
  and (_05383_, _05005_, _04991_);
  or (_05384_, _05383_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_26812_[15], _05384_, _22773_);
  and (_05385_, _05349_, _22773_);
  and (_05387_, _05385_, word_in[31]);
  and (_05388_, _05383_, _05120_);
  and (_05390_, _05385_, _05388_);
  and (_05391_, _05390_, _05387_);
  not (_05392_, _05390_);
  and (_05393_, _05238_, _04991_);
  and (_05394_, _05278_, _22773_);
  and (_05395_, _05394_, _05151_);
  and (_05396_, _05395_, _05393_);
  not (_05398_, _05396_);
  and (_05399_, _05170_, _22773_);
  and (_05400_, _05399_, _05161_);
  and (_05401_, _05400_, _05218_);
  and (_05402_, _05032_, _22773_);
  and (_05403_, _05402_, _04999_);
  nor (_05404_, _05063_, rst);
  and (_05405_, _05404_, _05383_);
  and (_05406_, _05405_, _05403_);
  and (_05407_, _05404_, word_in[7]);
  and (_05408_, _05407_, _05406_);
  nor (_05409_, _05406_, _05104_);
  nor (_05410_, _05409_, _05408_);
  nor (_05411_, _05410_, _05401_);
  and (_05412_, _05401_, word_in[15]);
  or (_05413_, _05412_, _05411_);
  and (_05414_, _05413_, _05398_);
  and (_05415_, _05394_, word_in[23]);
  and (_05416_, _05415_, _05396_);
  or (_05417_, _05416_, _05414_);
  and (_05418_, _05417_, _05392_);
  or (_26820_[7], _05418_, _05391_);
  or (_05419_, _05324_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_26830_, _05419_, _22773_);
  or (_05421_, _25931_, _25888_);
  or (_05422_, _25892_, _25889_);
  or (_05423_, _25929_, _25914_);
  or (_05424_, _05423_, _05422_);
  or (_05425_, _05424_, _05421_);
  not (_05426_, _25906_);
  and (_05428_, _24541_, _24503_);
  and (_05429_, _05428_, _24669_);
  and (_05430_, _05429_, _25887_);
  nor (_05431_, _05430_, _05426_);
  nand (_05432_, _05431_, _25878_);
  not (_05433_, _25900_);
  and (_05434_, _25849_, _24639_);
  or (_05435_, _05434_, _05433_);
  or (_05436_, _05435_, _05432_);
  or (_05437_, _05436_, _05425_);
  and (_05439_, _25924_, _24677_);
  or (_05441_, _05439_, _24710_);
  and (_05442_, _26167_, _24669_);
  or (_05443_, _05442_, _25902_);
  or (_05444_, _05443_, _05441_);
  or (_05445_, _05444_, _05437_);
  and (_05447_, _05445_, _01886_);
  and (_05448_, _25850_, _24733_);
  not (_05449_, _25859_);
  and (_05450_, _05449_, _04966_);
  or (_05452_, _05442_, _05434_);
  and (_05453_, _05452_, _24733_);
  or (_05454_, _05453_, _05450_);
  or (_05455_, _05454_, _05448_);
  and (_05456_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_05457_, _05456_, _05455_);
  and (_05458_, _05457_, _22773_);
  or (_26839_[0], _05458_, _05447_);
  and (_05459_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_05460_, _05459_, _05454_);
  and (_05462_, _05460_, _22773_);
  and (_05463_, _05429_, _24690_);
  or (_05464_, _05463_, _24725_);
  or (_05466_, _05464_, _25921_);
  and (_05467_, _25904_, _24670_);
  or (_05468_, _05467_, _24691_);
  or (_05470_, _05468_, _05466_);
  or (_05471_, _05470_, _05452_);
  and (_05473_, _05471_, _01886_);
  or (_26839_[1], _05473_, _05462_);
  not (_05474_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05475_, _05028_, _04991_);
  nand (_05477_, _05475_, _05474_);
  or (_05478_, _05477_, _05240_);
  and (_26812_[1], _05478_, _22773_);
  and (_05479_, _05359_, _05161_);
  nor (_05480_, _05479_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_05481_, _05141_);
  and (_05482_, _05475_, _05481_);
  nand (_05484_, _05482_, _05480_);
  and (_26812_[2], _05484_, _22773_);
  and (_05485_, _02531_, _23751_);
  and (_05486_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  or (_00919_, _05486_, _05485_);
  and (_05487_, _01709_, _23751_);
  and (_05489_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_00936_, _05489_, _05487_);
  and (_05491_, _02531_, _23900_);
  and (_05492_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  or (_00944_, _05492_, _05491_);
  not (_05494_, _05135_);
  and (_05496_, _05359_, _05123_);
  or (_05498_, _05005_, _04991_);
  or (_05499_, _05498_, _05161_);
  and (_05500_, _05499_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05501_, _05500_, _05496_);
  and (_05502_, _05501_, _05494_);
  and (_05504_, _05027_, _05012_);
  or (_05505_, _05504_, _05479_);
  or (_05507_, _05505_, _05502_);
  and (_05508_, _05507_, _05482_);
  not (_05509_, _05475_);
  or (_05510_, _05504_, _05501_);
  and (_05511_, _05510_, _05141_);
  or (_05512_, _05511_, _05509_);
  or (_05513_, _05512_, _05508_);
  and (_26812_[3], _05513_, _22773_);
  and (_05514_, _02531_, _24027_);
  and (_05515_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  or (_00954_, _05515_, _05514_);
  nand (_05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _22773_);
  nor (_01000_, _05516_, t2ex_i);
  and (_05517_, _05130_, _05120_);
  or (_05518_, _05517_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05519_, _05518_, _05498_);
  or (_05521_, _05519_, _05496_);
  and (_05523_, _05521_, _05494_);
  and (_05524_, _05518_, _05141_);
  and (_05526_, _05151_, _05359_);
  and (_05527_, _05307_, _05091_);
  and (_05529_, _05527_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_05530_, _05529_, _05526_);
  or (_05532_, _05530_, _05479_);
  or (_05534_, _05532_, _05524_);
  or (_05535_, _05534_, _05523_);
  and (_26812_[4], _05535_, _22773_);
  and (_05536_, _05498_, _05481_);
  not (_05537_, _05239_);
  or (_05538_, _05517_, _05496_);
  or (_05540_, _05538_, _05537_);
  and (_05541_, _05540_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05543_, _05509_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05544_, _05151_, _05130_);
  and (_05546_, _05479_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05547_, _05546_, _05544_);
  or (_05549_, _05547_, _05543_);
  or (_05550_, _05549_, _05541_);
  or (_05552_, _05129_, _05313_);
  and (_05553_, _05552_, _05550_);
  and (_05555_, _05359_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05556_, _05555_, _05517_);
  or (_05557_, _05556_, _05553_);
  and (_05559_, _05557_, _05536_);
  and (_05561_, _05550_, _05141_);
  and (_05563_, _05526_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05564_, _05527_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05566_, _05564_, _05479_);
  or (_05567_, _05566_, _05563_);
  or (_05569_, _05567_, _05496_);
  or (_05570_, _05569_, _05561_);
  or (_05571_, _05570_, _05559_);
  and (_26812_[5], _05571_, _22773_);
  nor (_05573_, t2_i, rst);
  and (_01097_, _05573_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and (_01107_, t2_i, _22773_);
  nand (_05575_, _02481_, _23976_);
  not (_05576_, _02473_);
  and (_05577_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_05578_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_05579_, _05578_, _05577_);
  or (_05582_, _05579_, _02481_);
  and (_05584_, _05582_, _05576_);
  and (_05585_, _05584_, _05575_);
  and (_05586_, _02473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_05587_, _05586_, _05585_);
  and (_01111_, _05587_, _22773_);
  and (_01115_, t2ex_i, _22773_);
  and (_05588_, _05538_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05589_, _05588_, _05544_);
  nand (_05590_, _05005_, _04985_);
  nand (_05591_, _05239_, _05590_);
  and (_05592_, _05161_, _05130_);
  or (_05593_, _05592_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_05594_, _05593_, _05591_);
  and (_05595_, _05594_, _05537_);
  or (_05596_, _05595_, _05589_);
  and (_05597_, _05596_, _05552_);
  and (_05598_, _05593_, _05141_);
  and (_05599_, _05479_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_05601_, _05509_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05602_, _05601_, _05496_);
  or (_05604_, _05602_, _05599_);
  or (_05605_, _05604_, _05517_);
  or (_05606_, _05605_, _05598_);
  or (_05607_, _05606_, _05597_);
  and (_26812_[6], _05607_, _22773_);
  not (_05609_, _02477_);
  or (_05610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_05611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_05613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _05611_);
  and (_05615_, _05613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_05616_, _05615_, _05610_);
  and (_05617_, _02472_, _23209_);
  and (_05618_, _02472_, _24191_);
  nor (_05619_, _05618_, _05617_);
  and (_05620_, _05619_, _05616_);
  and (_05621_, _05620_, _05609_);
  not (_05622_, _05621_);
  and (_05623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_05624_, _05623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_05625_, _05624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_05626_, _05625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_05627_, _05626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_05628_, _05627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_05629_, _05628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_05630_, _05629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_05631_, _05630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_05632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_05633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_05634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_05635_, _05634_, _05633_);
  and (_05636_, _05635_, _05632_);
  and (_05637_, _05636_, _05631_);
  or (_05639_, _05637_, _05622_);
  or (_05641_, _05621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_05643_, _05641_, _22773_);
  and (_01126_, _05643_, _05639_);
  nand (_05644_, _02473_, _23976_);
  or (_05645_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_05646_, _02482_);
  or (_05647_, _05646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_05648_, _05647_, _05645_);
  or (_05650_, _05648_, _02473_);
  and (_05651_, _05650_, _22773_);
  and (_01131_, _05651_, _05644_);
  and (_05652_, _05618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_05653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_05655_, _02476_, _05653_);
  nor (_05656_, _05655_, _05609_);
  not (_05657_, _02478_);
  and (_05658_, _05616_, _05657_);
  and (_05659_, _05658_, _05637_);
  and (_05660_, _05659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_05661_, _05660_, _05656_);
  and (_05662_, _05631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_05663_, _05662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_05664_, _05663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_05665_, _05616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_05667_, _05665_, _05664_);
  and (_05668_, _05667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand (_05670_, _05668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_05671_, _05668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_05672_, _05671_, _05670_);
  or (_05673_, _05672_, _05661_);
  not (_05674_, _05656_);
  or (_05675_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_05676_, _05675_, _05619_);
  and (_05677_, _05676_, _05673_);
  or (_05678_, _05677_, _05652_);
  not (_05679_, _05617_);
  nor (_05680_, _05679_, _23976_);
  or (_05681_, _05680_, _05678_);
  and (_01134_, _05681_, _22773_);
  not (_05682_, _05618_);
  nor (_05683_, _05682_, _23976_);
  or (_05684_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_05685_, _05616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_05686_, _05628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_05687_, _05629_, _05616_);
  and (_05688_, _05687_, _05686_);
  and (_05689_, _05657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_05691_, _05689_, _05637_);
  or (_05692_, _05691_, _05688_);
  and (_05693_, _05692_, _05685_);
  or (_05694_, _05693_, _05656_);
  and (_05696_, _05694_, _05684_);
  and (_05697_, _05696_, _05682_);
  or (_05698_, _05697_, _05617_);
  or (_05699_, _05698_, _05683_);
  or (_05700_, _05679_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_05702_, _05700_, _22773_);
  and (_01138_, _05702_, _05699_);
  or (_05704_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_05705_, _26279_, _24423_);
  or (_05706_, _05705_, _05704_);
  nand (_05708_, _03241_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_05709_, _05708_, _05705_);
  or (_05710_, _05709_, _03242_);
  and (_05711_, _05710_, _05706_);
  and (_05713_, _02472_, _24406_);
  or (_05714_, _05713_, _05711_);
  nand (_05716_, _05713_, _23976_);
  and (_05718_, _05716_, _22773_);
  and (_01147_, _05718_, _05714_);
  not (_05719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor (_05720_, _05619_, _05719_);
  and (_05721_, _05655_, _02477_);
  and (_05723_, _05721_, _05637_);
  and (_05724_, _05723_, _05620_);
  or (_05725_, _05724_, _05720_);
  and (_01150_, _05725_, _22773_);
  and (_05726_, _23909_, _23444_);
  and (_05727_, _05726_, _23751_);
  not (_05728_, _05726_);
  and (_05730_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_27103_, _05730_, _05727_);
  and (_05731_, _24274_, _23891_);
  and (_05732_, _05731_, _23715_);
  not (_05733_, _05731_);
  and (_05734_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or (_01165_, _05734_, _05732_);
  and (_05736_, _05731_, _23693_);
  and (_05737_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or (_27242_, _05737_, _05736_);
  and (_05738_, _05731_, _23751_);
  and (_05739_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or (_01182_, _05739_, _05738_);
  and (_05740_, _05726_, _23715_);
  and (_05741_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_01184_, _05741_, _05740_);
  and (_05742_, _05726_, _23920_);
  and (_05743_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_01190_, _05743_, _05742_);
  or (_05744_, _05517_, _05240_);
  or (_05745_, _05744_, _05241_);
  and (_05746_, _04991_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05747_, _05019_, _05006_);
  and (_05748_, _05130_, _05033_);
  or (_05749_, _05748_, _05131_);
  or (_05751_, _05749_, _05747_);
  or (_05752_, _05751_, _05746_);
  and (_05754_, _05752_, _05745_);
  and (_05755_, _05019_, _05040_);
  and (_05756_, _05517_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_05758_, _05756_, _05544_);
  or (_05759_, _05758_, _05755_);
  or (_05761_, _05759_, _05754_);
  and (_26812_[7], _05761_, _22773_);
  or (_05763_, _05576_, _23205_);
  and (_05765_, _05646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_05766_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_05768_, _05766_, _05765_);
  or (_05769_, _05768_, _02473_);
  and (_05770_, _05769_, _22773_);
  and (_01214_, _05770_, _05763_);
  and (_05771_, _26228_, _25876_);
  and (_05772_, _05771_, _24566_);
  or (_05773_, _05772_, _04210_);
  or (_05775_, _05773_, _05434_);
  or (_05776_, _04945_, _24706_);
  or (_05778_, _04949_, _04943_);
  or (_05779_, _05778_, _05776_);
  or (_05780_, _05779_, _05775_);
  and (_05781_, _04214_, _24670_);
  or (_05782_, _05781_, _26253_);
  and (_05783_, _24639_, _24704_);
  and (_05784_, _04213_, _24566_);
  or (_05785_, _05784_, _05783_);
  or (_05786_, _05785_, _05782_);
  and (_05787_, _04919_, _25887_);
  or (_05788_, _05463_, _05442_);
  or (_05790_, _05788_, _05787_);
  and (_05791_, _26231_, _05428_);
  or (_05793_, _05791_, _24693_);
  or (_05795_, _04923_, _04232_);
  or (_05796_, _05795_, _05793_);
  or (_05797_, _05796_, _05790_);
  or (_05798_, _05797_, _05786_);
  or (_05799_, _04228_, _26229_);
  or (_05801_, _04920_, _25857_);
  or (_05802_, _05801_, _05799_);
  or (_05803_, _05802_, _04938_);
  and (_05804_, _04214_, _24669_);
  or (_05805_, _03594_, _25858_);
  or (_05806_, _05805_, _01885_);
  or (_05807_, _05806_, _05804_);
  or (_05808_, _05807_, _05803_);
  or (_05809_, _05808_, _05798_);
  or (_05810_, _05809_, _05780_);
  and (_05811_, _05810_, _23760_);
  and (_05812_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_05813_, _04975_, _25860_);
  or (_05814_, _05813_, _05812_);
  or (_05815_, _05814_, _05811_);
  and (_26840_[0], _05815_, _22773_);
  not (_05816_, _05498_);
  or (_05817_, _05359_, _05317_);
  nor (_05819_, _05817_, _05527_);
  or (_05820_, _05819_, _05816_);
  and (_05821_, _05820_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05822_, _05307_, _04991_);
  and (_05823_, _05130_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_05824_, _05132_, _05122_);
  and (_05825_, _05824_, _05823_);
  or (_05826_, _05544_, _05131_);
  or (_05827_, _05826_, _05825_);
  or (_05828_, _05827_, _05592_);
  or (_05830_, _05828_, _05822_);
  or (_05831_, _05830_, _05821_);
  and (_26812_[8], _05831_, _22773_);
  and (_05832_, _05726_, _23983_);
  and (_05833_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_01257_, _05833_, _05832_);
  and (_05834_, _24068_, _23891_);
  and (_05835_, _05834_, _23920_);
  not (_05836_, _05834_);
  and (_05837_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_01263_, _05837_, _05835_);
  and (_05838_, _24053_, _23910_);
  and (_05840_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_01277_, _05840_, _05838_);
  and (_05841_, _05239_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05842_, _05129_, _05308_);
  and (_05844_, _05369_, _05151_);
  nor (_05846_, _05239_, _05024_);
  or (_05847_, _05846_, _05844_);
  and (_05849_, _05847_, _05842_);
  or (_05850_, _05849_, _05822_);
  and (_05851_, _05016_, _05091_);
  and (_05853_, _05847_, _05141_);
  or (_05854_, _05853_, _05851_);
  or (_05856_, _05854_, _05850_);
  or (_05858_, _05856_, _05841_);
  and (_26812_[9], _05858_, _22773_);
  and (_05859_, _24145_, _23909_);
  and (_05860_, _05859_, _24053_);
  not (_05862_, _05859_);
  and (_05863_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  or (_01329_, _05863_, _05860_);
  and (_05864_, _05731_, _24027_);
  and (_05866_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or (_27243_, _05866_, _05864_);
  and (_05867_, _05859_, _23693_);
  and (_05868_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  or (_01334_, _05868_, _05867_);
  and (_05869_, _05731_, _23920_);
  and (_05870_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or (_01337_, _05870_, _05869_);
  and (_05871_, _05859_, _23900_);
  and (_05872_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  or (_01354_, _05872_, _05871_);
  and (_05873_, _05731_, _23900_);
  and (_05874_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or (_01377_, _05874_, _05873_);
  and (_05876_, _05859_, _23920_);
  and (_05877_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  or (_01392_, _05877_, _05876_);
  and (_05878_, _23924_, _23909_);
  and (_05880_, _05878_, _23751_);
  not (_05881_, _05878_);
  and (_05882_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_01398_, _05882_, _05880_);
  and (_05883_, _23905_, _23891_);
  and (_05885_, _05883_, _23715_);
  not (_05886_, _05883_);
  and (_05887_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_01402_, _05887_, _05885_);
  and (_05888_, _05314_, _05161_);
  not (_05889_, _05125_);
  and (_05890_, _05889_, _05053_);
  or (_05891_, _05890_, _05888_);
  and (_05893_, _05238_, _05091_);
  and (_05894_, _05893_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05895_, _05509_, _05592_);
  and (_05896_, _05895_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05897_, _05896_, _05894_);
  or (_05898_, _05897_, _05131_);
  or (_05900_, _05898_, _05844_);
  or (_05902_, _05900_, _05891_);
  or (_05904_, _05902_, _05822_);
  and (_26812_[10], _05904_, _22773_);
  and (_05906_, _05883_, _23900_);
  and (_05908_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_27240_, _05908_, _05906_);
  and (_05909_, _02403_, _24053_);
  and (_05910_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_01424_, _05910_, _05909_);
  and (_05912_, _05314_, _05123_);
  and (_05913_, _05383_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05914_, _05913_, _05912_);
  and (_05915_, _05202_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05916_, _05173_, _05359_);
  and (_05917_, _05916_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05918_, _05131_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05919_, _04991_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05920_, _05919_, _05307_);
  or (_05921_, _05920_, _05918_);
  or (_05922_, _05921_, _05917_);
  or (_05923_, _05922_, _05888_);
  or (_05924_, _05923_, _05915_);
  or (_05925_, _05924_, _05844_);
  or (_05926_, _05925_, _05914_);
  and (_26812_[11], _05926_, _22773_);
  or (_05927_, _05778_, _05773_);
  or (_05929_, _05927_, _05776_);
  and (_05930_, _26231_, _24696_);
  or (_05932_, _05930_, _24693_);
  or (_05933_, _25902_, _25858_);
  or (_05934_, _05933_, _05932_);
  or (_05935_, _24715_, _24699_);
  and (_05936_, _05935_, _24648_);
  or (_05937_, _05936_, _25918_);
  or (_05938_, _05937_, _05934_);
  and (_05939_, _04919_, _24690_);
  or (_05941_, _05430_, _04231_);
  or (_05943_, _05941_, _05939_);
  or (_05944_, _05943_, _24684_);
  or (_05946_, _05944_, _05938_);
  or (_05947_, _05946_, _05803_);
  or (_05948_, _05947_, _05929_);
  and (_05949_, _05948_, _23760_);
  and (_05950_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_05951_, _05950_, _05813_);
  or (_05952_, _05951_, _05949_);
  and (_26840_[1], _05952_, _22773_);
  and (_05953_, _05878_, _23715_);
  and (_05955_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_01507_, _05955_, _05953_);
  and (_05956_, _01735_, _24341_);
  nand (_05957_, _05956_, _23681_);
  or (_05958_, _05956_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_05959_, _05958_, _01739_);
  and (_05960_, _05959_, _05957_);
  nor (_05961_, _01739_, _23976_);
  or (_05962_, _05961_, _05960_);
  and (_01519_, _05962_, _22773_);
  or (_05963_, _02331_, _02271_);
  and (_05965_, _05963_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_05966_, _05965_, _02296_);
  and (_01521_, _05966_, _22773_);
  nor (_01523_, _04172_, rst);
  and (_05967_, _05878_, _23900_);
  and (_05968_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_01540_, _05968_, _05967_);
  nor (_05969_, _05120_, _05041_);
  and (_05971_, _05969_, _05383_);
  and (_05973_, _04999_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05974_, _05973_, _05359_);
  nand (_05976_, _05475_, _05308_);
  and (_05977_, _05976_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05978_, _05130_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05979_, _05978_, _05369_);
  or (_05980_, _05979_, _05977_);
  or (_05982_, _05980_, _05974_);
  or (_05983_, _05982_, _05971_);
  and (_26812_[12], _05983_, _22773_);
  and (_05985_, _01749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_05987_, _01751_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_01547_, _05987_, _05985_);
  or (_05988_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_05989_, _05988_, _22773_);
  and (_05990_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_05991_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_05992_, _05991_, rxd_i);
  or (_05993_, _05992_, _05990_);
  and (_05994_, _05993_, _02186_);
  and (_05995_, _02209_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_05996_, _05995_, _05994_);
  and (_05997_, _02196_, rxd_i);
  or (_05998_, _05997_, _02207_);
  or (_05999_, _05998_, _05996_);
  and (_01549_, _05999_, _05989_);
  and (_06000_, _05878_, _23983_);
  and (_06001_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_01576_, _06001_, _06000_);
  and (_06003_, _05834_, _24027_);
  and (_06004_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_01581_, _06004_, _06003_);
  and (_06005_, _25175_, _23938_);
  and (_06006_, _06005_, _24053_);
  not (_06007_, _06005_);
  and (_06008_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_01593_, _06008_, _06006_);
  and (_06010_, _02283_, _02182_);
  and (_06011_, _02273_, _06010_);
  nand (_06012_, _06011_, _02298_);
  or (_06013_, _06011_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_06014_, _06013_, _22773_);
  and (_01596_, _06014_, _06012_);
  or (_06015_, _04266_, rxd_i);
  nand (_06016_, _06015_, _02190_);
  or (_06017_, _02191_, _02178_);
  and (_06018_, _06017_, _06016_);
  or (_06019_, _02195_, _02189_);
  or (_06020_, _06019_, _02179_);
  or (_06021_, _06020_, _06018_);
  and (_01598_, _06021_, _01751_);
  or (_06022_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_06023_, _06022_, _22773_);
  nand (_06024_, _01959_, _23976_);
  and (_01600_, _06024_, _06023_);
  nand (_06025_, _01983_, _01979_);
  and (_06026_, _06025_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_06027_, _06026_, _04194_);
  nor (_06028_, _01977_, _04195_);
  and (_06029_, _06028_, _06027_);
  or (_06030_, _06029_, _02142_);
  nand (_06031_, _06030_, _22773_);
  nor (_01603_, _06031_, _01970_);
  or (_06032_, _05393_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_26812_[13], _06032_, _22773_);
  and (_06033_, _06005_, _23693_);
  and (_06034_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_01623_, _06034_, _06033_);
  and (_06035_, _06005_, _23715_);
  and (_06036_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_01649_, _06036_, _06035_);
  and (_06037_, _01745_, _23751_);
  and (_06039_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or (_26913_, _06039_, _06037_);
  and (_06041_, _06005_, _24027_);
  and (_06042_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_27115_, _06042_, _06041_);
  or (_06043_, _05218_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_26812_[14], _06043_, _22773_);
  and (_06044_, _24901_, _23900_);
  and (_06045_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_01690_, _06045_, _06044_);
  and (_06047_, _04207_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_06048_, _26228_, _25849_);
  or (_06049_, _04935_, _06048_);
  and (_06051_, _25924_, _24687_);
  or (_06052_, _06051_, _04945_);
  or (_06053_, _06052_, _06049_);
  and (_06054_, _24712_, _24648_);
  or (_06055_, _25876_, _25849_);
  and (_06057_, _06055_, _24690_);
  or (_06058_, _06057_, _06054_);
  or (_06059_, _06058_, _06053_);
  or (_06060_, _24724_, _24687_);
  and (_06061_, _06060_, _26231_);
  or (_06063_, _25914_, _24693_);
  nor (_06065_, _06063_, _06061_);
  nand (_06066_, _06065_, _25882_);
  or (_06068_, _25888_, _24675_);
  or (_06069_, _06068_, _05433_);
  or (_06070_, _06069_, _06066_);
  or (_06071_, _06070_, _06059_);
  and (_06072_, _04949_, _24676_);
  and (_06073_, _06072_, _24669_);
  and (_06074_, _25898_, _24565_);
  nor (_06076_, _06074_, _04210_);
  nand (_06077_, _06076_, _02542_);
  or (_06079_, _06077_, _06073_);
  and (_06080_, _04949_, _24503_);
  or (_06081_, _04942_, _04214_);
  or (_06082_, _06081_, _04944_);
  or (_06084_, _06082_, _06080_);
  and (_06085_, _06084_, _24669_);
  or (_06086_, _06085_, _06079_);
  or (_06087_, _06086_, _06071_);
  and (_06088_, _06087_, _01886_);
  or (_26841_[0], _06088_, _06047_);
  and (_06090_, _24901_, _23920_);
  and (_06091_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_01696_, _06091_, _06090_);
  and (_06093_, _04207_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_06094_, _04935_, _25891_);
  and (_06095_, _24699_, _24690_);
  or (_06096_, _06095_, _05771_);
  or (_06097_, _06096_, _06094_);
  or (_06098_, _04222_, _24647_);
  or (_06100_, _06098_, _24691_);
  or (_06102_, _06100_, _24675_);
  or (_06103_, _06102_, _06097_);
  or (_06104_, _04232_, _25892_);
  or (_06105_, _06104_, _25879_);
  or (_06106_, _06105_, _03593_);
  or (_06107_, _06106_, _06103_);
  or (_06108_, _04943_, _24706_);
  or (_06109_, _06108_, _05782_);
  or (_06111_, _06109_, _05807_);
  and (_06112_, _06080_, _24669_);
  or (_06113_, _06112_, _06073_);
  or (_06115_, _06113_, _06111_);
  or (_06116_, _06115_, _06107_);
  or (_06117_, _25858_, _24646_);
  nor (_06118_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and (_06120_, _06118_, _06117_);
  and (_06121_, _06120_, _06116_);
  or (_26842_[0], _06121_, _06093_);
  and (_06122_, _05834_, _23983_);
  and (_06123_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_01706_, _06123_, _06122_);
  and (_06124_, _23900_, _23454_);
  and (_06126_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or (_01708_, _06126_, _06124_);
  and (_06128_, _02455_, _23751_);
  and (_06130_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or (_01710_, _06130_, _06128_);
  or (_06131_, _26240_, _25881_);
  or (_06132_, _04210_, _25858_);
  or (_06133_, _05771_, _04941_);
  or (_06134_, _06133_, _06132_);
  or (_06135_, _06134_, _06080_);
  or (_06136_, _06135_, _06131_);
  or (_06137_, _05799_, _24694_);
  or (_06138_, _03597_, _24725_);
  or (_06139_, _06138_, _06052_);
  nor (_06140_, _06139_, _06137_);
  nand (_06141_, _06140_, _03595_);
  or (_06142_, _05421_, _04932_);
  or (_06143_, _06142_, _06048_);
  or (_06144_, _06054_, _25875_);
  and (_06145_, _24724_, _24615_);
  or (_06146_, _06145_, _26232_);
  or (_06147_, _06146_, _04920_);
  or (_06148_, _06147_, _06144_);
  or (_06149_, _06148_, _06143_);
  or (_06150_, _06149_, _06141_);
  or (_06152_, _06150_, _06136_);
  and (_06154_, _06152_, _06120_);
  and (_06155_, _04207_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or (_26842_[1], _06155_, _06154_);
  and (_06156_, _02829_, _24053_);
  and (_06157_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or (_27122_, _06157_, _06156_);
  and (_06158_, _02829_, _23983_);
  and (_06159_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or (_01763_, _06159_, _06158_);
  and (_06160_, _04033_, _23751_);
  and (_06162_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or (_27124_, _06162_, _06160_);
  and (_06163_, _02455_, _24053_);
  and (_06164_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or (_01828_, _06164_, _06163_);
  and (_06165_, _01709_, _23983_);
  and (_06167_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_01845_, _06167_, _06165_);
  and (_06168_, _04033_, _23920_);
  and (_06169_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or (_01853_, _06169_, _06168_);
  and (_06171_, _02350_, _23900_);
  and (_06172_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_01884_, _06172_, _06171_);
  and (_06173_, _24389_, _23983_);
  and (_06174_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_01899_, _06174_, _06173_);
  and (_06175_, _02798_, _23920_);
  and (_06177_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_01912_, _06177_, _06175_);
  not (_06178_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_06179_, _05404_, _04999_);
  nor (_06180_, _06179_, _05402_);
  and (_06181_, _05404_, _05498_);
  not (_06182_, _06181_);
  and (_06183_, _06182_, _06180_);
  and (_06184_, _06183_, _05404_);
  nor (_06186_, _06184_, _06178_);
  and (_06187_, _05399_, _05141_);
  and (_06188_, _05404_, word_in[0]);
  and (_06189_, _06188_, _06183_);
  or (_06190_, _06189_, _06187_);
  or (_06191_, _06190_, _06186_);
  and (_06192_, _05383_, _05161_);
  and (_06194_, _05394_, _06192_);
  not (_06195_, _06194_);
  not (_06196_, _06187_);
  or (_06197_, _06196_, word_in[8]);
  and (_06198_, _06197_, _06195_);
  and (_06199_, _06198_, _06191_);
  and (_06200_, _05151_, _05383_);
  and (_06201_, _05385_, _06200_);
  and (_06202_, _06194_, word_in[16]);
  or (_06203_, _06202_, _06201_);
  or (_06204_, _06203_, _06199_);
  not (_06205_, _06201_);
  or (_06206_, _06205_, word_in[24]);
  and (_26814_[0], _06206_, _06204_);
  and (_06207_, _05385_, word_in[25]);
  and (_06208_, _06207_, _06200_);
  not (_06209_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_06210_, _06184_, _06209_);
  and (_06212_, _05404_, word_in[1]);
  and (_06213_, _06212_, _06183_);
  or (_06214_, _06213_, _06210_);
  and (_06215_, _06214_, _06196_);
  and (_06216_, _06187_, word_in[9]);
  or (_06217_, _06216_, _06215_);
  or (_06219_, _06217_, _06194_);
  or (_06220_, _06195_, word_in[17]);
  and (_06221_, _06220_, _06205_);
  and (_06222_, _06221_, _06219_);
  or (_26814_[1], _06222_, _06208_);
  and (_06223_, _02798_, _23715_);
  and (_06224_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_27125_, _06224_, _06223_);
  not (_06225_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_06226_, _06184_, _06225_);
  and (_06227_, _05404_, word_in[2]);
  and (_06228_, _06227_, _06183_);
  or (_06229_, _06228_, _06226_);
  or (_06230_, _06229_, _06187_);
  or (_06231_, _06196_, word_in[10]);
  and (_06232_, _06231_, _06195_);
  and (_06233_, _06232_, _06230_);
  and (_06234_, _06194_, word_in[18]);
  or (_06235_, _06234_, _06233_);
  and (_06236_, _06235_, _06205_);
  and (_06237_, _06201_, word_in[26]);
  or (_26814_[2], _06237_, _06236_);
  not (_06238_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_06239_, _06184_, _06238_);
  and (_06240_, _05404_, word_in[3]);
  and (_06241_, _06240_, _06183_);
  or (_06242_, _06241_, _06239_);
  and (_06243_, _06242_, _06196_);
  and (_06244_, _06187_, word_in[11]);
  or (_06245_, _06244_, _06243_);
  and (_06246_, _06245_, _06195_);
  and (_06247_, _05394_, word_in[19]);
  and (_06249_, _06247_, _06192_);
  or (_06250_, _06249_, _06246_);
  and (_06251_, _06250_, _06205_);
  and (_06252_, _06201_, word_in[27]);
  or (_26814_[3], _06252_, _06251_);
  and (_06253_, _25175_, _23444_);
  and (_06254_, _06253_, _23751_);
  not (_06255_, _06253_);
  and (_06256_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or (_01930_, _06256_, _06254_);
  not (_06257_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_06258_, _06184_, _06257_);
  and (_06259_, _05404_, word_in[4]);
  and (_06260_, _06259_, _06183_);
  or (_06261_, _06260_, _06258_);
  or (_06262_, _06261_, _06187_);
  or (_06263_, _06196_, word_in[12]);
  and (_06264_, _06263_, _06195_);
  and (_06265_, _06264_, _06262_);
  and (_06266_, _06194_, word_in[20]);
  or (_06268_, _06266_, _06265_);
  and (_06269_, _06268_, _06205_);
  and (_06271_, _06201_, word_in[28]);
  or (_26814_[4], _06271_, _06269_);
  and (_06273_, _05385_, word_in[29]);
  and (_06274_, _06273_, _06200_);
  not (_06275_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_06276_, _06184_, _06275_);
  and (_06278_, _05404_, word_in[5]);
  and (_06279_, _06278_, _06183_);
  or (_06281_, _06279_, _06187_);
  or (_06282_, _06281_, _06276_);
  or (_06284_, _06196_, word_in[13]);
  and (_06285_, _06284_, _06195_);
  and (_06286_, _06285_, _06282_);
  and (_06287_, _06194_, word_in[21]);
  or (_06288_, _06287_, _06286_);
  and (_06289_, _06288_, _06205_);
  or (_26814_[5], _06289_, _06274_);
  and (_06290_, _06194_, word_in[22]);
  not (_06291_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_06292_, _06184_, _06291_);
  and (_06294_, _05404_, word_in[6]);
  and (_06295_, _06294_, _06183_);
  or (_06296_, _06295_, _06292_);
  or (_06297_, _06296_, _06187_);
  or (_06298_, _06196_, word_in[14]);
  and (_06299_, _06298_, _06195_);
  and (_06300_, _06299_, _06297_);
  or (_06301_, _06300_, _06290_);
  and (_06302_, _06301_, _06205_);
  and (_06303_, _06201_, word_in[30]);
  or (_26814_[6], _06303_, _06302_);
  or (_06304_, _06051_, _04941_);
  or (_06305_, _03594_, _25914_);
  nor (_06306_, _06305_, _06304_);
  nand (_06307_, _06306_, _02542_);
  or (_06308_, _06142_, _06072_);
  or (_06309_, _06308_, _06307_);
  or (_06310_, _25902_, _24691_);
  or (_06312_, _06138_, _06049_);
  or (_06313_, _06312_, _06310_);
  or (_06314_, _06313_, _06148_);
  or (_06315_, _06314_, _06309_);
  and (_06316_, _06315_, _23760_);
  and (_06317_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06318_, _25857_, _22781_);
  or (_06319_, _06318_, _06317_);
  or (_06320_, _06319_, _06316_);
  and (_26842_[2], _06320_, _22773_);
  and (_06321_, _06194_, word_in[23]);
  or (_06322_, _06196_, word_in[15]);
  and (_06323_, _06322_, _06195_);
  and (_06324_, _06184_, word_in[7]);
  nor (_06325_, _06184_, _05180_);
  or (_06326_, _06325_, _06324_);
  or (_06327_, _06326_, _06187_);
  and (_06328_, _06327_, _06323_);
  or (_06329_, _06328_, _06321_);
  and (_06330_, _06329_, _06205_);
  and (_06331_, _06201_, word_in[31]);
  or (_26814_[7], _06331_, _06330_);
  and (_06332_, _06253_, _23920_);
  and (_06334_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or (_01950_, _06334_, _06332_);
  and (_06335_, _02794_, _24027_);
  and (_06336_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or (_01956_, _06336_, _06335_);
  and (_06337_, _04033_, _23983_);
  and (_06338_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or (_01968_, _06338_, _06337_);
  and (_06339_, _02789_, _23751_);
  and (_06341_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_01973_, _06341_, _06339_);
  and (_06342_, _02789_, _23983_);
  and (_06343_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_01985_, _06343_, _06342_);
  and (_06344_, _02853_, _24053_);
  and (_06345_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or (_01989_, _06345_, _06344_);
  and (_06347_, _02779_, _23920_);
  and (_06348_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_01993_, _06348_, _06347_);
  and (_06349_, _05385_, _05161_);
  and (_06350_, _06349_, _05324_);
  and (_06351_, _05399_, _05120_);
  and (_06352_, _06351_, _05135_);
  not (_06353_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_06354_, _05402_, _05001_);
  and (_06355_, _06354_, _06182_);
  nor (_06356_, _06355_, _06353_);
  and (_06357_, _06355_, _06188_);
  nor (_06358_, _06357_, _06356_);
  nor (_06360_, _06358_, _06352_);
  and (_06361_, _05394_, _05123_);
  and (_06362_, _06361_, _05242_);
  and (_06363_, _06352_, word_in[8]);
  or (_06364_, _06363_, _06362_);
  or (_06365_, _06364_, _06360_);
  not (_06367_, _06362_);
  or (_06368_, _06367_, word_in[16]);
  and (_06369_, _06368_, _06365_);
  or (_06370_, _06369_, _06350_);
  not (_06372_, _06350_);
  or (_06373_, _06372_, word_in[24]);
  and (_26821_[0], _06373_, _06370_);
  not (_06376_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_06377_, _06355_, _06376_);
  and (_06378_, _06355_, _06212_);
  nor (_06379_, _06378_, _06377_);
  nor (_06380_, _06379_, _06352_);
  and (_06381_, _06352_, word_in[9]);
  or (_06383_, _06381_, _06362_);
  or (_06384_, _06383_, _06380_);
  or (_06385_, _06367_, word_in[17]);
  and (_06386_, _06385_, _06384_);
  or (_06387_, _06386_, _06350_);
  or (_06388_, _06372_, word_in[25]);
  and (_26821_[1], _06388_, _06387_);
  and (_06389_, _04767_, _24053_);
  and (_06390_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_02002_, _06390_, _06389_);
  not (_06391_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_06392_, _06355_, _06391_);
  and (_06393_, _06355_, _06227_);
  nor (_06394_, _06393_, _06392_);
  nor (_06395_, _06394_, _06352_);
  and (_06396_, _06352_, word_in[10]);
  or (_06397_, _06396_, _06362_);
  or (_06398_, _06397_, _06395_);
  or (_06399_, _06367_, word_in[18]);
  and (_06400_, _06399_, _06398_);
  or (_06401_, _06400_, _06350_);
  or (_06402_, _06372_, word_in[26]);
  and (_26821_[2], _06402_, _06401_);
  or (_06403_, _06367_, word_in[19]);
  not (_06404_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_06405_, _06355_, _06404_);
  and (_06406_, _06355_, _06240_);
  nor (_06408_, _06406_, _06405_);
  nor (_06409_, _06408_, _06352_);
  and (_06410_, _06352_, word_in[11]);
  or (_06411_, _06410_, _06362_);
  or (_06412_, _06411_, _06409_);
  and (_06413_, _06412_, _06403_);
  or (_06414_, _06413_, _06350_);
  or (_06415_, _06372_, word_in[27]);
  and (_26821_[3], _06415_, _06414_);
  and (_06416_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and (_06417_, _02838_, _23983_);
  or (_27140_, _06417_, _06416_);
  or (_06418_, _06367_, word_in[20]);
  not (_06419_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_06420_, _06355_, _06419_);
  and (_06421_, _06355_, _06259_);
  nor (_06422_, _06421_, _06420_);
  nor (_06423_, _06422_, _06352_);
  and (_06424_, _06352_, word_in[12]);
  or (_06425_, _06424_, _06362_);
  or (_06426_, _06425_, _06423_);
  and (_06427_, _06426_, _06418_);
  or (_06428_, _06427_, _06350_);
  or (_06429_, _06372_, word_in[28]);
  and (_26821_[4], _06429_, _06428_);
  not (_06430_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_06431_, _06355_, _06430_);
  and (_06432_, _06355_, _06278_);
  nor (_06434_, _06432_, _06431_);
  nor (_06435_, _06434_, _06352_);
  and (_06437_, _06352_, word_in[13]);
  or (_06438_, _06437_, _06362_);
  or (_06439_, _06438_, _06435_);
  or (_06440_, _06367_, word_in[21]);
  and (_06442_, _06440_, _06439_);
  or (_06443_, _06442_, _06350_);
  or (_06444_, _06372_, word_in[29]);
  and (_26821_[5], _06444_, _06443_);
  and (_06445_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_06446_, _02775_, _24027_);
  or (_27142_, _06446_, _06445_);
  not (_06447_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_06448_, _06355_, _06447_);
  and (_06449_, _06355_, _06294_);
  nor (_06450_, _06449_, _06448_);
  nor (_06451_, _06450_, _06352_);
  and (_06452_, _06352_, word_in[14]);
  or (_06453_, _06452_, _06362_);
  or (_06455_, _06453_, _06451_);
  or (_06456_, _06367_, word_in[22]);
  and (_06457_, _06456_, _06455_);
  or (_06458_, _06457_, _06350_);
  or (_06459_, _06372_, word_in[30]);
  and (_26821_[6], _06459_, _06458_);
  nor (_06461_, _06355_, _05065_);
  and (_06462_, _06355_, _05407_);
  nor (_06463_, _06462_, _06461_);
  nor (_06464_, _06463_, _06352_);
  and (_06466_, _06352_, word_in[15]);
  or (_06467_, _06466_, _06362_);
  or (_06468_, _06467_, _06464_);
  or (_06469_, _06367_, word_in[23]);
  and (_06470_, _06469_, _06468_);
  and (_06471_, _06470_, _06372_);
  and (_06472_, _06350_, word_in[31]);
  or (_26821_[7], _06472_, _06471_);
  and (_06473_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  and (_06474_, _03169_, _24053_);
  or (_02042_, _06474_, _06473_);
  and (_06475_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and (_06476_, _03169_, _23920_);
  or (_02057_, _06476_, _06475_);
  and (_06478_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  and (_06479_, _03165_, _24027_);
  or (_02061_, _06479_, _06478_);
  and (_06482_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  and (_06484_, _03165_, _23715_);
  or (_02065_, _06484_, _06482_);
  and (_06485_, _05385_, _05123_);
  and (_06486_, _06485_, _05324_);
  and (_06487_, _05399_, _05151_);
  and (_06488_, _06487_, _05135_);
  not (_06489_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not (_06490_, _05402_);
  and (_06491_, _06179_, _06490_);
  and (_06492_, _06491_, _05816_);
  nor (_06493_, _06492_, _06489_);
  and (_06494_, _06492_, _06188_);
  nor (_06495_, _06494_, _06493_);
  nor (_06496_, _06495_, _06488_);
  and (_06497_, _05394_, _05120_);
  and (_06498_, _06497_, _05242_);
  and (_06499_, _06488_, word_in[8]);
  or (_06500_, _06499_, _06498_);
  or (_06501_, _06500_, _06496_);
  not (_06502_, _06498_);
  or (_06503_, _06502_, word_in[16]);
  and (_06504_, _06503_, _06501_);
  or (_06505_, _06504_, _06486_);
  not (_06506_, _06486_);
  or (_06507_, _06506_, word_in[24]);
  and (_26822_[0], _06507_, _06505_);
  not (_06508_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_06509_, _06492_, _06508_);
  and (_06510_, _06492_, _06212_);
  nor (_06511_, _06510_, _06509_);
  nor (_06512_, _06511_, _06488_);
  and (_06513_, _06488_, word_in[9]);
  or (_06514_, _06513_, _06498_);
  or (_06515_, _06514_, _06512_);
  or (_06516_, _06502_, word_in[17]);
  and (_06517_, _06516_, _06515_);
  or (_06518_, _06517_, _06486_);
  or (_06519_, _06506_, word_in[25]);
  and (_26822_[1], _06519_, _06518_);
  or (_06521_, _06502_, word_in[18]);
  not (_06522_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_06524_, _06492_, _06522_);
  and (_06525_, _06492_, _06227_);
  nor (_06527_, _06525_, _06524_);
  nor (_06529_, _06527_, _06488_);
  and (_06530_, _06488_, word_in[10]);
  or (_06531_, _06530_, _06498_);
  or (_06532_, _06531_, _06529_);
  and (_06533_, _06532_, _06521_);
  or (_06534_, _06533_, _06486_);
  or (_06536_, _06506_, word_in[26]);
  and (_26822_[2], _06536_, _06534_);
  not (_06539_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_06540_, _06492_, _06539_);
  and (_06541_, _06492_, _06240_);
  nor (_06542_, _06541_, _06540_);
  nor (_06543_, _06542_, _06488_);
  and (_06544_, _06488_, word_in[11]);
  or (_06545_, _06544_, _06498_);
  or (_06547_, _06545_, _06543_);
  or (_06548_, _06502_, word_in[19]);
  and (_06549_, _06548_, _06547_);
  or (_06551_, _06549_, _06486_);
  or (_06552_, _06506_, word_in[27]);
  and (_26822_[3], _06552_, _06551_);
  not (_06553_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_06554_, _06492_, _06553_);
  and (_06555_, _06492_, _06259_);
  nor (_06557_, _06555_, _06554_);
  nor (_06558_, _06557_, _06488_);
  and (_06560_, _06488_, word_in[12]);
  or (_06561_, _06560_, _06498_);
  or (_06562_, _06561_, _06558_);
  or (_06563_, _06502_, word_in[20]);
  and (_06566_, _06563_, _06562_);
  or (_06567_, _06566_, _06486_);
  or (_06568_, _06506_, word_in[28]);
  and (_26822_[4], _06568_, _06567_);
  not (_06569_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_06570_, _06492_, _06569_);
  and (_06571_, _06492_, _06278_);
  nor (_06572_, _06571_, _06570_);
  nor (_06573_, _06572_, _06488_);
  and (_06574_, _06488_, word_in[13]);
  or (_06575_, _06574_, _06498_);
  or (_06576_, _06575_, _06573_);
  or (_06577_, _06502_, word_in[21]);
  and (_06578_, _06577_, _06576_);
  or (_06579_, _06578_, _06486_);
  or (_06580_, _06506_, word_in[29]);
  and (_26822_[5], _06580_, _06579_);
  or (_06581_, _06502_, word_in[22]);
  not (_06582_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_06583_, _06492_, _06582_);
  and (_06584_, _06492_, _06294_);
  nor (_06585_, _06584_, _06583_);
  nor (_06586_, _06585_, _06488_);
  and (_06587_, _06488_, word_in[14]);
  or (_06588_, _06587_, _06498_);
  or (_06589_, _06588_, _06586_);
  and (_06590_, _06589_, _06581_);
  or (_06591_, _06590_, _06486_);
  or (_06592_, _06506_, word_in[30]);
  and (_26822_[6], _06592_, _06591_);
  and (_06593_, _04207_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and (_06594_, _25876_, _24648_);
  or (_06595_, _06054_, _25920_);
  or (_06596_, _06595_, _06594_);
  or (_06597_, _04935_, _26229_);
  or (_06598_, _06597_, _25879_);
  or (_06599_, _06598_, _06131_);
  or (_06600_, _06599_, _06596_);
  or (_06602_, _06081_, _24693_);
  or (_06603_, _06602_, _04947_);
  or (_06605_, _06603_, _06112_);
  or (_06606_, _06605_, _06600_);
  or (_06607_, _06606_, _06079_);
  and (_06608_, _06607_, _01886_);
  or (_26843_[0], _06608_, _06593_);
  nor (_06609_, _06492_, _05174_);
  and (_06610_, _06492_, _05407_);
  nor (_06611_, _06610_, _06609_);
  nor (_06612_, _06611_, _06488_);
  and (_06613_, _06488_, word_in[15]);
  or (_06614_, _06613_, _06498_);
  or (_06615_, _06614_, _06612_);
  or (_06616_, _06502_, word_in[23]);
  and (_06617_, _06616_, _06615_);
  or (_06618_, _06617_, _06486_);
  or (_06619_, _06506_, word_in[31]);
  and (_26822_[7], _06619_, _06618_);
  and (_06621_, _02717_, _24061_);
  not (_06623_, _06621_);
  and (_06625_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_06626_, _06621_, _23900_);
  or (_02095_, _06626_, _06625_);
  and (_06627_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_06628_, _06621_, _24053_);
  or (_02102_, _06628_, _06627_);
  and (_06629_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_06630_, _03161_, _23693_);
  or (_02108_, _06630_, _06629_);
  and (_06631_, _23930_, _23706_);
  and (_06632_, _06631_, _23983_);
  not (_06633_, _06631_);
  and (_06635_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or (_26924_, _06635_, _06632_);
  and (_06636_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and (_06637_, _03157_, _24053_);
  or (_02131_, _06637_, _06636_);
  and (_06639_, _05385_, _05527_);
  and (_06641_, _05400_, _05135_);
  not (_06642_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_06643_, _06182_, _05403_);
  nor (_06645_, _06643_, _06642_);
  and (_06646_, _06643_, _06188_);
  nor (_06648_, _06646_, _06645_);
  nor (_06649_, _06648_, _06641_);
  and (_06651_, _05395_, _05242_);
  and (_06653_, _06641_, word_in[8]);
  or (_06654_, _06653_, _06651_);
  or (_06655_, _06654_, _06649_);
  not (_06656_, _06651_);
  or (_06657_, _06656_, word_in[16]);
  and (_06658_, _06657_, _06655_);
  or (_06659_, _06658_, _06639_);
  not (_06661_, _06639_);
  or (_06663_, _06661_, word_in[24]);
  and (_26823_[0], _06663_, _06659_);
  not (_06664_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_06666_, _06643_, _06664_);
  and (_06667_, _06643_, _06212_);
  nor (_06669_, _06667_, _06666_);
  nor (_06670_, _06669_, _06641_);
  and (_06672_, _06641_, word_in[9]);
  or (_06674_, _06672_, _06651_);
  or (_06675_, _06674_, _06670_);
  or (_06676_, _06656_, word_in[17]);
  and (_06678_, _06676_, _06661_);
  and (_06679_, _06678_, _06675_);
  and (_06681_, _06639_, word_in[25]);
  or (_26823_[1], _06681_, _06679_);
  nand (_26833_[0], _04973_, _01886_);
  or (_06684_, _06656_, word_in[18]);
  not (_06686_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_06688_, _06643_, _06686_);
  and (_06689_, _06643_, _06227_);
  nor (_06690_, _06689_, _06688_);
  nor (_06691_, _06690_, _06641_);
  and (_06692_, _06641_, word_in[10]);
  or (_06694_, _06692_, _06651_);
  or (_06696_, _06694_, _06691_);
  and (_06698_, _06696_, _06684_);
  and (_06699_, _06698_, _06661_);
  and (_06700_, _06639_, word_in[26]);
  or (_26823_[2], _06700_, _06699_);
  or (_06702_, _06656_, word_in[19]);
  not (_06703_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_06704_, _06643_, _06703_);
  and (_06705_, _06643_, _06240_);
  nor (_06706_, _06705_, _06704_);
  nor (_06707_, _06706_, _06641_);
  and (_06709_, _06641_, word_in[11]);
  or (_06710_, _06709_, _06651_);
  or (_06711_, _06710_, _06707_);
  and (_06712_, _06711_, _06702_);
  or (_06713_, _06712_, _06639_);
  or (_06714_, _06661_, word_in[27]);
  and (_26823_[3], _06714_, _06713_);
  or (_06715_, _06656_, word_in[20]);
  not (_06716_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_06717_, _06643_, _06716_);
  and (_06718_, _06643_, _06259_);
  nor (_06719_, _06718_, _06717_);
  nor (_06720_, _06719_, _06641_);
  and (_06721_, _06641_, word_in[12]);
  or (_06722_, _06721_, _06651_);
  or (_06723_, _06722_, _06720_);
  and (_06724_, _06723_, _06715_);
  or (_06725_, _06724_, _06639_);
  or (_06726_, _06661_, word_in[28]);
  and (_26823_[4], _06726_, _06725_);
  and (_06727_, _06639_, word_in[29]);
  not (_06728_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_06730_, _06643_, _06728_);
  and (_06732_, _06643_, _06278_);
  nor (_06733_, _06732_, _06730_);
  nor (_06735_, _06733_, _06641_);
  and (_06736_, _06641_, word_in[13]);
  or (_06737_, _06736_, _06651_);
  or (_06738_, _06737_, _06735_);
  or (_06739_, _06656_, word_in[21]);
  and (_06740_, _06739_, _06661_);
  and (_06741_, _06740_, _06738_);
  or (_26823_[5], _06741_, _06727_);
  or (_06743_, _06656_, word_in[22]);
  not (_06745_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_06747_, _06643_, _06745_);
  and (_06748_, _06643_, _06294_);
  nor (_06750_, _06748_, _06747_);
  nor (_06751_, _06750_, _06641_);
  and (_06752_, _06641_, word_in[14]);
  or (_06753_, _06752_, _06651_);
  or (_06754_, _06753_, _06751_);
  and (_06755_, _06754_, _06743_);
  or (_06756_, _06755_, _06639_);
  or (_06758_, _06661_, word_in[30]);
  and (_26823_[6], _06758_, _06756_);
  or (_06760_, _06656_, word_in[23]);
  nor (_06762_, _06643_, _05083_);
  and (_06764_, _06643_, _05407_);
  nor (_06765_, _06764_, _06762_);
  nor (_06767_, _06765_, _06641_);
  and (_06768_, _06641_, word_in[15]);
  or (_06769_, _06768_, _06651_);
  or (_06771_, _06769_, _06767_);
  and (_06772_, _06771_, _06760_);
  or (_06773_, _06772_, _06639_);
  or (_06775_, _06661_, word_in[31]);
  and (_26823_[7], _06775_, _06773_);
  and (_06776_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_06777_, _02722_, _23751_);
  or (_02169_, _06777_, _06776_);
  and (_06778_, _01932_, _23715_);
  and (_06779_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_27031_, _06779_, _06778_);
  and (_06782_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_06783_, _02722_, _24027_);
  or (_02180_, _06783_, _06782_);
  and (_06785_, _05385_, _05310_);
  and (_06786_, _06785_, _05316_);
  and (_06788_, _06786_, _05151_);
  and (_06789_, _05394_, _05479_);
  not (_06791_, _06789_);
  or (_06792_, _06791_, word_in[16]);
  and (_06794_, _05399_, _05496_);
  not (_06795_, _06794_);
  not (_06797_, word_in[0]);
  and (_06798_, _05404_, _05130_);
  and (_06799_, _06798_, _06180_);
  nand (_06800_, _06799_, _06797_);
  or (_06801_, _06799_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_06802_, _06801_, _06800_);
  and (_06803_, _06802_, _06795_);
  and (_06804_, _06794_, word_in[8]);
  or (_06805_, _06804_, _06789_);
  or (_06807_, _06805_, _06803_);
  and (_06808_, _06807_, _06792_);
  or (_06809_, _06808_, _06788_);
  and (_06810_, _05385_, word_in[24]);
  not (_06811_, _06788_);
  or (_06812_, _06811_, _06810_);
  and (_26824_[0], _06812_, _06809_);
  or (_06813_, _06791_, word_in[17]);
  or (_06814_, _06799_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  not (_06815_, word_in[1]);
  nand (_06816_, _06799_, _06815_);
  and (_06817_, _06816_, _06814_);
  or (_06818_, _06817_, _06794_);
  or (_06819_, _06795_, word_in[9]);
  and (_06820_, _06819_, _06818_);
  or (_06821_, _06820_, _06789_);
  and (_06822_, _06821_, _06813_);
  or (_06823_, _06822_, _06788_);
  or (_06824_, _06811_, _06207_);
  and (_26824_[1], _06824_, _06823_);
  or (_06825_, _06791_, word_in[18]);
  not (_06827_, word_in[2]);
  nand (_06828_, _06799_, _06827_);
  or (_06830_, _06799_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_06831_, _06830_, _06828_);
  or (_06832_, _06831_, _06794_);
  or (_06833_, _06795_, word_in[10]);
  and (_06834_, _06833_, _06832_);
  or (_06836_, _06834_, _06789_);
  and (_06838_, _06836_, _06825_);
  or (_06840_, _06838_, _06788_);
  and (_06842_, _05385_, word_in[26]);
  or (_06844_, _06811_, _06842_);
  and (_26824_[2], _06844_, _06840_);
  not (_06845_, word_in[3]);
  nand (_06846_, _06799_, _06845_);
  or (_06847_, _06799_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_06849_, _06847_, _06846_);
  or (_06850_, _06849_, _06794_);
  or (_06851_, _06795_, word_in[11]);
  and (_06853_, _06851_, _06850_);
  or (_06855_, _06853_, _06789_);
  nor (_06856_, _06791_, _06247_);
  nor (_06858_, _06856_, _06788_);
  and (_06860_, _06858_, _06855_);
  and (_06861_, _05385_, word_in[27]);
  and (_06862_, _06788_, _06861_);
  or (_26813_, _06862_, _06860_);
  or (_06863_, _06791_, word_in[20]);
  not (_06864_, word_in[4]);
  nand (_06865_, _06799_, _06864_);
  or (_06867_, _06799_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_06868_, _06867_, _06865_);
  or (_06869_, _06868_, _06794_);
  or (_06870_, _06795_, word_in[12]);
  and (_06871_, _06870_, _06869_);
  or (_06872_, _06871_, _06789_);
  and (_06873_, _06872_, _06863_);
  or (_06874_, _06873_, _06788_);
  and (_06876_, _05385_, word_in[28]);
  or (_06878_, _06811_, _06876_);
  and (_26824_[4], _06878_, _06874_);
  or (_06880_, _06791_, word_in[21]);
  not (_06881_, word_in[5]);
  nand (_06882_, _06799_, _06881_);
  or (_06883_, _06799_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_06885_, _06883_, _06882_);
  or (_06886_, _06885_, _06794_);
  or (_06889_, _06795_, word_in[13]);
  and (_06891_, _06889_, _06886_);
  or (_06892_, _06891_, _06789_);
  and (_06894_, _06892_, _06880_);
  or (_06896_, _06894_, _06788_);
  or (_06897_, _06811_, _06273_);
  and (_26824_[5], _06897_, _06896_);
  not (_06900_, word_in[6]);
  nand (_06901_, _06799_, _06900_);
  or (_06903_, _06799_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_06904_, _06903_, _06901_);
  or (_06905_, _06904_, _06794_);
  or (_06906_, _06795_, word_in[14]);
  and (_06907_, _06906_, _06905_);
  or (_06908_, _06907_, _06789_);
  nor (_06909_, _06791_, word_in[22]);
  nor (_06910_, _06909_, _06788_);
  and (_06911_, _06910_, _06908_);
  and (_06912_, _05385_, word_in[30]);
  and (_06913_, _06788_, _06912_);
  or (_26824_[6], _06913_, _06911_);
  nor (_06915_, _06799_, _05209_);
  and (_06916_, _06799_, _05407_);
  or (_06917_, _06916_, _06915_);
  or (_06918_, _06917_, _06794_);
  or (_06919_, _06795_, word_in[15]);
  and (_06920_, _06919_, _06918_);
  or (_06921_, _06920_, _06789_);
  or (_06922_, _06791_, word_in[23]);
  and (_06923_, _06922_, _06921_);
  or (_06924_, _06923_, _06788_);
  or (_06925_, _06811_, _05387_);
  and (_26824_[7], _06925_, _06924_);
  and (_06926_, _06361_, _05893_);
  not (_06927_, _06926_);
  and (_06928_, _06351_, _05202_);
  not (_06929_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_06930_, _06798_, _06354_);
  nor (_06931_, _06930_, _06929_);
  and (_06932_, _06930_, _06188_);
  nor (_06933_, _06932_, _06931_);
  nor (_06934_, _06933_, _06928_);
  and (_06935_, _06928_, word_in[8]);
  or (_06936_, _06935_, _06934_);
  and (_06937_, _06936_, _06927_);
  and (_06938_, _06786_, _05161_);
  and (_06939_, _06926_, word_in[16]);
  or (_06940_, _06939_, _06938_);
  or (_06941_, _06940_, _06937_);
  not (_06942_, _06938_);
  or (_06943_, _06942_, word_in[24]);
  and (_26825_[0], _06943_, _06941_);
  not (_06944_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_06945_, _06930_, _06944_);
  and (_06946_, _06930_, _06212_);
  or (_06947_, _06946_, _06945_);
  or (_06949_, _06947_, _06928_);
  not (_06950_, _06928_);
  or (_06951_, _06950_, word_in[9]);
  and (_06952_, _06951_, _06949_);
  or (_06953_, _06952_, _06926_);
  or (_06954_, _06927_, word_in[17]);
  and (_06955_, _06954_, _06953_);
  or (_06956_, _06955_, _06938_);
  or (_06957_, _06942_, word_in[25]);
  and (_26825_[1], _06957_, _06956_);
  not (_06958_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_06959_, _06930_, _06958_);
  and (_06960_, _06930_, _06227_);
  nor (_06961_, _06960_, _06959_);
  nor (_06962_, _06961_, _06928_);
  and (_06963_, _06928_, word_in[10]);
  or (_06964_, _06963_, _06962_);
  and (_06966_, _06964_, _06927_);
  and (_06967_, _06926_, word_in[18]);
  or (_06968_, _06967_, _06938_);
  or (_06969_, _06968_, _06966_);
  or (_06970_, _06942_, word_in[26]);
  and (_26825_[2], _06970_, _06969_);
  not (_06972_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_06974_, _06930_, _06972_);
  and (_06975_, _06930_, _06240_);
  or (_06976_, _06975_, _06974_);
  or (_06977_, _06976_, _06928_);
  or (_06979_, _06950_, word_in[11]);
  and (_06980_, _06979_, _06977_);
  or (_06981_, _06980_, _06926_);
  or (_06982_, _06927_, word_in[19]);
  and (_06983_, _06982_, _06981_);
  or (_06984_, _06983_, _06938_);
  or (_06985_, _06942_, word_in[27]);
  and (_26825_[3], _06985_, _06984_);
  not (_06987_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_06988_, _06930_, _06987_);
  and (_06989_, _06930_, _06259_);
  nor (_06990_, _06989_, _06988_);
  nor (_06991_, _06990_, _06928_);
  and (_06993_, _06928_, word_in[12]);
  or (_06994_, _06993_, _06991_);
  and (_06995_, _06994_, _06927_);
  and (_06996_, _06926_, word_in[20]);
  or (_06997_, _06996_, _06938_);
  or (_06998_, _06997_, _06995_);
  or (_06999_, _06942_, word_in[28]);
  and (_26825_[4], _06999_, _06998_);
  not (_07000_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_07001_, _06930_, _07000_);
  and (_07002_, _06930_, _06278_);
  or (_07003_, _07002_, _07001_);
  or (_07004_, _07003_, _06928_);
  or (_07005_, _06950_, word_in[13]);
  and (_07006_, _07005_, _07004_);
  or (_07007_, _07006_, _06926_);
  or (_07008_, _06927_, word_in[21]);
  and (_07009_, _07008_, _07007_);
  and (_07010_, _07009_, _06942_);
  and (_07011_, _06938_, word_in[29]);
  or (_26825_[5], _07011_, _07010_);
  not (_07013_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_07014_, _06930_, _07013_);
  and (_07015_, _06930_, _06294_);
  or (_07016_, _07015_, _07014_);
  or (_07018_, _07016_, _06928_);
  or (_07019_, _06950_, word_in[14]);
  and (_07020_, _07019_, _07018_);
  or (_07021_, _07020_, _06926_);
  or (_07022_, _06927_, word_in[22]);
  and (_07024_, _07022_, _07021_);
  or (_07025_, _07024_, _06938_);
  or (_07026_, _06942_, word_in[30]);
  and (_26825_[6], _07026_, _07025_);
  nor (_07027_, _06930_, _05077_);
  and (_07028_, _06930_, _05407_);
  nor (_07029_, _07028_, _07027_);
  nor (_07030_, _07029_, _06928_);
  and (_07032_, _06928_, word_in[15]);
  or (_07033_, _07032_, _07030_);
  and (_07034_, _07033_, _06927_);
  and (_07036_, _06926_, word_in[23]);
  or (_07037_, _07036_, _06938_);
  or (_07038_, _07037_, _07034_);
  or (_07040_, _06942_, word_in[31]);
  and (_26825_[7], _07040_, _07038_);
  and (_07041_, _06786_, _05123_);
  and (_07042_, _06497_, _05893_);
  not (_07043_, _07042_);
  or (_07044_, _07043_, word_in[16]);
  and (_07046_, _06487_, _05202_);
  and (_07047_, _06798_, _06491_);
  nand (_07048_, _07047_, _06797_);
  or (_07049_, _07047_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand (_07050_, _07049_, _07048_);
  nor (_07051_, _07050_, _07046_);
  and (_07052_, _07046_, word_in[8]);
  or (_07053_, _07052_, _07042_);
  or (_07054_, _07053_, _07051_);
  and (_07055_, _07054_, _07044_);
  or (_07056_, _07055_, _07041_);
  not (_07057_, _07041_);
  or (_07058_, _07057_, word_in[24]);
  and (_26826_[0], _07058_, _07056_);
  or (_07059_, _07047_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nand (_07060_, _07047_, _06815_);
  and (_07062_, _07060_, _07059_);
  or (_07064_, _07062_, _07046_);
  not (_07066_, _07046_);
  or (_07067_, _07066_, word_in[9]);
  and (_07068_, _07067_, _07064_);
  or (_07069_, _07068_, _07042_);
  nor (_07071_, _07043_, word_in[17]);
  nor (_07072_, _07071_, _07041_);
  and (_07073_, _07072_, _07069_);
  and (_07075_, _07041_, word_in[25]);
  or (_26826_[1], _07075_, _07073_);
  or (_07076_, _07047_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand (_07077_, _07047_, _06827_);
  and (_07078_, _07077_, _07076_);
  or (_07079_, _07078_, _07046_);
  or (_07080_, _07066_, word_in[10]);
  and (_07081_, _07080_, _07079_);
  or (_07082_, _07081_, _07042_);
  or (_07083_, _07043_, word_in[18]);
  and (_07084_, _07083_, _07082_);
  or (_07085_, _07084_, _07041_);
  or (_07086_, _07057_, word_in[26]);
  and (_26826_[2], _07086_, _07085_);
  and (_07087_, _23924_, _23719_);
  and (_07088_, _07087_, _23693_);
  not (_07089_, _07087_);
  and (_07090_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_02294_, _07090_, _07088_);
  or (_07091_, _07047_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nand (_07092_, _07047_, _06845_);
  and (_07093_, _07092_, _07091_);
  or (_07094_, _07093_, _07046_);
  or (_07095_, _07066_, word_in[11]);
  and (_07096_, _07095_, _07094_);
  or (_07097_, _07096_, _07042_);
  or (_07098_, _07043_, word_in[19]);
  and (_07100_, _07098_, _07097_);
  or (_07101_, _07100_, _07041_);
  or (_07102_, _07057_, word_in[27]);
  and (_26826_[3], _07102_, _07101_);
  or (_07103_, _07047_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nand (_07104_, _07047_, _06864_);
  and (_07105_, _07104_, _07103_);
  or (_07106_, _07105_, _07046_);
  or (_07107_, _07066_, word_in[12]);
  and (_07108_, _07107_, _07106_);
  or (_07109_, _07108_, _07042_);
  nor (_07110_, _07043_, word_in[20]);
  nor (_07111_, _07110_, _07041_);
  and (_07112_, _07111_, _07109_);
  and (_07113_, _07041_, word_in[28]);
  or (_26826_[4], _07113_, _07112_);
  and (_07114_, _07087_, _23900_);
  and (_07115_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_02299_, _07115_, _07114_);
  or (_07116_, _07047_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nand (_07117_, _07047_, _06881_);
  and (_07118_, _07117_, _07116_);
  or (_07119_, _07118_, _07046_);
  or (_07120_, _07066_, word_in[13]);
  and (_07121_, _07120_, _07119_);
  or (_07122_, _07121_, _07042_);
  or (_07123_, _07043_, word_in[21]);
  and (_07124_, _07123_, _07122_);
  or (_07125_, _07124_, _07041_);
  or (_07126_, _07057_, word_in[29]);
  and (_26826_[5], _07126_, _07125_);
  or (_07127_, _07047_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nand (_07128_, _07047_, _06900_);
  and (_07129_, _07128_, _07127_);
  or (_07130_, _07129_, _07046_);
  or (_07131_, _07066_, word_in[14]);
  and (_07132_, _07131_, _07130_);
  or (_07133_, _07132_, _07042_);
  or (_07134_, _07043_, word_in[22]);
  and (_07135_, _07134_, _07133_);
  or (_07136_, _07135_, _07041_);
  or (_07137_, _07057_, word_in[30]);
  and (_26826_[6], _07137_, _07136_);
  nor (_07138_, _07047_, _05204_);
  and (_07139_, _07047_, _05407_);
  or (_07140_, _07139_, _07138_);
  or (_07141_, _07140_, _07046_);
  or (_07142_, _07066_, word_in[15]);
  and (_07144_, _07142_, _07141_);
  or (_07145_, _07144_, _07042_);
  or (_07146_, _07043_, word_in[23]);
  and (_07147_, _07146_, _07145_);
  or (_07148_, _07147_, _07041_);
  or (_07149_, _07057_, word_in[31]);
  and (_26826_[7], _07149_, _07148_);
  and (_07151_, _05883_, _23983_);
  and (_07152_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_02342_, _07152_, _07151_);
  and (_07155_, _05893_, _05395_);
  and (_07156_, _05400_, _05202_);
  not (_07157_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_07158_, _06798_, _05403_);
  nor (_07160_, _07158_, _07157_);
  and (_07162_, _07158_, _06188_);
  or (_07164_, _07162_, _07160_);
  or (_07166_, _07164_, _07156_);
  not (_07167_, _07156_);
  or (_07168_, _07167_, word_in[8]);
  and (_07169_, _07168_, _07166_);
  or (_07170_, _07169_, _07155_);
  and (_07171_, _05385_, _05517_);
  not (_07172_, _07171_);
  and (_07174_, _05394_, word_in[16]);
  not (_07175_, _07155_);
  or (_07177_, _07175_, _07174_);
  and (_07179_, _07177_, _07172_);
  and (_07181_, _07179_, _07170_);
  and (_07183_, _07171_, word_in[24]);
  or (_26827_[0], _07183_, _07181_);
  and (_07184_, _07171_, _06207_);
  not (_07185_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_07187_, _07158_, _07185_);
  and (_07188_, _07158_, _06212_);
  nor (_07189_, _07188_, _07187_);
  nor (_07190_, _07189_, _07156_);
  and (_07191_, _07156_, word_in[9]);
  or (_07192_, _07191_, _07190_);
  and (_07193_, _07192_, _07175_);
  and (_07194_, _05394_, word_in[17]);
  and (_07195_, _07155_, _07194_);
  or (_07196_, _07195_, _07193_);
  and (_07197_, _07196_, _07172_);
  or (_26827_[1], _07197_, _07184_);
  and (_07198_, _05394_, word_in[18]);
  and (_07199_, _07155_, _07198_);
  not (_07200_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_07201_, _07158_, _07200_);
  and (_07202_, _07158_, _06227_);
  nor (_07203_, _07202_, _07201_);
  nor (_07205_, _07203_, _07156_);
  and (_07207_, _07156_, word_in[10]);
  or (_07208_, _07207_, _07205_);
  and (_07210_, _07208_, _07175_);
  or (_07212_, _07210_, _07199_);
  and (_07213_, _07212_, _07172_);
  and (_07215_, _07171_, word_in[26]);
  or (_26827_[2], _07215_, _07213_);
  and (_07216_, _07171_, _06861_);
  not (_07218_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_07219_, _07158_, _07218_);
  and (_07221_, _07158_, _06240_);
  nor (_07222_, _07221_, _07219_);
  nor (_07223_, _07222_, _07156_);
  and (_07225_, _07156_, word_in[11]);
  or (_07226_, _07225_, _07223_);
  and (_07228_, _07226_, _07175_);
  and (_07230_, _07155_, _06247_);
  or (_07232_, _07230_, _07228_);
  and (_07234_, _07232_, _07172_);
  or (_26827_[3], _07234_, _07216_);
  and (_07235_, _05394_, word_in[20]);
  and (_07237_, _07155_, _07235_);
  not (_07238_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_07239_, _07158_, _07238_);
  and (_07240_, _07158_, _06259_);
  nor (_07241_, _07240_, _07239_);
  nor (_07242_, _07241_, _07156_);
  and (_07244_, _07156_, word_in[12]);
  or (_07245_, _07244_, _07242_);
  and (_07247_, _07245_, _07175_);
  or (_07249_, _07247_, _07237_);
  and (_07251_, _07249_, _07172_);
  and (_07253_, _07171_, word_in[28]);
  or (_26827_[4], _07253_, _07251_);
  and (_07254_, _07171_, _06273_);
  and (_07255_, _07158_, _06278_);
  not (_07257_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_07258_, _07158_, _07257_);
  nor (_07260_, _07258_, _07255_);
  nor (_07262_, _07260_, _07156_);
  and (_07263_, _07156_, word_in[13]);
  or (_07265_, _07263_, _07262_);
  or (_07267_, _07265_, _07155_);
  and (_07268_, _05394_, word_in[21]);
  or (_07270_, _07175_, _07268_);
  and (_07272_, _07270_, _07172_);
  and (_07274_, _07272_, _07267_);
  or (_26827_[5], _07274_, _07254_);
  and (_07276_, _07171_, _06912_);
  and (_07278_, _07158_, _06294_);
  not (_07279_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_07280_, _07158_, _07279_);
  nor (_07281_, _07280_, _07278_);
  nor (_07283_, _07281_, _07156_);
  and (_07284_, _07156_, word_in[14]);
  or (_07285_, _07284_, _07283_);
  and (_07286_, _07285_, _07175_);
  and (_07287_, _05394_, word_in[22]);
  and (_07289_, _07155_, _07287_);
  or (_07290_, _07289_, _07286_);
  and (_07291_, _07290_, _07172_);
  or (_26827_[6], _07291_, _07276_);
  or (_07293_, _07175_, _05415_);
  nor (_07294_, _07158_, _05072_);
  and (_07296_, _07158_, _05407_);
  or (_07297_, _07296_, _07294_);
  or (_07298_, _07297_, _07156_);
  or (_07300_, _07167_, word_in[15]);
  and (_07301_, _07300_, _07298_);
  or (_07302_, _07301_, _07155_);
  and (_07303_, _07302_, _07293_);
  or (_07304_, _07303_, _07171_);
  or (_07305_, _07172_, word_in[31]);
  and (_26827_[7], _07305_, _07304_);
  and (_07307_, _07087_, _23715_);
  and (_07309_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_02374_, _07309_, _07307_);
  not (_07311_, _24192_);
  or (_07312_, _07311_, _23744_);
  and (_07313_, _24984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_07314_, _07313_, _25011_);
  and (_07315_, _07314_, _25000_);
  or (_07316_, _07315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_07317_, _07315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_07318_, _07317_, _25003_);
  and (_07319_, _07318_, _07316_);
  and (_07320_, _24193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_07321_, _07320_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_07322_, _24200_, _24193_);
  not (_07323_, _07322_);
  and (_07324_, _07323_, _24196_);
  and (_07325_, _07324_, _07321_);
  and (_07326_, _07313_, _25007_);
  nor (_07327_, _07326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_07328_, _07326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_07329_, _07328_, _07327_);
  and (_07330_, _07329_, _24975_);
  or (_07331_, _07330_, _07325_);
  or (_07333_, _07331_, _07319_);
  or (_07334_, _07333_, _24192_);
  and (_07336_, _07334_, _24188_);
  and (_07338_, _07336_, _07312_);
  and (_07339_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_07340_, _07339_, _07338_);
  and (_02389_, _07340_, _22773_);
  and (_07342_, _05883_, _24027_);
  and (_07343_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_02398_, _07343_, _07342_);
  and (_07346_, _05385_, _05317_);
  and (_07347_, _07346_, _05151_);
  and (_07349_, _05394_, _05592_);
  not (_07351_, _07349_);
  or (_07352_, _07351_, word_in[16]);
  and (_07354_, _05399_, _05131_);
  and (_07355_, _05040_, _04991_);
  and (_07356_, _05404_, _07355_);
  and (_07357_, _07356_, _06180_);
  or (_07358_, _07357_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nand (_07359_, _07357_, _06797_);
  and (_07361_, _07359_, _07358_);
  or (_07362_, _07361_, _07354_);
  not (_07364_, _07354_);
  or (_07365_, _07364_, word_in[8]);
  and (_07366_, _07365_, _07362_);
  or (_07367_, _07366_, _07349_);
  and (_07369_, _07367_, _07352_);
  or (_07370_, _07369_, _07347_);
  not (_07372_, _07347_);
  or (_07373_, _07372_, word_in[24]);
  and (_26828_[0], _07373_, _07370_);
  nand (_07376_, _07357_, _06815_);
  or (_07377_, _07357_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_07379_, _07377_, _07376_);
  or (_07381_, _07379_, _07354_);
  or (_07382_, _07364_, word_in[9]);
  and (_07383_, _07382_, _07381_);
  or (_07384_, _07383_, _07349_);
  nor (_07386_, _07351_, word_in[17]);
  nor (_07388_, _07386_, _07347_);
  and (_07389_, _07388_, _07384_);
  and (_07390_, _07347_, word_in[25]);
  or (_26828_[1], _07390_, _07389_);
  nand (_07391_, _07357_, _06827_);
  or (_07392_, _07357_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_07393_, _07392_, _07391_);
  or (_07394_, _07393_, _07354_);
  or (_07396_, _07364_, word_in[10]);
  and (_07397_, _07396_, _07394_);
  or (_07398_, _07397_, _07349_);
  nor (_07399_, _07351_, word_in[18]);
  nor (_07400_, _07399_, _07347_);
  and (_07401_, _07400_, _07398_);
  and (_07402_, _07347_, word_in[26]);
  or (_26828_[2], _07402_, _07401_);
  nand (_07404_, _07357_, _06845_);
  or (_07406_, _07357_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_07408_, _07406_, _07404_);
  or (_07410_, _07408_, _07354_);
  or (_07411_, _07364_, word_in[11]);
  and (_07413_, _07411_, _07410_);
  or (_07415_, _07413_, _07349_);
  nor (_07416_, _07351_, word_in[19]);
  nor (_07418_, _07416_, _07347_);
  and (_07419_, _07418_, _07415_);
  and (_07421_, _07347_, word_in[27]);
  or (_26828_[3], _07421_, _07419_);
  nand (_07422_, _07357_, _06864_);
  or (_07423_, _07357_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_07424_, _07423_, _07422_);
  or (_07425_, _07424_, _07354_);
  or (_07426_, _07364_, word_in[12]);
  and (_07427_, _07426_, _07425_);
  or (_07428_, _07427_, _07349_);
  nor (_07429_, _07351_, word_in[20]);
  nor (_07430_, _07429_, _07347_);
  and (_07431_, _07430_, _07428_);
  and (_07432_, _07347_, word_in[28]);
  or (_26828_[4], _07432_, _07431_);
  nand (_07433_, _07357_, _06881_);
  or (_07434_, _07357_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_07435_, _07434_, _07433_);
  or (_07436_, _07435_, _07354_);
  or (_07437_, _07364_, word_in[13]);
  and (_07438_, _07437_, _07436_);
  or (_07440_, _07438_, _07349_);
  nor (_07442_, _07351_, word_in[21]);
  nor (_07443_, _07442_, _07347_);
  and (_07444_, _07443_, _07440_);
  and (_07445_, _07347_, word_in[29]);
  or (_26828_[5], _07445_, _07444_);
  nand (_07447_, _07357_, _06900_);
  or (_07449_, _07357_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_07451_, _07449_, _07447_);
  or (_07453_, _07451_, _07354_);
  or (_07455_, _07364_, word_in[14]);
  and (_07456_, _07455_, _07453_);
  or (_07457_, _07456_, _07349_);
  nor (_07459_, _07351_, word_in[22]);
  nor (_07461_, _07459_, _07347_);
  and (_07463_, _07461_, _07457_);
  and (_07465_, _07347_, word_in[30]);
  or (_26828_[6], _07465_, _07463_);
  nor (_07467_, _07357_, _05193_);
  and (_07469_, _07357_, _05407_);
  or (_07471_, _07469_, _07467_);
  or (_07472_, _07471_, _07354_);
  or (_07474_, _07364_, word_in[15]);
  and (_07476_, _07474_, _07472_);
  or (_07478_, _07476_, _07349_);
  nor (_07479_, _07351_, word_in[23]);
  nor (_07481_, _07479_, _07347_);
  and (_07482_, _07481_, _07478_);
  and (_07483_, _07347_, word_in[31]);
  or (_26828_[7], _07483_, _07482_);
  and (_07484_, _23891_, _23700_);
  and (_07485_, _07484_, _23983_);
  not (_07487_, _07484_);
  and (_07488_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_02433_, _07488_, _07485_);
  and (_07489_, _01701_, _23920_);
  and (_07490_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or (_02442_, _07490_, _07489_);
  and (_07491_, _07484_, _24027_);
  and (_07492_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_02449_, _07492_, _07491_);
  and (_07494_, _07484_, _23920_);
  and (_07495_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_02459_, _07495_, _07494_);
  and (_07496_, _07346_, _05161_);
  and (_07497_, _06351_, _05133_);
  not (_07498_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_07500_, _07356_, _06354_);
  nor (_07501_, _07500_, _07498_);
  and (_07502_, _07500_, _06188_);
  nor (_07504_, _07502_, _07501_);
  nor (_07505_, _07504_, _07497_);
  and (_07506_, _06361_, _05246_);
  and (_07507_, _07497_, word_in[8]);
  or (_07509_, _07507_, _07506_);
  or (_07511_, _07509_, _07505_);
  not (_07512_, _07506_);
  or (_07513_, _07512_, _07174_);
  and (_07515_, _07513_, _07511_);
  or (_07516_, _07515_, _07496_);
  not (_07517_, _07496_);
  or (_07518_, _07517_, word_in[24]);
  and (_26829_[0], _07518_, _07516_);
  or (_07519_, _07512_, _07194_);
  not (_07520_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_07521_, _07500_, _07520_);
  and (_07522_, _07500_, _06212_);
  nor (_07523_, _07522_, _07521_);
  nor (_07524_, _07523_, _07497_);
  and (_07525_, _07497_, word_in[9]);
  or (_07526_, _07525_, _07506_);
  or (_07527_, _07526_, _07524_);
  and (_07528_, _07527_, _07519_);
  or (_07529_, _07528_, _07496_);
  or (_07530_, _07517_, word_in[25]);
  and (_26829_[1], _07530_, _07529_);
  not (_07531_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_07532_, _07500_, _07531_);
  and (_07534_, _07500_, _06227_);
  nor (_07536_, _07534_, _07532_);
  nor (_07537_, _07536_, _07497_);
  and (_07538_, _07497_, word_in[10]);
  or (_07539_, _07538_, _07506_);
  or (_07541_, _07539_, _07537_);
  or (_07542_, _07512_, _07198_);
  and (_07543_, _07542_, _07541_);
  or (_07545_, _07543_, _07496_);
  or (_07547_, _07517_, word_in[26]);
  and (_26829_[2], _07547_, _07545_);
  or (_07548_, _07512_, _06247_);
  not (_07549_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_07550_, _07500_, _07549_);
  and (_07551_, _07500_, _06240_);
  nor (_07552_, _07551_, _07550_);
  nor (_07553_, _07552_, _07497_);
  and (_07554_, _07497_, word_in[11]);
  or (_07555_, _07554_, _07506_);
  or (_07556_, _07555_, _07553_);
  and (_07557_, _07556_, _07548_);
  or (_07558_, _07557_, _07496_);
  or (_07560_, _07517_, word_in[27]);
  and (_26829_[3], _07560_, _07558_);
  not (_07561_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_07563_, _07500_, _07561_);
  and (_07564_, _07500_, _06259_);
  nor (_07566_, _07564_, _07563_);
  nor (_07567_, _07566_, _07497_);
  and (_07568_, _07497_, word_in[12]);
  or (_07569_, _07568_, _07506_);
  or (_07571_, _07569_, _07567_);
  or (_07573_, _07512_, _07235_);
  and (_07574_, _07573_, _07571_);
  or (_07576_, _07574_, _07496_);
  or (_07578_, _07517_, word_in[28]);
  and (_26829_[4], _07578_, _07576_);
  or (_07580_, _07512_, _07268_);
  not (_07581_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_07582_, _07500_, _07581_);
  and (_07583_, _07500_, _06278_);
  nor (_07584_, _07583_, _07582_);
  nor (_07585_, _07584_, _07497_);
  and (_07587_, _07497_, word_in[13]);
  or (_07588_, _07587_, _07506_);
  or (_07589_, _07588_, _07585_);
  and (_07590_, _07589_, _07580_);
  or (_07592_, _07590_, _07496_);
  or (_07593_, _07517_, word_in[29]);
  and (_26829_[5], _07593_, _07592_);
  not (_07597_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_07598_, _07500_, _07597_);
  and (_07599_, _07500_, _06294_);
  nor (_07600_, _07599_, _07598_);
  nor (_07601_, _07600_, _07497_);
  and (_07602_, _07497_, word_in[14]);
  or (_07604_, _07602_, _07506_);
  or (_07605_, _07604_, _07601_);
  or (_07607_, _07512_, _07287_);
  and (_07609_, _07607_, _07605_);
  or (_07610_, _07609_, _07496_);
  or (_07612_, _07517_, word_in[30]);
  and (_26829_[6], _07612_, _07610_);
  nor (_07614_, _07500_, _05092_);
  and (_07615_, _07500_, _05407_);
  nor (_07616_, _07615_, _07614_);
  nor (_07617_, _07616_, _07497_);
  and (_07618_, _07497_, word_in[15]);
  or (_07619_, _07618_, _07506_);
  or (_07620_, _07619_, _07617_);
  or (_07621_, _07512_, _05415_);
  and (_07622_, _07621_, _07620_);
  or (_07623_, _07622_, _07496_);
  or (_07624_, _07517_, word_in[31]);
  and (_26829_[7], _07624_, _07623_);
  and (_07625_, _07346_, _05123_);
  and (_07626_, _06497_, _05246_);
  not (_07627_, _07626_);
  or (_07628_, _07627_, _07174_);
  and (_07629_, _06487_, _05133_);
  not (_07630_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_07631_, _07356_, _06491_);
  nor (_07632_, _07631_, _07630_);
  and (_07633_, _07631_, _06188_);
  nor (_07634_, _07633_, _07632_);
  nor (_07635_, _07634_, _07629_);
  and (_07636_, _07629_, word_in[8]);
  or (_07637_, _07636_, _07626_);
  or (_07638_, _07637_, _07635_);
  and (_07639_, _07638_, _07628_);
  or (_07640_, _07639_, _07625_);
  not (_07642_, _07625_);
  or (_07644_, _07642_, word_in[24]);
  and (_26815_[0], _07644_, _07640_);
  or (_07645_, _07627_, _07194_);
  not (_07646_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_07648_, _07631_, _07646_);
  and (_07650_, _07631_, _06212_);
  nor (_07652_, _07650_, _07648_);
  nor (_07653_, _07652_, _07629_);
  and (_07655_, _07629_, word_in[9]);
  or (_07656_, _07655_, _07626_);
  or (_07658_, _07656_, _07653_);
  and (_07659_, _07658_, _07645_);
  or (_07660_, _07659_, _07625_);
  or (_07661_, _07642_, word_in[25]);
  and (_26815_[1], _07661_, _07660_);
  or (_07663_, _07627_, _07198_);
  not (_07665_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_07666_, _07631_, _07665_);
  and (_07668_, _07631_, _06227_);
  nor (_07669_, _07668_, _07666_);
  nor (_07670_, _07669_, _07629_);
  and (_07671_, _07629_, word_in[10]);
  or (_07672_, _07671_, _07626_);
  or (_07674_, _07672_, _07670_);
  and (_07675_, _07674_, _07663_);
  or (_07676_, _07675_, _07625_);
  or (_07677_, _07642_, word_in[26]);
  and (_26815_[2], _07677_, _07676_);
  or (_07680_, _07627_, _06247_);
  not (_07681_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_07683_, _07631_, _07681_);
  and (_07684_, _07631_, _06240_);
  nor (_07685_, _07684_, _07683_);
  nor (_07686_, _07685_, _07629_);
  and (_07687_, _07629_, word_in[11]);
  or (_07689_, _07687_, _07626_);
  or (_07690_, _07689_, _07686_);
  and (_07691_, _07690_, _07680_);
  or (_07693_, _07691_, _07625_);
  or (_07694_, _07642_, word_in[27]);
  and (_26815_[3], _07694_, _07693_);
  not (_07697_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_07698_, _07631_, _07697_);
  and (_07699_, _07631_, _06259_);
  nor (_07701_, _07699_, _07698_);
  nor (_07703_, _07701_, _07629_);
  and (_07704_, _07629_, word_in[12]);
  or (_07706_, _07704_, _07626_);
  or (_07708_, _07706_, _07703_);
  or (_07709_, _07627_, _07235_);
  and (_07711_, _07709_, _07708_);
  or (_07712_, _07711_, _07625_);
  or (_07713_, _07642_, word_in[28]);
  and (_26815_[4], _07713_, _07712_);
  or (_07714_, _07627_, _07268_);
  not (_07715_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_07717_, _07631_, _07715_);
  and (_07718_, _07631_, _06278_);
  nor (_07720_, _07718_, _07717_);
  nor (_07721_, _07720_, _07629_);
  and (_07722_, _07629_, word_in[13]);
  or (_07723_, _07722_, _07626_);
  or (_07724_, _07723_, _07721_);
  and (_07725_, _07724_, _07714_);
  or (_07726_, _07725_, _07625_);
  or (_07727_, _07642_, word_in[29]);
  and (_26815_[5], _07727_, _07726_);
  or (_07728_, _07627_, _07287_);
  not (_07729_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_07730_, _07631_, _07729_);
  and (_07731_, _07631_, _06294_);
  nor (_07732_, _07731_, _07730_);
  nor (_07733_, _07732_, _07629_);
  and (_07734_, _07629_, word_in[14]);
  or (_07735_, _07734_, _07626_);
  or (_07736_, _07735_, _07733_);
  and (_07737_, _07736_, _07728_);
  or (_07739_, _07737_, _07625_);
  or (_07740_, _07642_, word_in[30]);
  and (_26815_[6], _07740_, _07739_);
  or (_07741_, _07627_, _05415_);
  nor (_07743_, _07631_, _05187_);
  and (_07745_, _07631_, _05407_);
  nor (_07746_, _07745_, _07743_);
  nor (_07747_, _07746_, _07629_);
  and (_07749_, _07629_, word_in[15]);
  or (_07750_, _07749_, _07626_);
  or (_07752_, _07750_, _07747_);
  and (_07753_, _07752_, _07741_);
  or (_07754_, _07753_, _07625_);
  or (_07755_, _07642_, word_in[31]);
  and (_26815_[7], _07755_, _07754_);
  and (_07756_, _07346_, _05120_);
  and (_07757_, _05400_, _05133_);
  not (_07758_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_07759_, _07356_, _05403_);
  nor (_07760_, _07759_, _07758_);
  and (_07762_, _07759_, _06188_);
  nor (_07764_, _07762_, _07760_);
  nor (_07766_, _07764_, _07757_);
  and (_07768_, _05395_, _05246_);
  and (_07769_, _07757_, word_in[8]);
  or (_07770_, _07769_, _07768_);
  or (_07771_, _07770_, _07766_);
  not (_07772_, _07768_);
  or (_07773_, _07772_, _07174_);
  and (_07774_, _07773_, _07771_);
  or (_07775_, _07774_, _07756_);
  not (_07776_, _07756_);
  or (_07777_, _07776_, word_in[24]);
  and (_26816_[0], _07777_, _07775_);
  not (_07778_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_07779_, _07759_, _07778_);
  and (_07780_, _07759_, _06212_);
  nor (_07781_, _07780_, _07779_);
  nor (_07782_, _07781_, _07757_);
  and (_07783_, _07757_, word_in[9]);
  or (_07785_, _07783_, _07768_);
  or (_07786_, _07785_, _07782_);
  or (_07787_, _07772_, _07194_);
  and (_07788_, _07787_, _07786_);
  or (_07789_, _07788_, _07756_);
  or (_07790_, _07776_, word_in[25]);
  and (_26816_[1], _07790_, _07789_);
  not (_07791_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_07792_, _07759_, _07791_);
  and (_07793_, _07759_, _06227_);
  nor (_07794_, _07793_, _07792_);
  nor (_07795_, _07794_, _07757_);
  and (_07796_, _07757_, word_in[10]);
  or (_07797_, _07796_, _07768_);
  or (_07798_, _07797_, _07795_);
  or (_07799_, _07772_, _07198_);
  and (_07800_, _07799_, _07798_);
  or (_07802_, _07800_, _07756_);
  or (_07804_, _07776_, word_in[26]);
  and (_26816_[2], _07804_, _07802_);
  not (_07806_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_07807_, _07759_, _07806_);
  and (_07808_, _07759_, _06240_);
  nor (_07809_, _07808_, _07807_);
  nor (_07810_, _07809_, _07757_);
  and (_07811_, _07757_, word_in[11]);
  or (_07812_, _07811_, _07768_);
  or (_07813_, _07812_, _07810_);
  or (_07814_, _07772_, _06247_);
  and (_07815_, _07814_, _07813_);
  or (_07816_, _07815_, _07756_);
  or (_07817_, _07776_, word_in[27]);
  and (_26816_[3], _07817_, _07816_);
  not (_07818_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_07819_, _07759_, _07818_);
  and (_07820_, _07759_, _06259_);
  nor (_07821_, _07820_, _07819_);
  nor (_07822_, _07821_, _07757_);
  and (_07823_, _07757_, word_in[12]);
  or (_07824_, _07823_, _07768_);
  or (_07825_, _07824_, _07822_);
  or (_07826_, _07772_, _07235_);
  and (_07827_, _07826_, _07825_);
  or (_07828_, _07827_, _07756_);
  or (_07829_, _07776_, word_in[28]);
  and (_26816_[4], _07829_, _07828_);
  not (_07830_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_07831_, _07759_, _07830_);
  and (_07832_, _07759_, _06278_);
  nor (_07833_, _07832_, _07831_);
  nor (_07834_, _07833_, _07757_);
  and (_07835_, _07757_, word_in[13]);
  or (_07836_, _07835_, _07768_);
  or (_07837_, _07836_, _07834_);
  or (_07838_, _07772_, _07268_);
  and (_07839_, _07838_, _07837_);
  or (_07840_, _07839_, _07756_);
  or (_07841_, _07776_, word_in[29]);
  and (_26816_[5], _07841_, _07840_);
  not (_07842_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_07843_, _07759_, _07842_);
  and (_07844_, _07759_, _06294_);
  nor (_07845_, _07844_, _07843_);
  nor (_07846_, _07845_, _07757_);
  and (_07847_, _07757_, word_in[14]);
  or (_07848_, _07847_, _07768_);
  or (_07849_, _07848_, _07846_);
  or (_07850_, _07772_, _07287_);
  and (_07851_, _07850_, _07849_);
  or (_07852_, _07851_, _07756_);
  or (_07853_, _07776_, word_in[30]);
  and (_26816_[6], _07853_, _07852_);
  or (_07854_, _07772_, _05415_);
  nor (_07855_, _07759_, _05111_);
  and (_07856_, _07759_, _05407_);
  nor (_07857_, _07856_, _07855_);
  nor (_07858_, _07857_, _07757_);
  and (_07859_, _07757_, word_in[15]);
  or (_07860_, _07859_, _07768_);
  or (_07861_, _07860_, _07858_);
  and (_07862_, _07861_, _07854_);
  or (_07863_, _07862_, _07756_);
  or (_07864_, _07776_, word_in[31]);
  and (_26816_[7], _07864_, _07863_);
  and (_07865_, _23758_, _22781_);
  and (_07866_, _07865_, _24732_);
  and (_07867_, _01215_, _01152_);
  and (_07868_, _01231_, _01145_);
  and (_07869_, _01163_, _01146_);
  and (_07870_, _07869_, _01128_);
  or (_07871_, _07870_, _07868_);
  or (_07872_, _07871_, _07867_);
  and (_07873_, _01189_, _01128_);
  or (_07874_, _07873_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_07875_, _07874_, _07872_);
  and (_07876_, _07875_, _07866_);
  nor (_07877_, _07865_, _24732_);
  or (_07878_, _07877_, rst);
  or (_26834_[0], _07878_, _07876_);
  and (_07879_, _05834_, _23751_);
  and (_07880_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_02635_, _07880_, _07879_);
  nor (_07881_, _24989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_07882_, _07881_, _07326_);
  and (_07883_, _07882_, _24975_);
  and (_07884_, _25012_, _25000_);
  or (_07885_, _07884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not (_07886_, _07315_);
  and (_07887_, _07886_, _25003_);
  and (_07888_, _07887_, _07885_);
  or (_07890_, _24193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_07891_, _07890_, _24196_);
  nor (_07892_, _07891_, _07320_);
  or (_07893_, _07892_, _07888_);
  or (_07894_, _07893_, _07883_);
  or (_07895_, _07894_, _24192_);
  nand (_07896_, _24192_, _24047_);
  and (_07897_, _07896_, _24188_);
  and (_07898_, _07897_, _07895_);
  and (_07899_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_07900_, _07899_, _07898_);
  and (_02645_, _07900_, _22773_);
  and (_07901_, _05399_, _05912_);
  and (_07902_, _06180_, _05405_);
  and (_07903_, _07902_, word_in[0]);
  not (_07904_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_07905_, _07902_, _07904_);
  or (_07906_, _07905_, _07903_);
  or (_07907_, _07906_, _07901_);
  and (_07908_, _05394_, _05888_);
  not (_07909_, _07908_);
  not (_07910_, _07901_);
  or (_07911_, _07910_, word_in[8]);
  and (_07912_, _07911_, _07909_);
  and (_07913_, _07912_, _07907_);
  not (_07914_, _05316_);
  and (_07915_, _06785_, _07914_);
  and (_07916_, _07915_, _05151_);
  and (_07917_, _07908_, word_in[16]);
  or (_07918_, _07917_, _07916_);
  or (_07919_, _07918_, _07913_);
  not (_07920_, _07916_);
  or (_07921_, _07920_, _06810_);
  and (_26817_[0], _07921_, _07919_);
  nand (_07922_, _07902_, _06815_);
  or (_07923_, _07902_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_07924_, _07923_, _07922_);
  or (_07925_, _07924_, _07901_);
  or (_07926_, _07910_, word_in[9]);
  and (_07927_, _07926_, _07925_);
  or (_07928_, _07927_, _07908_);
  nor (_07929_, _07909_, word_in[17]);
  nor (_07930_, _07929_, _07916_);
  and (_07931_, _07930_, _07928_);
  and (_07932_, _07916_, _06207_);
  or (_26817_[1], _07932_, _07931_);
  or (_07933_, _07909_, word_in[18]);
  nand (_07934_, _07902_, _06827_);
  or (_07935_, _07902_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_07936_, _07935_, _07934_);
  or (_07937_, _07936_, _07901_);
  or (_07938_, _07910_, word_in[10]);
  and (_07939_, _07938_, _07937_);
  or (_07940_, _07939_, _07908_);
  and (_07941_, _07940_, _07933_);
  or (_07942_, _07941_, _07916_);
  or (_07943_, _07920_, _06842_);
  and (_26817_[2], _07943_, _07942_);
  nand (_07944_, _07902_, _06845_);
  or (_07945_, _07902_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_07946_, _07945_, _07944_);
  or (_07947_, _07946_, _07901_);
  or (_07948_, _07910_, word_in[11]);
  and (_07949_, _07948_, _07947_);
  or (_07950_, _07949_, _07908_);
  nor (_07951_, _07909_, word_in[19]);
  nor (_07952_, _07951_, _07916_);
  and (_07953_, _07952_, _07950_);
  and (_07954_, _07916_, _06861_);
  or (_26817_[3], _07954_, _07953_);
  or (_07955_, _07902_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand (_07956_, _07902_, _06864_);
  and (_07957_, _07956_, _07955_);
  or (_07958_, _07957_, _07901_);
  or (_07959_, _07910_, word_in[12]);
  and (_07960_, _07959_, _07958_);
  or (_07961_, _07960_, _07908_);
  or (_07962_, _07909_, word_in[20]);
  and (_07963_, _07962_, _07961_);
  or (_07964_, _07963_, _07916_);
  or (_07965_, _07920_, _06876_);
  and (_26817_[4], _07965_, _07964_);
  or (_07966_, _07909_, word_in[21]);
  nand (_07967_, _07902_, _06881_);
  or (_07968_, _07902_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_07969_, _07968_, _07967_);
  or (_07970_, _07969_, _07901_);
  or (_07971_, _07910_, word_in[13]);
  and (_07972_, _07971_, _07970_);
  or (_07973_, _07972_, _07908_);
  and (_07974_, _07973_, _07966_);
  or (_07975_, _07974_, _07916_);
  or (_07976_, _07920_, _06273_);
  and (_26817_[5], _07976_, _07975_);
  nand (_07977_, _07902_, _06900_);
  or (_07978_, _07902_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_07979_, _07978_, _07977_);
  or (_07980_, _07979_, _07901_);
  or (_07981_, _07910_, word_in[14]);
  and (_07982_, _07981_, _07980_);
  or (_07983_, _07982_, _07908_);
  nor (_07984_, _07909_, word_in[22]);
  nor (_07985_, _07984_, _07916_);
  and (_07986_, _07985_, _07983_);
  and (_07987_, _07916_, _06912_);
  or (_26817_[6], _07987_, _07986_);
  nor (_07988_, _07902_, _05224_);
  and (_07989_, _07902_, _05407_);
  or (_07990_, _07989_, _07988_);
  or (_07991_, _07990_, _07901_);
  or (_07992_, _07910_, word_in[15]);
  and (_07993_, _07992_, _07991_);
  or (_07994_, _07993_, _07908_);
  or (_07995_, _07909_, word_in[23]);
  and (_07996_, _07995_, _07994_);
  or (_07997_, _07996_, _07916_);
  or (_07998_, _07920_, _05387_);
  and (_26817_[7], _07998_, _07997_);
  and (_07999_, _25175_, _23890_);
  and (_08000_, _07999_, _23900_);
  not (_08001_, _07999_);
  and (_08002_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_02673_, _08002_, _08000_);
  and (_08003_, _07999_, _24053_);
  and (_08004_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_02678_, _08004_, _08003_);
  and (_08005_, _25175_, _24097_);
  and (_08006_, _08005_, _23920_);
  not (_08007_, _08005_);
  and (_08008_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_02690_, _08008_, _08006_);
  and (_08009_, _08005_, _23693_);
  and (_08010_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_02692_, _08010_, _08009_);
  and (_08011_, _25175_, _24068_);
  and (_08012_, _08011_, _23983_);
  not (_08013_, _08011_);
  and (_08014_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or (_02698_, _08014_, _08012_);
  and (_08015_, _08011_, _23715_);
  and (_08016_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or (_02703_, _08016_, _08015_);
  and (_08017_, _25175_, _23700_);
  and (_08018_, _08017_, _23715_);
  not (_08019_, _08017_);
  and (_08020_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or (_02713_, _08020_, _08018_);
  and (_08021_, _07915_, _05161_);
  and (_08022_, _06361_, _05393_);
  and (_08023_, _06351_, _05218_);
  not (_08025_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_08027_, _06354_, _05405_);
  nor (_08028_, _08027_, _08025_);
  and (_08030_, _08027_, _06188_);
  or (_08031_, _08030_, _08028_);
  or (_08032_, _08031_, _08023_);
  not (_08033_, _08023_);
  or (_08034_, _08033_, word_in[8]);
  and (_08035_, _08034_, _08032_);
  or (_08037_, _08035_, _08022_);
  not (_08038_, _08022_);
  or (_08040_, _08038_, _07174_);
  and (_08042_, _08040_, _08037_);
  or (_08043_, _08042_, _08021_);
  not (_08045_, _08021_);
  or (_08046_, _08045_, word_in[24]);
  and (_26818_[0], _08046_, _08043_);
  and (_08048_, _06005_, _23900_);
  and (_08049_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_27114_, _08049_, _08048_);
  not (_08052_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_08053_, _08027_, _08052_);
  and (_08054_, _08027_, _06212_);
  nor (_08056_, _08054_, _08053_);
  nor (_08057_, _08056_, _08023_);
  and (_08058_, _08023_, word_in[9]);
  or (_08059_, _08058_, _08057_);
  and (_08060_, _08059_, _08038_);
  and (_08061_, _08022_, _07194_);
  or (_08062_, _08061_, _08021_);
  or (_08063_, _08062_, _08060_);
  or (_08064_, _08045_, word_in[25]);
  and (_26818_[1], _08064_, _08063_);
  not (_08065_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_08066_, _08027_, _08065_);
  and (_08067_, _08027_, _06227_);
  nor (_08068_, _08067_, _08066_);
  nor (_08069_, _08068_, _08023_);
  and (_08070_, _08023_, word_in[10]);
  or (_08071_, _08070_, _08069_);
  and (_08072_, _08071_, _08038_);
  and (_08073_, _08022_, _07198_);
  or (_08074_, _08073_, _08021_);
  or (_08075_, _08074_, _08072_);
  or (_08076_, _08045_, word_in[26]);
  and (_26818_[2], _08076_, _08075_);
  not (_08077_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_08078_, _08027_, _08077_);
  and (_08079_, _08027_, _06240_);
  nor (_08080_, _08079_, _08078_);
  nor (_08081_, _08080_, _08023_);
  and (_08082_, _08023_, word_in[11]);
  or (_08083_, _08082_, _08081_);
  and (_08084_, _08083_, _08038_);
  and (_08085_, _08022_, _06247_);
  or (_08086_, _08085_, _08021_);
  or (_08087_, _08086_, _08084_);
  or (_08088_, _08045_, word_in[27]);
  and (_26818_[3], _08088_, _08087_);
  not (_08089_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_08090_, _08027_, _08089_);
  and (_08091_, _08027_, _06259_);
  or (_08092_, _08091_, _08090_);
  or (_08093_, _08092_, _08023_);
  or (_08094_, _08033_, word_in[12]);
  and (_08095_, _08094_, _08093_);
  or (_08096_, _08095_, _08022_);
  or (_08097_, _08038_, _07235_);
  and (_08098_, _08097_, _08096_);
  or (_08099_, _08098_, _08021_);
  or (_08100_, _08045_, word_in[28]);
  and (_26818_[4], _08100_, _08099_);
  and (_08101_, _05878_, _23920_);
  and (_08102_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_02729_, _08102_, _08101_);
  not (_08103_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_08104_, _08027_, _08103_);
  and (_08105_, _08027_, _06278_);
  nor (_08106_, _08105_, _08104_);
  nor (_08107_, _08106_, _08023_);
  and (_08108_, _08023_, word_in[13]);
  or (_08109_, _08108_, _08107_);
  and (_08111_, _08109_, _08038_);
  and (_08112_, _08022_, _07268_);
  or (_08113_, _08112_, _08021_);
  or (_08114_, _08113_, _08111_);
  or (_08115_, _08045_, word_in[29]);
  and (_26818_[5], _08115_, _08114_);
  or (_08117_, _08038_, _07287_);
  not (_08118_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_08119_, _08027_, _08118_);
  and (_08120_, _08027_, _06294_);
  or (_08121_, _08120_, _08119_);
  or (_08122_, _08121_, _08023_);
  or (_08124_, _08033_, word_in[14]);
  and (_08126_, _08124_, _08122_);
  or (_08127_, _08126_, _08022_);
  and (_08128_, _08127_, _08117_);
  or (_08130_, _08128_, _08021_);
  or (_08131_, _08045_, word_in[30]);
  and (_26818_[6], _08131_, _08130_);
  nor (_08133_, _08027_, _05099_);
  and (_08134_, _08027_, _05407_);
  nor (_08135_, _08134_, _08133_);
  nor (_08137_, _08135_, _08023_);
  and (_08138_, _08023_, word_in[15]);
  or (_08140_, _08138_, _08137_);
  and (_08141_, _08140_, _08038_);
  and (_08143_, _08022_, _05415_);
  or (_08144_, _08143_, _08021_);
  or (_08145_, _08144_, _08141_);
  or (_08146_, _08045_, word_in[31]);
  and (_26818_[7], _08146_, _08145_);
  and (_08147_, _05878_, _24053_);
  and (_08149_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_02743_, _08149_, _08147_);
  and (_08151_, _05859_, _24027_);
  and (_08152_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  or (_02747_, _08152_, _08151_);
  and (_08153_, _05859_, _23751_);
  and (_08155_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  or (_02757_, _08155_, _08153_);
  and (_08157_, _05726_, _23900_);
  and (_08158_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_02770_, _08158_, _08157_);
  and (_08159_, _05726_, _24053_);
  and (_08161_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_02774_, _08161_, _08159_);
  and (_08163_, _02531_, _23920_);
  and (_08164_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  or (_02781_, _08164_, _08163_);
  and (_08165_, _02531_, _23693_);
  and (_08167_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  or (_02784_, _08167_, _08165_);
  and (_08168_, _02464_, _23983_);
  and (_08170_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  or (_02788_, _08170_, _08168_);
  and (_08171_, _02464_, _23715_);
  and (_08173_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  or (_02793_, _08173_, _08171_);
  and (_08174_, _06497_, _05393_);
  and (_08175_, _06487_, _05218_);
  and (_08176_, _06491_, _05405_);
  nand (_08177_, _08176_, _06797_);
  or (_08178_, _08176_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_08179_, _08178_, _08177_);
  or (_08180_, _08179_, _08175_);
  not (_08181_, _08175_);
  or (_08182_, _08181_, word_in[8]);
  and (_08183_, _08182_, _08180_);
  or (_08184_, _08183_, _08174_);
  and (_08185_, _07915_, _05123_);
  not (_08186_, _08174_);
  nor (_08187_, _08186_, _07174_);
  nor (_08188_, _08187_, _08185_);
  and (_08189_, _08188_, _08184_);
  and (_08190_, _08185_, word_in[24]);
  or (_26819_[0], _08190_, _08189_);
  nand (_08191_, _08176_, _06815_);
  or (_08192_, _08176_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_08193_, _08192_, _08191_);
  or (_08194_, _08193_, _08175_);
  or (_08195_, _08181_, word_in[9]);
  and (_08196_, _08195_, _08194_);
  or (_08197_, _08196_, _08174_);
  nor (_08198_, _08186_, _07194_);
  nor (_08199_, _08198_, _08185_);
  and (_08200_, _08199_, _08197_);
  and (_08201_, _08185_, word_in[25]);
  or (_26819_[1], _08201_, _08200_);
  nand (_08202_, _08176_, _06827_);
  or (_08203_, _08176_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_08204_, _08203_, _08202_);
  nor (_08205_, _08204_, _08175_);
  and (_08206_, _08175_, word_in[10]);
  or (_08207_, _08206_, _08205_);
  or (_08208_, _08207_, _08174_);
  nor (_08209_, _08186_, _07198_);
  nor (_08210_, _08209_, _08185_);
  and (_08211_, _08210_, _08208_);
  and (_08212_, _08185_, word_in[26]);
  or (_26819_[2], _08212_, _08211_);
  and (_08213_, _01759_, _24027_);
  and (_08214_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  or (_27112_, _08214_, _08213_);
  not (_08215_, _08185_);
  or (_08216_, _08186_, _06247_);
  or (_08217_, _08176_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nand (_08218_, _08176_, _06845_);
  and (_08219_, _08218_, _08217_);
  or (_08220_, _08219_, _08175_);
  or (_08221_, _08181_, word_in[11]);
  and (_08222_, _08221_, _08220_);
  or (_08223_, _08222_, _08174_);
  and (_08224_, _08223_, _08216_);
  and (_08225_, _08224_, _08215_);
  and (_08226_, _08185_, word_in[27]);
  or (_26819_[3], _08226_, _08225_);
  and (_08227_, _02829_, _23900_);
  and (_08228_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or (_02804_, _08228_, _08227_);
  or (_08229_, _08186_, _07235_);
  nand (_08230_, _08176_, _06864_);
  or (_08231_, _08176_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_08232_, _08231_, _08230_);
  or (_08233_, _08232_, _08175_);
  or (_08234_, _08181_, word_in[12]);
  and (_08235_, _08234_, _08233_);
  or (_08236_, _08235_, _08174_);
  and (_08237_, _08236_, _08229_);
  or (_08238_, _08237_, _08185_);
  or (_08239_, _08215_, word_in[28]);
  and (_26819_[4], _08239_, _08238_);
  and (_08240_, _23706_, _23444_);
  and (_08241_, _08240_, _23751_);
  not (_08242_, _08240_);
  and (_08243_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_02808_, _08243_, _08241_);
  nand (_08244_, _08176_, _06881_);
  or (_08245_, _08176_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_08246_, _08245_, _08244_);
  or (_08247_, _08246_, _08175_);
  or (_08248_, _08181_, word_in[13]);
  and (_08249_, _08248_, _08247_);
  or (_08250_, _08249_, _08174_);
  nor (_08251_, _08186_, _07268_);
  nor (_08252_, _08251_, _08185_);
  and (_08253_, _08252_, _08250_);
  and (_08254_, _08185_, word_in[29]);
  or (_26819_[5], _08254_, _08253_);
  and (_08255_, _01759_, _23751_);
  and (_08256_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  or (_02812_, _08256_, _08255_);
  or (_08257_, _08186_, _07287_);
  nand (_08258_, _08176_, _06900_);
  or (_08259_, _08176_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_08260_, _08259_, _08258_);
  or (_08261_, _08260_, _08175_);
  or (_08262_, _08181_, word_in[14]);
  and (_08263_, _08262_, _08261_);
  or (_08264_, _08263_, _08174_);
  and (_08265_, _08264_, _08257_);
  or (_08266_, _08265_, _08185_);
  or (_08267_, _08215_, word_in[30]);
  and (_26819_[6], _08267_, _08266_);
  or (_08268_, _08186_, _05415_);
  nor (_08269_, _08176_, _05219_);
  and (_08270_, _08176_, _05407_);
  or (_08271_, _08270_, _08269_);
  or (_08272_, _08271_, _08175_);
  or (_08273_, _08181_, word_in[15]);
  and (_08274_, _08273_, _08272_);
  or (_08275_, _08274_, _08174_);
  and (_08276_, _08275_, _08268_);
  or (_08277_, _08276_, _08185_);
  or (_08278_, _08215_, word_in[31]);
  and (_26819_[7], _08278_, _08277_);
  and (_08279_, _23910_, _23900_);
  and (_08280_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_02824_, _08280_, _08279_);
  and (_08281_, _25176_, _23751_);
  and (_08282_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or (_02830_, _08282_, _08281_);
  and (_08283_, _07999_, _24027_);
  and (_08284_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_02834_, _08284_, _08283_);
  and (_08285_, _07999_, _23693_);
  and (_08286_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_27118_, _08286_, _08285_);
  and (_08287_, _08005_, _23983_);
  and (_08288_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_27117_, _08288_, _08287_);
  and (_08289_, _08240_, _24053_);
  and (_08290_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_02852_, _08290_, _08289_);
  and (_08291_, _08011_, _24053_);
  and (_08292_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or (_02854_, _08292_, _08291_);
  and (_08293_, _08017_, _24053_);
  and (_08294_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or (_02859_, _08294_, _08293_);
  and (_08295_, _06005_, _23751_);
  and (_08296_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_02868_, _08296_, _08295_);
  and (_08297_, _05878_, _23693_);
  and (_08298_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_02875_, _08298_, _08297_);
  and (_08299_, _05859_, _23715_);
  and (_08300_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  or (_02878_, _08300_, _08299_);
  and (_08301_, _23910_, _23751_);
  and (_08302_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_02881_, _08302_, _08301_);
  not (_08303_, _05401_);
  or (_08304_, _08303_, word_in[8]);
  not (_08305_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_08306_, _05406_, _08305_);
  and (_08307_, _06188_, _05406_);
  or (_08308_, _08307_, _08306_);
  or (_08309_, _08308_, _05401_);
  and (_08310_, _08309_, _08304_);
  or (_08311_, _08310_, _05396_);
  or (_08312_, _07174_, _05398_);
  and (_08313_, _08312_, _08311_);
  and (_08314_, _08313_, _05392_);
  and (_08315_, _05390_, word_in[24]);
  or (_26820_[0], _08315_, _08314_);
  and (_08316_, _05726_, _24027_);
  and (_08317_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_27104_, _08317_, _08316_);
  and (_08318_, _05390_, word_in[25]);
  not (_08319_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_08320_, _05406_, _08319_);
  and (_08321_, _06212_, _05406_);
  or (_08322_, _08321_, _08320_);
  or (_08323_, _08322_, _05401_);
  or (_08324_, _08303_, word_in[9]);
  and (_08325_, _08324_, _08323_);
  or (_08326_, _08325_, _05396_);
  or (_08327_, _07194_, _05398_);
  and (_08328_, _08327_, _05392_);
  and (_08329_, _08328_, _08326_);
  or (_26820_[1], _08329_, _08318_);
  and (_08330_, _05726_, _23693_);
  and (_08331_, _05728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_02887_, _08331_, _08330_);
  or (_08332_, _08303_, word_in[10]);
  not (_08333_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_08334_, _05406_, _08333_);
  and (_08335_, _06227_, _05406_);
  or (_08336_, _08335_, _08334_);
  or (_08337_, _08336_, _05401_);
  and (_08338_, _08337_, _08332_);
  or (_08339_, _08338_, _05396_);
  or (_08340_, _07198_, _05398_);
  and (_08341_, _08340_, _08339_);
  and (_08342_, _08341_, _05392_);
  and (_08343_, _05390_, word_in[26]);
  or (_26820_[2], _08343_, _08342_);
  and (_08344_, _02531_, _23983_);
  and (_08345_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  or (_02890_, _08345_, _08344_);
  not (_08346_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_08347_, _05406_, _08346_);
  and (_08348_, _06240_, _05406_);
  or (_08349_, _08348_, _08347_);
  or (_08350_, _08349_, _05401_);
  or (_08351_, _08303_, word_in[11]);
  and (_08352_, _08351_, _08350_);
  or (_08353_, _08352_, _05396_);
  or (_08354_, _06247_, _05398_);
  and (_08355_, _08354_, _05392_);
  and (_08356_, _08355_, _08353_);
  and (_08357_, _05390_, word_in[27]);
  or (_26820_[3], _08357_, _08356_);
  and (_08358_, _05390_, word_in[28]);
  not (_08359_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_08360_, _05406_, _08359_);
  and (_08361_, _06259_, _05406_);
  or (_08362_, _08361_, _08360_);
  or (_08363_, _08362_, _05401_);
  or (_08364_, _08303_, word_in[12]);
  and (_08365_, _08364_, _08363_);
  or (_08366_, _08365_, _05396_);
  or (_08367_, _07235_, _05398_);
  and (_08368_, _08367_, _05392_);
  and (_08369_, _08368_, _08366_);
  or (_26820_[4], _08369_, _08358_);
  not (_08370_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_08371_, _05406_, _08370_);
  and (_08372_, _06278_, _05406_);
  or (_08373_, _08372_, _08371_);
  or (_08374_, _08373_, _05401_);
  or (_08375_, _08303_, word_in[13]);
  and (_08376_, _08375_, _08374_);
  or (_08377_, _08376_, _05396_);
  or (_08378_, _07268_, _05398_);
  and (_08379_, _08378_, _05392_);
  and (_08380_, _08379_, _08377_);
  and (_08381_, _05390_, word_in[29]);
  or (_26820_[5], _08381_, _08380_);
  and (_08382_, _06294_, _05406_);
  not (_08383_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_08384_, _05406_, _08383_);
  nor (_08385_, _08384_, _08382_);
  nor (_08387_, _08385_, _05401_);
  and (_08388_, _05401_, word_in[14]);
  or (_08390_, _08388_, _08387_);
  and (_08391_, _08390_, _05398_);
  and (_08393_, _07287_, _05396_);
  or (_08395_, _08393_, _08391_);
  and (_08396_, _08395_, _05392_);
  and (_08397_, _05390_, word_in[30]);
  or (_26820_[6], _08397_, _08396_);
  and (_08400_, _02464_, _24053_);
  and (_08401_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  or (_02915_, _08401_, _08400_);
  and (_08402_, _24237_, _24157_);
  and (_08404_, _08402_, _23751_);
  not (_08405_, _08402_);
  and (_08407_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_27060_, _08407_, _08404_);
  and (_08408_, _01759_, _23715_);
  and (_08409_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  or (_27111_, _08409_, _08408_);
  and (_08410_, _24027_, _23910_);
  and (_08411_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_02946_, _08411_, _08410_);
  and (_08413_, _08402_, _24053_);
  and (_08415_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_02948_, _08415_, _08413_);
  and (_08416_, _04901_, _23983_);
  and (_08417_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or (_02955_, _08417_, _08416_);
  and (_08418_, _05834_, _23715_);
  and (_08419_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_02961_, _08419_, _08418_);
  and (_08421_, _06005_, _23983_);
  and (_08422_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_02965_, _08422_, _08421_);
  and (_08423_, _08005_, _23715_);
  and (_08424_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_02969_, _08424_, _08423_);
  and (_08425_, _08011_, _23900_);
  and (_08426_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or (_02972_, _08426_, _08425_);
  and (_08427_, _08017_, _23900_);
  and (_08428_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or (_27116_, _08428_, _08427_);
  and (_08429_, _06005_, _23920_);
  and (_08430_, _06007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_02979_, _08430_, _08429_);
  and (_08431_, _05878_, _24027_);
  and (_08432_, _05881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_27113_, _08432_, _08431_);
  and (_08433_, _24053_, _23988_);
  and (_08434_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_02987_, _08434_, _08433_);
  and (_08435_, _23890_, _23706_);
  and (_08436_, _08435_, _23900_);
  not (_08437_, _08435_);
  and (_08438_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or (_02990_, _08438_, _08436_);
  and (_08439_, _05859_, _23983_);
  and (_08440_, _05862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  or (_02993_, _08440_, _08439_);
  nor (_08441_, _05063_, _06797_);
  nand (_08442_, _04985_, _06642_);
  or (_08443_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_08444_, _08443_, _08442_);
  and (_08445_, _08444_, _05009_);
  or (_08446_, _08445_, _04991_);
  nand (_08447_, _04985_, _06929_);
  or (_08448_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_08449_, _08448_, _08447_);
  and (_08450_, _08449_, _05006_);
  nand (_08451_, _04985_, _07157_);
  or (_08452_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_08453_, _08452_, _08451_);
  and (_08454_, _08453_, _05016_);
  nand (_08455_, _04985_, _06353_);
  or (_08456_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_08457_, _08456_, _08455_);
  and (_08458_, _08457_, _05027_);
  or (_08459_, _08458_, _08454_);
  or (_08460_, _08459_, _08450_);
  or (_08461_, _08460_, _08446_);
  nand (_08462_, _04985_, _07758_);
  or (_08463_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_08464_, _08463_, _08462_);
  and (_08465_, _08464_, _05009_);
  or (_08466_, _08465_, _05091_);
  nand (_08467_, _04985_, _08305_);
  or (_08468_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_08469_, _08468_, _08467_);
  and (_08470_, _08469_, _05016_);
  nand (_08471_, _04985_, _08025_);
  or (_08472_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_08473_, _08472_, _08471_);
  and (_08474_, _08473_, _05006_);
  or (_08475_, _08474_, _08470_);
  nand (_08476_, _04985_, _07498_);
  or (_08477_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_08478_, _08477_, _08476_);
  and (_08479_, _08478_, _05027_);
  or (_08480_, _08479_, _08475_);
  or (_08481_, _08480_, _08466_);
  and (_08482_, _08481_, _08461_);
  and (_08483_, _08482_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _08483_, _08441_);
  nor (_08484_, _05063_, _06815_);
  nand (_08485_, _04985_, _06376_);
  or (_08486_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_08487_, _08486_, _08485_);
  and (_08488_, _08487_, _05027_);
  or (_08489_, _08488_, _04991_);
  nand (_08490_, _04985_, _06944_);
  or (_08491_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_08492_, _08491_, _08490_);
  and (_08493_, _08492_, _05006_);
  nand (_08494_, _04985_, _07185_);
  or (_08495_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_08496_, _08495_, _08494_);
  and (_08497_, _08496_, _05016_);
  nand (_08498_, _04985_, _06664_);
  or (_08499_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_08500_, _08499_, _08498_);
  and (_08501_, _08500_, _05009_);
  or (_08502_, _08501_, _08497_);
  or (_08503_, _08502_, _08493_);
  or (_08504_, _08503_, _08489_);
  nand (_08505_, _04985_, _07520_);
  or (_08506_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_08507_, _08506_, _08505_);
  and (_08508_, _08507_, _05027_);
  or (_08509_, _08508_, _05091_);
  nand (_08510_, _04985_, _08052_);
  or (_08511_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_08512_, _08511_, _08510_);
  and (_08513_, _08512_, _05006_);
  nand (_08514_, _04985_, _08319_);
  or (_08515_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_08516_, _08515_, _08514_);
  and (_08517_, _08516_, _05016_);
  nand (_08518_, _04985_, _07778_);
  or (_08519_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_08520_, _08519_, _08518_);
  and (_08521_, _08520_, _05009_);
  or (_08522_, _08521_, _08517_);
  or (_08523_, _08522_, _08513_);
  or (_08524_, _08523_, _08509_);
  and (_08525_, _08524_, _08504_);
  and (_08526_, _08525_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _08526_, _08484_);
  nor (_08527_, _05063_, _06827_);
  nand (_08528_, _04985_, _06391_);
  or (_08529_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_08530_, _08529_, _08528_);
  and (_08531_, _08530_, _05027_);
  or (_08532_, _08531_, _04991_);
  nand (_08533_, _04985_, _06958_);
  or (_08534_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_08535_, _08534_, _08533_);
  and (_08536_, _08535_, _05006_);
  nand (_08537_, _04985_, _07200_);
  or (_08538_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_08539_, _08538_, _08537_);
  and (_08540_, _08539_, _05016_);
  nand (_08541_, _04985_, _06686_);
  or (_08542_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_08543_, _08542_, _08541_);
  and (_08544_, _08543_, _05009_);
  or (_08545_, _08544_, _08540_);
  or (_08546_, _08545_, _08536_);
  or (_08547_, _08546_, _08532_);
  nand (_08548_, _04985_, _07531_);
  or (_08549_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_08550_, _08549_, _08548_);
  and (_08551_, _08550_, _05027_);
  or (_08552_, _08551_, _05091_);
  nand (_08553_, _04985_, _08065_);
  or (_08555_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_08556_, _08555_, _08553_);
  and (_08557_, _08556_, _05006_);
  nand (_08558_, _04985_, _08333_);
  or (_08559_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_08560_, _08559_, _08558_);
  and (_08561_, _08560_, _05016_);
  nand (_08562_, _04985_, _07791_);
  or (_08563_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_08564_, _08563_, _08562_);
  and (_08565_, _08564_, _05009_);
  or (_08566_, _08565_, _08561_);
  or (_08567_, _08566_, _08557_);
  or (_08568_, _08567_, _08552_);
  and (_08569_, _08568_, _08547_);
  and (_08570_, _08569_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _08570_, _08527_);
  nor (_08571_, _05063_, _06845_);
  nand (_08572_, _04985_, _06703_);
  or (_08573_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_08574_, _08573_, _08572_);
  and (_08575_, _08574_, _05009_);
  or (_08576_, _08575_, _04991_);
  nand (_08578_, _04985_, _06972_);
  or (_08579_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_08580_, _08579_, _08578_);
  and (_08581_, _08580_, _05006_);
  nand (_08582_, _04985_, _07218_);
  or (_08583_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_08584_, _08583_, _08582_);
  and (_08585_, _08584_, _05016_);
  nand (_08586_, _04985_, _06404_);
  or (_08587_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_08588_, _08587_, _08586_);
  and (_08589_, _08588_, _05027_);
  or (_08590_, _08589_, _08585_);
  or (_08591_, _08590_, _08581_);
  or (_08592_, _08591_, _08576_);
  nand (_08594_, _04985_, _07806_);
  or (_08595_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_08596_, _08595_, _08594_);
  and (_08597_, _08596_, _05009_);
  or (_08598_, _08597_, _05091_);
  nand (_08599_, _04985_, _08346_);
  or (_08600_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_08601_, _08600_, _08599_);
  and (_08602_, _08601_, _05016_);
  nand (_08603_, _04985_, _08077_);
  or (_08605_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_08606_, _08605_, _08603_);
  and (_08607_, _08606_, _05006_);
  or (_08608_, _08607_, _08602_);
  nand (_08609_, _04985_, _07549_);
  or (_08610_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_08611_, _08610_, _08609_);
  and (_08612_, _08611_, _05027_);
  or (_08613_, _08612_, _08608_);
  or (_08614_, _08613_, _08598_);
  and (_08615_, _08614_, _08592_);
  and (_08616_, _08615_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _08616_, _08571_);
  nor (_08618_, _05063_, _06864_);
  nand (_08619_, _04985_, _06716_);
  or (_08620_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_08621_, _08620_, _08619_);
  and (_08622_, _08621_, _05009_);
  or (_08623_, _08622_, _04991_);
  nand (_08624_, _04985_, _06987_);
  or (_08625_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_08626_, _08625_, _08624_);
  and (_08627_, _08626_, _05006_);
  nand (_08628_, _04985_, _07238_);
  or (_08629_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_08630_, _08629_, _08628_);
  and (_08631_, _08630_, _05016_);
  nand (_08632_, _04985_, _06419_);
  or (_08633_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_08634_, _08633_, _08632_);
  and (_08635_, _08634_, _05027_);
  or (_08636_, _08635_, _08631_);
  or (_08637_, _08636_, _08627_);
  or (_08638_, _08637_, _08623_);
  nand (_08639_, _04985_, _07818_);
  or (_08640_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_08641_, _08640_, _08639_);
  and (_08642_, _08641_, _05009_);
  or (_08643_, _08642_, _05091_);
  nand (_08644_, _04985_, _08359_);
  or (_08645_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_08646_, _08645_, _08644_);
  and (_08647_, _08646_, _05016_);
  nand (_08648_, _04985_, _08089_);
  or (_08650_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_08651_, _08650_, _08648_);
  and (_08652_, _08651_, _05006_);
  or (_08653_, _08652_, _08647_);
  nand (_08654_, _04985_, _07561_);
  or (_08655_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_08656_, _08655_, _08654_);
  and (_08657_, _08656_, _05027_);
  or (_08658_, _08657_, _08653_);
  or (_08659_, _08658_, _08643_);
  and (_08660_, _08659_, _08638_);
  and (_08661_, _08660_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _08661_, _08618_);
  nor (_08662_, _05063_, _06881_);
  nand (_08664_, _04985_, _06728_);
  or (_08665_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_08666_, _08665_, _08664_);
  and (_08668_, _08666_, _05009_);
  or (_08669_, _08668_, _04991_);
  nand (_08670_, _04985_, _07000_);
  or (_08671_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_08672_, _08671_, _08670_);
  and (_08673_, _08672_, _05006_);
  nand (_08674_, _04985_, _07257_);
  or (_08675_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_08676_, _08675_, _08674_);
  and (_08677_, _08676_, _05016_);
  nand (_08678_, _04985_, _06430_);
  or (_08679_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_08680_, _08679_, _08678_);
  and (_08681_, _08680_, _05027_);
  or (_08682_, _08681_, _08677_);
  or (_08683_, _08682_, _08673_);
  or (_08684_, _08683_, _08669_);
  nand (_08686_, _04985_, _07830_);
  or (_08687_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_08688_, _08687_, _08686_);
  and (_08690_, _08688_, _05009_);
  or (_08691_, _08690_, _05091_);
  nand (_08692_, _04985_, _08370_);
  or (_08693_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_08694_, _08693_, _08692_);
  and (_08695_, _08694_, _05016_);
  nand (_08696_, _04985_, _08103_);
  or (_08697_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_08698_, _08697_, _08696_);
  and (_08699_, _08698_, _05006_);
  or (_08700_, _08699_, _08695_);
  nand (_08701_, _04985_, _07581_);
  or (_08703_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_08704_, _08703_, _08701_);
  and (_08705_, _08704_, _05027_);
  or (_08706_, _08705_, _08700_);
  or (_08708_, _08706_, _08691_);
  and (_08709_, _08708_, _08684_);
  and (_08710_, _08709_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _08710_, _08662_);
  nor (_08711_, _05063_, _06900_);
  nand (_08712_, _04985_, _06447_);
  or (_08713_, _04985_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_08714_, _08713_, _08712_);
  and (_08715_, _08714_, _05027_);
  or (_08716_, _08715_, _04991_);
  nand (_08717_, _04985_, _07013_);
  or (_08718_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_08719_, _08718_, _08717_);
  and (_08720_, _08719_, _05006_);
  nand (_08721_, _04985_, _07279_);
  or (_08722_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_08723_, _08722_, _08721_);
  and (_08724_, _08723_, _05016_);
  nand (_08725_, _04985_, _06745_);
  or (_08726_, _04985_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_08727_, _08726_, _08725_);
  and (_08728_, _08727_, _05009_);
  or (_08730_, _08728_, _08724_);
  or (_08731_, _08730_, _08720_);
  or (_08732_, _08731_, _08716_);
  nand (_08733_, _04985_, _07597_);
  or (_08734_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_08735_, _08734_, _08733_);
  and (_08736_, _08735_, _05027_);
  or (_08737_, _08736_, _05091_);
  nand (_08738_, _04985_, _08118_);
  or (_08739_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_08740_, _08739_, _08738_);
  and (_08741_, _08740_, _05006_);
  nand (_08742_, _04985_, _08383_);
  or (_08743_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_08744_, _08743_, _08742_);
  and (_08745_, _08744_, _05016_);
  nand (_08746_, _04985_, _07842_);
  or (_08747_, _04985_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_08748_, _08747_, _08746_);
  and (_08749_, _08748_, _05009_);
  or (_08750_, _08749_, _08745_);
  or (_08751_, _08750_, _08741_);
  or (_08752_, _08751_, _08737_);
  and (_08753_, _08752_, _08732_);
  and (_08754_, _08753_, _05063_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _08754_, _08711_);
  and (_08755_, _05170_, word_in[8]);
  nand (_08756_, _04985_, _06489_);
  or (_08757_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_08758_, _08757_, _08756_);
  and (_08759_, _08758_, _05173_);
  nand (_08760_, _04985_, _06178_);
  or (_08761_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_08762_, _08761_, _08760_);
  and (_08763_, _08762_, _05172_);
  or (_08764_, _08763_, _08759_);
  and (_08765_, _08764_, _05135_);
  nand (_08766_, _04985_, _07630_);
  or (_08767_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_08768_, _08767_, _08766_);
  and (_08769_, _08768_, _05173_);
  and (_08770_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_08771_, _04985_, _07498_);
  or (_08772_, _08771_, _08770_);
  and (_08773_, _08772_, _05172_);
  or (_08774_, _08773_, _08769_);
  and (_08775_, _08774_, _05133_);
  and (_08776_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_08777_, _04985_, _07157_);
  or (_08778_, _08777_, _08776_);
  and (_08779_, _08778_, _05173_);
  and (_08780_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_08781_, _04985_, _06929_);
  or (_08782_, _08781_, _08780_);
  and (_08783_, _08782_, _05172_);
  or (_08784_, _08783_, _08779_);
  and (_08785_, _08784_, _05202_);
  and (_08786_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_08787_, _04985_, _08305_);
  or (_08788_, _08787_, _08786_);
  and (_08789_, _08788_, _05173_);
  nand (_08791_, _04985_, _07904_);
  or (_08792_, _04985_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_08793_, _08792_, _08791_);
  and (_08794_, _08793_, _05172_);
  or (_08795_, _08794_, _08789_);
  and (_08796_, _08795_, _05218_);
  or (_08797_, _08796_, _08785_);
  or (_08798_, _08797_, _08775_);
  nor (_08799_, _08798_, _08765_);
  nor (_08800_, _08799_, _05170_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _08800_, _08755_);
  and (_08801_, _05170_, word_in[9]);
  nand (_08802_, _04985_, _06508_);
  or (_08803_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_08804_, _08803_, _08802_);
  and (_08805_, _08804_, _05173_);
  nand (_08806_, _04985_, _06209_);
  or (_08807_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_08808_, _08807_, _08806_);
  and (_08809_, _08808_, _05172_);
  or (_08810_, _08809_, _08805_);
  and (_08811_, _08810_, _05135_);
  nand (_08813_, _04985_, _07646_);
  or (_08814_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_08815_, _08814_, _08813_);
  and (_08816_, _08815_, _05173_);
  and (_08818_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_08819_, _04985_, _07520_);
  or (_08820_, _08819_, _08818_);
  and (_08821_, _08820_, _05172_);
  or (_08822_, _08821_, _08816_);
  and (_08823_, _08822_, _05133_);
  and (_08824_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_08825_, _04985_, _07185_);
  or (_08826_, _08825_, _08824_);
  and (_08827_, _08826_, _05173_);
  and (_08828_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_08829_, _04985_, _06944_);
  or (_08830_, _08829_, _08828_);
  and (_08831_, _08830_, _05172_);
  or (_08832_, _08831_, _08827_);
  and (_08833_, _08832_, _05202_);
  and (_08834_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_08835_, _04985_, _08319_);
  or (_08836_, _08835_, _08834_);
  and (_08837_, _08836_, _05173_);
  and (_08838_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_08839_, _04985_, _08052_);
  or (_08840_, _08839_, _08838_);
  and (_08841_, _08840_, _05172_);
  or (_08842_, _08841_, _08837_);
  and (_08843_, _08842_, _05218_);
  or (_08844_, _08843_, _08833_);
  or (_08845_, _08844_, _08823_);
  nor (_08846_, _08845_, _08811_);
  nor (_08847_, _08846_, _05170_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _08847_, _08801_);
  and (_08848_, _05170_, word_in[10]);
  nand (_08849_, _04985_, _06522_);
  or (_08850_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_08851_, _08850_, _08849_);
  and (_08852_, _08851_, _05173_);
  nand (_08853_, _04985_, _06225_);
  or (_08855_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_08856_, _08855_, _08853_);
  and (_08857_, _08856_, _05172_);
  or (_08858_, _08857_, _08852_);
  and (_08859_, _08858_, _05135_);
  nand (_08860_, _04985_, _07665_);
  or (_08861_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_08862_, _08861_, _08860_);
  and (_08863_, _08862_, _05173_);
  and (_08864_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_08865_, _04985_, _07531_);
  or (_08866_, _08865_, _08864_);
  and (_08867_, _08866_, _05172_);
  or (_08868_, _08867_, _08863_);
  and (_08869_, _08868_, _05133_);
  and (_08870_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_08871_, _04985_, _07200_);
  or (_08872_, _08871_, _08870_);
  and (_08873_, _08872_, _05173_);
  and (_08874_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_08875_, _04985_, _06958_);
  or (_08876_, _08875_, _08874_);
  and (_08877_, _08876_, _05172_);
  or (_08878_, _08877_, _08873_);
  and (_08879_, _08878_, _05202_);
  and (_08880_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_08881_, _04985_, _08333_);
  or (_08882_, _08881_, _08880_);
  and (_08883_, _08882_, _05173_);
  and (_08885_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_08887_, _04985_, _08065_);
  or (_08888_, _08887_, _08885_);
  and (_08889_, _08888_, _05172_);
  or (_08890_, _08889_, _08883_);
  and (_08891_, _08890_, _05218_);
  or (_08892_, _08891_, _08879_);
  or (_08893_, _08892_, _08869_);
  nor (_08894_, _08893_, _08859_);
  nor (_08896_, _08894_, _05170_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _08896_, _08848_);
  and (_08897_, _05170_, word_in[11]);
  nand (_08898_, _04985_, _06539_);
  or (_08899_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_08900_, _08899_, _08898_);
  and (_08901_, _08900_, _05173_);
  nand (_08902_, _04985_, _06238_);
  or (_08903_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_08904_, _08903_, _08902_);
  and (_08905_, _08904_, _05172_);
  or (_08906_, _08905_, _08901_);
  and (_08907_, _08906_, _05135_);
  nand (_08908_, _04985_, _07681_);
  or (_08909_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_08910_, _08909_, _08908_);
  and (_08911_, _08910_, _05173_);
  and (_08913_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_08915_, _04985_, _07549_);
  or (_08916_, _08915_, _08913_);
  and (_08918_, _08916_, _05172_);
  or (_08919_, _08918_, _08911_);
  and (_08921_, _08919_, _05133_);
  and (_08922_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_08923_, _04985_, _07218_);
  or (_08924_, _08923_, _08922_);
  and (_08926_, _08924_, _05173_);
  and (_08928_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_08929_, _04985_, _06972_);
  or (_08931_, _08929_, _08928_);
  and (_08932_, _08931_, _05172_);
  or (_08933_, _08932_, _08926_);
  and (_08935_, _08933_, _05202_);
  and (_08936_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_08937_, _04985_, _08346_);
  or (_08939_, _08937_, _08936_);
  and (_08940_, _08939_, _05173_);
  and (_08941_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_08942_, _04985_, _08077_);
  or (_08943_, _08942_, _08941_);
  and (_08944_, _08943_, _05172_);
  or (_08945_, _08944_, _08940_);
  and (_08946_, _08945_, _05218_);
  or (_08947_, _08946_, _08935_);
  or (_08948_, _08947_, _08921_);
  nor (_08949_, _08948_, _08907_);
  nor (_08951_, _08949_, _05170_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _08951_, _08897_);
  and (_08952_, _05170_, word_in[12]);
  nand (_08953_, _04985_, _06553_);
  or (_08954_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_08955_, _08954_, _08953_);
  and (_08956_, _08955_, _05173_);
  nand (_08957_, _04985_, _06257_);
  or (_08958_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_08959_, _08958_, _08957_);
  and (_08960_, _08959_, _05172_);
  or (_08961_, _08960_, _08956_);
  and (_08962_, _08961_, _05135_);
  nand (_08964_, _04985_, _07697_);
  or (_08965_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_08966_, _08965_, _08964_);
  and (_08967_, _08966_, _05173_);
  and (_08968_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_08969_, _04985_, _07561_);
  or (_08970_, _08969_, _08968_);
  and (_08971_, _08970_, _05172_);
  or (_08972_, _08971_, _08967_);
  and (_08974_, _08972_, _05133_);
  and (_08975_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_08976_, _04985_, _07238_);
  or (_08977_, _08976_, _08975_);
  and (_08978_, _08977_, _05173_);
  and (_08980_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_08981_, _04985_, _06987_);
  or (_08983_, _08981_, _08980_);
  and (_08984_, _08983_, _05172_);
  or (_08985_, _08984_, _08978_);
  and (_08986_, _08985_, _05202_);
  and (_08987_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_08988_, _04985_, _08359_);
  or (_08990_, _08988_, _08987_);
  and (_08992_, _08990_, _05173_);
  and (_08993_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_08994_, _04985_, _08089_);
  or (_08995_, _08994_, _08993_);
  and (_08996_, _08995_, _05172_);
  or (_08997_, _08996_, _08992_);
  and (_08998_, _08997_, _05218_);
  or (_08999_, _08998_, _08986_);
  or (_09000_, _08999_, _08974_);
  nor (_09001_, _09000_, _08962_);
  nor (_09002_, _09001_, _05170_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _09002_, _08952_);
  and (_09003_, _05170_, word_in[13]);
  nand (_09004_, _04985_, _06569_);
  or (_09005_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_09006_, _09005_, _09004_);
  and (_09007_, _09006_, _05173_);
  nand (_09008_, _04985_, _06275_);
  or (_09011_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_09012_, _09011_, _09008_);
  and (_09014_, _09012_, _05172_);
  or (_09016_, _09014_, _09007_);
  and (_09017_, _09016_, _05135_);
  nand (_09018_, _04985_, _07715_);
  or (_09020_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_09021_, _09020_, _09018_);
  and (_09023_, _09021_, _05173_);
  and (_09024_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_09026_, _04985_, _07581_);
  or (_09027_, _09026_, _09024_);
  and (_09028_, _09027_, _05172_);
  or (_09030_, _09028_, _09023_);
  and (_09031_, _09030_, _05133_);
  and (_09033_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_09035_, _04985_, _07257_);
  or (_09036_, _09035_, _09033_);
  and (_09037_, _09036_, _05173_);
  and (_09038_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_09039_, _04985_, _07000_);
  or (_09040_, _09039_, _09038_);
  and (_09041_, _09040_, _05172_);
  or (_09042_, _09041_, _09037_);
  and (_09043_, _09042_, _05202_);
  and (_09044_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_09046_, _04985_, _08370_);
  or (_09047_, _09046_, _09044_);
  and (_09048_, _09047_, _05173_);
  and (_09049_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_09050_, _04985_, _08103_);
  or (_09051_, _09050_, _09049_);
  and (_09052_, _09051_, _05172_);
  or (_09053_, _09052_, _09048_);
  and (_09054_, _09053_, _05218_);
  or (_09055_, _09054_, _09043_);
  or (_09056_, _09055_, _09031_);
  nor (_09057_, _09056_, _09017_);
  nor (_09058_, _09057_, _05170_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _09058_, _09003_);
  and (_09059_, _05170_, word_in[14]);
  nand (_09060_, _04985_, _06582_);
  or (_09061_, _04985_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_09062_, _09061_, _09060_);
  and (_09063_, _09062_, _05173_);
  nand (_09064_, _04985_, _06291_);
  or (_09065_, _04985_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_09066_, _09065_, _09064_);
  and (_09067_, _09066_, _05172_);
  or (_09068_, _09067_, _09063_);
  and (_09069_, _09068_, _05135_);
  nand (_09070_, _04985_, _07729_);
  or (_09071_, _04985_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_09072_, _09071_, _09070_);
  and (_09074_, _09072_, _05173_);
  and (_09075_, _04985_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_09076_, _04985_, _07597_);
  or (_09077_, _09076_, _09075_);
  and (_09078_, _09077_, _05172_);
  or (_09079_, _09078_, _09074_);
  and (_09080_, _09079_, _05133_);
  and (_09081_, _04985_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_09082_, _04985_, _07279_);
  or (_09084_, _09082_, _09081_);
  and (_09086_, _09084_, _05173_);
  and (_09087_, _04985_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_09088_, _04985_, _07013_);
  or (_09089_, _09088_, _09087_);
  and (_09090_, _09089_, _05172_);
  or (_09091_, _09090_, _09086_);
  and (_09093_, _09091_, _05202_);
  and (_09094_, _04985_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_09095_, _04985_, _08383_);
  or (_09096_, _09095_, _09094_);
  and (_09097_, _09096_, _05173_);
  and (_09098_, _04985_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_09099_, _04985_, _08118_);
  or (_09100_, _09099_, _09098_);
  and (_09101_, _09100_, _05172_);
  or (_09102_, _09101_, _09097_);
  and (_09103_, _09102_, _05218_);
  or (_09105_, _09103_, _09093_);
  or (_09106_, _09105_, _09080_);
  nor (_09107_, _09106_, _09069_);
  nor (_09109_, _09107_, _05170_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _09109_, _09059_);
  and (_09111_, _02531_, _23715_);
  and (_09112_, _02533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  or (_03041_, _09112_, _09111_);
  and (_09113_, _02464_, _23900_);
  and (_09115_, _02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  or (_27102_, _09115_, _09113_);
  and (_09116_, _01759_, _23983_);
  and (_09117_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  or (_03045_, _09117_, _09116_);
  and (_09119_, _05278_, word_in[16]);
  and (_09120_, _08449_, _05009_);
  and (_09121_, _08457_, _05016_);
  or (_09122_, _09121_, _09120_);
  and (_09123_, _08453_, _05006_);
  and (_09124_, _08444_, _05027_);
  or (_09125_, _09124_, _09123_);
  or (_09126_, _09125_, _09122_);
  or (_09127_, _09126_, _05241_);
  and (_09129_, _08473_, _05009_);
  and (_09130_, _08478_, _05016_);
  or (_09132_, _09130_, _09129_);
  and (_09133_, _08469_, _05006_);
  and (_09135_, _08464_, _05027_);
  or (_09136_, _09135_, _09133_);
  or (_09138_, _09136_, _09132_);
  or (_09139_, _09138_, _05289_);
  nand (_09140_, _09139_, _09127_);
  nor (_09141_, _09140_, _05278_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _09141_, _09119_);
  and (_09143_, _05278_, word_in[17]);
  and (_09144_, _08487_, _05016_);
  and (_09145_, _08496_, _05006_);
  or (_09146_, _09145_, _09144_);
  and (_09148_, _08492_, _05009_);
  and (_09150_, _08500_, _05027_);
  or (_09152_, _09150_, _09148_);
  or (_09153_, _09152_, _09146_);
  or (_09154_, _09153_, _05241_);
  and (_09156_, _08512_, _05009_);
  and (_09158_, _08507_, _05016_);
  or (_09159_, _09158_, _09156_);
  and (_09160_, _08516_, _05006_);
  and (_09161_, _08520_, _05027_);
  or (_09163_, _09161_, _09160_);
  or (_09164_, _09163_, _09159_);
  or (_09166_, _09164_, _05289_);
  nand (_09168_, _09166_, _09154_);
  nor (_09170_, _09168_, _05278_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _09170_, _09143_);
  and (_09172_, _05278_, word_in[18]);
  and (_09174_, _08535_, _05009_);
  and (_09175_, _08530_, _05016_);
  or (_09176_, _09175_, _09174_);
  and (_09177_, _08539_, _05006_);
  and (_09178_, _08543_, _05027_);
  or (_09179_, _09178_, _09177_);
  or (_09180_, _09179_, _09176_);
  or (_09181_, _09180_, _05241_);
  and (_09182_, _08550_, _05016_);
  and (_09183_, _08560_, _05006_);
  or (_09184_, _09183_, _09182_);
  and (_09185_, _08556_, _05009_);
  and (_09186_, _08564_, _05027_);
  or (_09188_, _09186_, _09185_);
  or (_09189_, _09188_, _09184_);
  or (_09191_, _09189_, _05289_);
  nand (_09192_, _09191_, _09181_);
  nor (_09193_, _09192_, _05278_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _09193_, _09172_);
  and (_09194_, _05278_, word_in[19]);
  and (_09195_, _08580_, _05009_);
  and (_09196_, _08588_, _05016_);
  or (_09197_, _09196_, _09195_);
  and (_09198_, _08584_, _05006_);
  and (_09199_, _08574_, _05027_);
  or (_09201_, _09199_, _09198_);
  or (_09202_, _09201_, _09197_);
  or (_09203_, _09202_, _05241_);
  and (_09204_, _08606_, _05009_);
  and (_09205_, _08611_, _05016_);
  or (_09206_, _09205_, _09204_);
  and (_09207_, _08601_, _05006_);
  and (_09209_, _08596_, _05027_);
  or (_09210_, _09209_, _09207_);
  or (_09211_, _09210_, _09206_);
  or (_09212_, _09211_, _05289_);
  nand (_09213_, _09212_, _09203_);
  nor (_09214_, _09213_, _05278_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _09214_, _09194_);
  and (_09215_, _05278_, word_in[20]);
  and (_09216_, _08626_, _05009_);
  and (_09217_, _08634_, _05016_);
  or (_09218_, _09217_, _09216_);
  and (_09219_, _08630_, _05006_);
  and (_09220_, _08621_, _05027_);
  or (_09221_, _09220_, _09219_);
  or (_09222_, _09221_, _09218_);
  or (_09223_, _09222_, _05241_);
  and (_09224_, _08651_, _05009_);
  and (_09225_, _08656_, _05016_);
  or (_09226_, _09225_, _09224_);
  and (_09227_, _08646_, _05006_);
  and (_09228_, _08641_, _05027_);
  or (_09229_, _09228_, _09227_);
  or (_09230_, _09229_, _09226_);
  or (_09232_, _09230_, _05289_);
  nand (_09233_, _09232_, _09223_);
  nor (_09234_, _09233_, _05278_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _09234_, _09215_);
  and (_09236_, _05278_, word_in[21]);
  and (_09237_, _08672_, _05009_);
  and (_09238_, _08680_, _05016_);
  or (_09239_, _09238_, _09237_);
  and (_09240_, _08676_, _05006_);
  and (_09242_, _08666_, _05027_);
  or (_09243_, _09242_, _09240_);
  or (_09244_, _09243_, _09239_);
  or (_09246_, _09244_, _05241_);
  and (_09247_, _08698_, _05009_);
  and (_09248_, _08704_, _05016_);
  or (_09250_, _09248_, _09247_);
  and (_09252_, _08694_, _05006_);
  and (_09253_, _08688_, _05027_);
  or (_09254_, _09253_, _09252_);
  or (_09256_, _09254_, _09250_);
  or (_09257_, _09256_, _05289_);
  nand (_09258_, _09257_, _09246_);
  nor (_09259_, _09258_, _05278_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _09259_, _09236_);
  and (_09260_, _05278_, word_in[22]);
  and (_09261_, _08719_, _05009_);
  and (_09262_, _08714_, _05016_);
  or (_09263_, _09262_, _09261_);
  and (_09264_, _08723_, _05006_);
  and (_09266_, _08727_, _05027_);
  or (_09267_, _09266_, _09264_);
  or (_09269_, _09267_, _09263_);
  or (_09270_, _09269_, _05241_);
  and (_09271_, _08740_, _05009_);
  and (_09272_, _08735_, _05016_);
  or (_09273_, _09272_, _09271_);
  and (_09274_, _08744_, _05006_);
  and (_09276_, _08748_, _05027_);
  or (_09277_, _09276_, _09274_);
  or (_09278_, _09277_, _09273_);
  or (_09279_, _09278_, _05289_);
  nand (_09281_, _09279_, _09270_);
  nor (_09282_, _09281_, _05278_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _09282_, _09260_);
  and (_09284_, _05349_, word_in[24]);
  and (_09285_, _08772_, _05173_);
  and (_09286_, _08768_, _05172_);
  or (_09287_, _09286_, _09285_);
  and (_09288_, _09287_, _05317_);
  and (_09289_, _08762_, _05173_);
  and (_09290_, _08758_, _05172_);
  or (_09292_, _09290_, _09289_);
  and (_09294_, _09292_, _05324_);
  and (_09295_, _08782_, _05173_);
  and (_09297_, _08778_, _05172_);
  or (_09298_, _09297_, _09295_);
  and (_09299_, _09298_, _05359_);
  and (_09300_, _08793_, _05173_);
  and (_09301_, _08788_, _05172_);
  or (_09303_, _09301_, _09300_);
  and (_09304_, _09303_, _05369_);
  or (_09306_, _09304_, _09299_);
  or (_09308_, _09306_, _09294_);
  nor (_09310_, _09308_, _09288_);
  nor (_09312_, _09310_, _05349_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _09312_, _09284_);
  and (_09314_, _05349_, word_in[25]);
  and (_09315_, _08820_, _05173_);
  and (_09316_, _08815_, _05172_);
  or (_09318_, _09316_, _09315_);
  and (_09320_, _09318_, _05317_);
  and (_09322_, _08808_, _05173_);
  and (_09323_, _08804_, _05172_);
  or (_09324_, _09323_, _09322_);
  and (_09325_, _09324_, _05324_);
  and (_09327_, _08830_, _05173_);
  and (_09328_, _08826_, _05172_);
  or (_09329_, _09328_, _09327_);
  and (_09330_, _09329_, _05359_);
  and (_09332_, _08840_, _05173_);
  and (_09333_, _08836_, _05172_);
  or (_09334_, _09333_, _09332_);
  and (_09335_, _09334_, _05369_);
  or (_09336_, _09335_, _09330_);
  or (_09337_, _09336_, _09325_);
  nor (_09338_, _09337_, _09320_);
  nor (_09339_, _09338_, _05349_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _09339_, _09314_);
  and (_09340_, _05349_, word_in[26]);
  and (_09341_, _08856_, _05173_);
  and (_09342_, _08851_, _05172_);
  or (_09343_, _09342_, _09341_);
  and (_09344_, _09343_, _05324_);
  and (_09345_, _08866_, _05173_);
  and (_09346_, _08862_, _05172_);
  or (_09347_, _09346_, _09345_);
  and (_09348_, _09347_, _05317_);
  and (_09349_, _08876_, _05173_);
  and (_09350_, _08872_, _05172_);
  or (_09352_, _09350_, _09349_);
  and (_09353_, _09352_, _05359_);
  and (_09354_, _08888_, _05173_);
  and (_09355_, _08882_, _05172_);
  or (_09356_, _09355_, _09354_);
  and (_09357_, _09356_, _05369_);
  or (_09358_, _09357_, _09353_);
  or (_09359_, _09358_, _09348_);
  nor (_09360_, _09359_, _09344_);
  nor (_09361_, _09360_, _05349_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _09361_, _09340_);
  and (_09362_, _05349_, word_in[27]);
  and (_09364_, _08916_, _05173_);
  and (_09365_, _08910_, _05172_);
  or (_09366_, _09365_, _09364_);
  and (_09367_, _09366_, _05317_);
  and (_09368_, _08904_, _05173_);
  and (_09370_, _08900_, _05172_);
  or (_09371_, _09370_, _09368_);
  and (_09372_, _09371_, _05324_);
  and (_09374_, _08931_, _05173_);
  and (_09375_, _08924_, _05172_);
  or (_09376_, _09375_, _09374_);
  and (_09377_, _09376_, _05359_);
  and (_09378_, _08943_, _05173_);
  and (_09379_, _08939_, _05172_);
  or (_09381_, _09379_, _09378_);
  and (_09382_, _09381_, _05369_);
  or (_09383_, _09382_, _09377_);
  or (_09384_, _09383_, _09372_);
  nor (_09385_, _09384_, _09367_);
  nor (_09386_, _09385_, _05349_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _09386_, _09362_);
  and (_09388_, _05349_, word_in[28]);
  and (_09389_, _08959_, _05173_);
  and (_09390_, _08955_, _05172_);
  or (_09391_, _09390_, _09389_);
  and (_09392_, _09391_, _05324_);
  and (_09393_, _08970_, _05173_);
  and (_09394_, _08966_, _05172_);
  or (_09395_, _09394_, _09393_);
  and (_09396_, _09395_, _05317_);
  and (_09397_, _08983_, _05173_);
  and (_09398_, _08977_, _05172_);
  or (_09399_, _09398_, _09397_);
  and (_09400_, _09399_, _05359_);
  and (_09401_, _08995_, _05173_);
  and (_09402_, _08990_, _05172_);
  or (_09403_, _09402_, _09401_);
  and (_09404_, _09403_, _05369_);
  or (_09405_, _09404_, _09400_);
  or (_09406_, _09405_, _09396_);
  nor (_09407_, _09406_, _09392_);
  nor (_09408_, _09407_, _05349_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _09408_, _09388_);
  and (_09409_, _05349_, word_in[29]);
  and (_09410_, _09012_, _05173_);
  and (_09411_, _09006_, _05172_);
  or (_09412_, _09411_, _09410_);
  and (_09413_, _09412_, _05324_);
  and (_09414_, _09027_, _05173_);
  and (_09415_, _09021_, _05172_);
  or (_09416_, _09415_, _09414_);
  and (_09417_, _09416_, _05317_);
  and (_09418_, _09040_, _05173_);
  and (_09419_, _09036_, _05172_);
  or (_09420_, _09419_, _09418_);
  and (_09421_, _09420_, _05359_);
  and (_09422_, _09051_, _05173_);
  and (_09423_, _09047_, _05172_);
  or (_09424_, _09423_, _09422_);
  and (_09425_, _09424_, _05369_);
  or (_09426_, _09425_, _09421_);
  or (_09427_, _09426_, _09417_);
  nor (_09428_, _09427_, _09413_);
  nor (_09429_, _09428_, _05349_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _09429_, _09409_);
  and (_09430_, _05349_, word_in[30]);
  and (_09431_, _09077_, _05173_);
  and (_09432_, _09072_, _05172_);
  or (_09434_, _09432_, _09431_);
  and (_09435_, _09434_, _05317_);
  and (_09436_, _09066_, _05173_);
  and (_09437_, _09062_, _05172_);
  or (_09438_, _09437_, _09436_);
  and (_09439_, _09438_, _05324_);
  and (_09440_, _09089_, _05173_);
  and (_09441_, _09084_, _05172_);
  or (_09442_, _09441_, _09440_);
  and (_09443_, _09442_, _05359_);
  and (_09444_, _09100_, _05173_);
  and (_09445_, _09096_, _05172_);
  or (_09446_, _09445_, _09444_);
  and (_09448_, _09446_, _05369_);
  or (_09449_, _09448_, _09443_);
  or (_09450_, _09449_, _09439_);
  nor (_09451_, _09450_, _09435_);
  nor (_09452_, _09451_, _05349_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _09452_, _09430_);
  and (_09453_, _25176_, _23693_);
  and (_09454_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or (_03129_, _09454_, _09453_);
  and (_09455_, _04901_, _24053_);
  and (_09456_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_03144_, _09456_, _09455_);
  and (_09457_, _23910_, _23693_);
  and (_09458_, _23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_03177_, _09458_, _09457_);
  and (_09459_, _08017_, _23751_);
  and (_09460_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or (_03187_, _09460_, _09459_);
  and (_09461_, _08017_, _23920_);
  and (_09462_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or (_03193_, _09462_, _09461_);
  and (_09463_, _24237_, _23890_);
  and (_09465_, _09463_, _23715_);
  not (_09466_, _09463_);
  and (_09467_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_27054_, _09467_, _09465_);
  nand (_09468_, _25868_, _22773_);
  nor (_26880_, _09468_, _25871_);
  and (_09469_, _24305_, _23751_);
  and (_09470_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or (_27047_, _09470_, _09469_);
  and (_09471_, _08017_, _23693_);
  and (_09472_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or (_03245_, _09472_, _09471_);
  and (_09475_, _07087_, _23751_);
  and (_09476_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_03248_, _09476_, _09475_);
  and (_09478_, _08017_, _24027_);
  and (_09479_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or (_03254_, _09479_, _09478_);
  and (_09480_, _24145_, _23719_);
  and (_09481_, _09480_, _23693_);
  not (_09482_, _09480_);
  and (_09483_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or (_03257_, _09483_, _09481_);
  and (_09485_, _23905_, _23719_);
  and (_09486_, _09485_, _23920_);
  not (_09487_, _09485_);
  and (_09488_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_03264_, _09488_, _09486_);
  and (_09489_, _02337_, _23983_);
  and (_09490_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_03269_, _09490_, _09489_);
  and (_09491_, _02337_, _23751_);
  and (_09492_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_03272_, _09492_, _09491_);
  and (_09493_, _04901_, _23715_);
  and (_09494_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or (_03281_, _09494_, _09493_);
  and (_09495_, _02509_, _23693_);
  and (_09496_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_03284_, _09496_, _09495_);
  and (_09497_, _01932_, _23920_);
  and (_09498_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_03286_, _09498_, _09497_);
  and (_09499_, _04901_, _23693_);
  and (_09500_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or (_03291_, _09500_, _09499_);
  and (_09501_, _01701_, _23983_);
  and (_09502_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or (_03304_, _09502_, _09501_);
  and (_09503_, _24098_, _24053_);
  and (_09504_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or (_03308_, _09504_, _09503_);
  and (_09505_, _04901_, _23751_);
  and (_09506_, _04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or (_27059_, _09506_, _09505_);
  and (_09507_, _24157_, _23453_);
  and (_09508_, _09507_, _23983_);
  not (_09509_, _09507_);
  and (_09510_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_03317_, _09510_, _09508_);
  and (_09511_, _25169_, _23693_);
  and (_09512_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_03320_, _09512_, _09511_);
  and (_09513_, _23900_, _23721_);
  and (_09514_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_03328_, _09514_, _09513_);
  and (_09515_, _05834_, _23693_);
  and (_09516_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_03348_, _09516_, _09515_);
  and (_09517_, _24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_09518_, _24085_, _23715_);
  or (_03372_, _09518_, _09517_);
  and (_09519_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and (_09520_, _24146_, _24027_);
  or (_03381_, _09520_, _09519_);
  and (_09522_, _07087_, _23983_);
  and (_09523_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_03409_, _09523_, _09522_);
  and (_09524_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_09525_, _25153_, _23983_);
  or (_03434_, _09525_, _09524_);
  and (_09526_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_09527_, _25153_, _23751_);
  or (_03437_, _09527_, _09526_);
  and (_09528_, _08402_, _23900_);
  and (_09529_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_03439_, _09529_, _09528_);
  and (_09530_, _25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  and (_09531_, _25308_, _23715_);
  or (_27005_, _09531_, _09530_);
  and (_09532_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_09533_, _25490_, _24053_);
  or (_03457_, _09533_, _09532_);
  and (_09534_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_09535_, _01768_, _23900_);
  or (_26997_, _09535_, _09534_);
  and (_09537_, _08402_, _23715_);
  and (_09538_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_03464_, _09538_, _09537_);
  and (_09540_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and (_09541_, _02170_, _23983_);
  or (_03470_, _09541_, _09540_);
  and (_09542_, _08402_, _23693_);
  and (_09543_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_03472_, _09543_, _09542_);
  and (_09544_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and (_09545_, _02170_, _23715_);
  or (_03475_, _09545_, _09544_);
  and (_09546_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and (_09547_, _02362_, _23715_);
  or (_03480_, _09547_, _09546_);
  and (_09548_, _09507_, _24027_);
  and (_09549_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_03505_, _09549_, _09548_);
  and (_09550_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_09551_, _02499_, _23920_);
  or (_26986_, _09551_, _09550_);
  and (_09552_, _23891_, _23444_);
  and (_09553_, _09552_, _23900_);
  not (_09554_, _09552_);
  and (_09555_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_03519_, _09555_, _09553_);
  and (_09556_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and (_09557_, _24275_, _24053_);
  or (_03536_, _09557_, _09556_);
  and (_09558_, _25364_, _23693_);
  and (_09559_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or (_03542_, _09559_, _09558_);
  and (_09560_, _08402_, _24027_);
  and (_09561_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_03545_, _09561_, _09560_);
  and (_09562_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_09563_, _02752_, _23751_);
  or (_03553_, _09563_, _09562_);
  and (_09564_, _02753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_09565_, _02752_, _24027_);
  or (_03575_, _09565_, _09564_);
  and (_09566_, _24238_, _23983_);
  and (_09567_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or (_03577_, _09567_, _09566_);
  and (_09568_, _08402_, _23920_);
  and (_09569_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_03579_, _09569_, _09568_);
  and (_09570_, _24237_, _24097_);
  and (_09572_, _09570_, _24053_);
  not (_09574_, _09570_);
  and (_09575_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_03591_, _09575_, _09572_);
  and (_09576_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and (_09577_, _24795_, _23715_);
  or (_03663_, _09577_, _09576_);
  and (_09578_, _23906_, _22856_);
  and (_09579_, _09578_, _23890_);
  not (_09580_, _09579_);
  and (_09581_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_09582_, _09579_, _24053_);
  or (_03678_, _09582_, _09581_);
  and (_09583_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and (_09584_, _24275_, _23900_);
  or (_03691_, _09584_, _09583_);
  and (_09585_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_09586_, _02687_, _24027_);
  or (_03693_, _09586_, _09585_);
  and (_09587_, _24901_, _24053_);
  and (_09588_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_03722_, _09588_, _09587_);
  and (_09589_, _02248_, _23920_);
  and (_09590_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or (_03726_, _09590_, _09589_);
  and (_09592_, _01932_, _24027_);
  and (_09593_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_03729_, _09593_, _09592_);
  and (_09595_, _07087_, _24027_);
  and (_09596_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_03744_, _09596_, _09595_);
  and (_09597_, _09578_, _24061_);
  not (_09598_, _09597_);
  and (_09599_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_09600_, _09597_, _23920_);
  or (_03799_, _09600_, _09599_);
  and (_09601_, _09552_, _24027_);
  and (_09602_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_03822_, _09602_, _09601_);
  and (_09603_, _09578_, _24108_);
  not (_09604_, _09603_);
  and (_09605_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and (_09606_, _09603_, _24027_);
  or (_03833_, _09606_, _09605_);
  and (_09608_, _24235_, _23909_);
  and (_09609_, _09608_, _23983_);
  not (_09610_, _09608_);
  and (_09611_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_03850_, _09611_, _09609_);
  and (_09612_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_09613_, _09597_, _23751_);
  or (_03863_, _09613_, _09612_);
  and (_09614_, _09608_, _23900_);
  and (_09615_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_03866_, _09615_, _09614_);
  and (_09616_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_09617_, _09597_, _23693_);
  or (_03868_, _09617_, _09616_);
  and (_09618_, _09608_, _23751_);
  and (_09619_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_03876_, _09619_, _09618_);
  and (_09620_, _09578_, _24235_);
  not (_09621_, _09620_);
  and (_09622_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  and (_09624_, _09620_, _23751_);
  or (_03889_, _09624_, _09622_);
  and (_09625_, _23909_, _23890_);
  and (_09626_, _09625_, _23715_);
  not (_09627_, _09625_);
  and (_09628_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  or (_03899_, _09628_, _09626_);
  and (_09629_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  and (_09630_, _09620_, _23715_);
  or (_03901_, _09630_, _09629_);
  and (_09631_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and (_09632_, _09620_, _23920_);
  or (_03915_, _09632_, _09631_);
  and (_09634_, _24097_, _23909_);
  and (_09635_, _09634_, _23715_);
  not (_09636_, _09634_);
  and (_09637_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  or (_03932_, _09637_, _09635_);
  and (_09638_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  and (_09639_, _09620_, _24027_);
  or (_03937_, _09639_, _09638_);
  and (_09640_, _09634_, _24053_);
  and (_09641_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  or (_03947_, _09641_, _09640_);
  and (_09642_, _24068_, _23909_);
  and (_09643_, _09642_, _23920_);
  not (_09644_, _09642_);
  and (_09645_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_27091_, _09645_, _09643_);
  and (_09647_, _09578_, _24123_);
  not (_09648_, _09647_);
  and (_09649_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  and (_09650_, _09647_, _24053_);
  or (_03966_, _09650_, _09649_);
  and (_09651_, _09642_, _23693_);
  and (_09652_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_03969_, _09652_, _09651_);
  and (_09653_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and (_09654_, _09647_, _23693_);
  or (_03972_, _09654_, _09653_);
  and (_09655_, _06631_, _23900_);
  and (_09656_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or (_03981_, _09656_, _09655_);
  and (_09657_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  and (_09658_, _09647_, _23900_);
  or (_03984_, _09658_, _09657_);
  and (_09660_, _23909_, _23700_);
  and (_09662_, _09660_, _23715_);
  not (_09663_, _09660_);
  and (_09664_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_03995_, _09664_, _09662_);
  and (_09665_, _09552_, _23920_);
  and (_09666_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_04003_, _09666_, _09665_);
  and (_09667_, _09660_, _23751_);
  and (_09668_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_04005_, _09668_, _09667_);
  and (_09669_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  and (_09670_, _09647_, _23920_);
  or (_04009_, _09670_, _09669_);
  and (_09671_, _08017_, _23983_);
  and (_09672_, _08019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or (_04011_, _09672_, _09671_);
  and (_09673_, _08011_, _23751_);
  and (_09674_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or (_04013_, _09674_, _09673_);
  and (_09676_, _23938_, _23909_);
  and (_09677_, _09676_, _23693_);
  not (_09678_, _09676_);
  and (_09679_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  or (_04026_, _09679_, _09677_);
  nand (_09680_, _24192_, _24017_);
  not (_09681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_09683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_09684_, _24989_, _24202_);
  or (_09685_, _09684_, _09683_);
  or (_09686_, _09685_, _09682_);
  nand (_09687_, _09686_, _09681_);
  and (_09688_, _24990_, _24975_);
  and (_09690_, _09688_, _09687_);
  and (_09691_, _24203_, _24193_);
  and (_09692_, _09691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_09693_, _09692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_09694_, _24995_);
  and (_09695_, _09694_, _24196_);
  and (_09696_, _09695_, _09693_);
  or (_09697_, _25014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_09698_, _25015_);
  and (_09699_, _09698_, _25003_);
  and (_09700_, _09699_, _09697_);
  or (_09701_, _09700_, _09696_);
  or (_09702_, _09701_, _09690_);
  or (_09703_, _09702_, _24192_);
  and (_09704_, _09703_, _24188_);
  and (_09705_, _09704_, _09680_);
  and (_09706_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_09707_, _09706_, _09705_);
  and (_04028_, _09707_, _22773_);
  nand (_09709_, _02481_, _23357_);
  and (_09710_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_09711_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_09712_, _09711_, _09710_);
  or (_09713_, _09712_, _02481_);
  and (_09714_, _09713_, _05576_);
  and (_09715_, _09714_, _09709_);
  and (_09716_, _02473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_09717_, _09716_, _09715_);
  and (_04031_, _09717_, _22773_);
  and (_09718_, _24237_, _24145_);
  and (_09719_, _09718_, _23900_);
  not (_09720_, _09718_);
  and (_09721_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_04034_, _09721_, _09719_);
  and (_09722_, _09578_, _24157_);
  not (_09723_, _09722_);
  and (_09724_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_09725_, _09722_, _23751_);
  or (_04037_, _09725_, _09724_);
  and (_09726_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_09727_, _09722_, _23715_);
  or (_04043_, _09727_, _09726_);
  and (_09728_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_09729_, _09722_, _23900_);
  or (_04048_, _09729_, _09728_);
  and (_09730_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_09731_, _09722_, _23983_);
  or (_04055_, _09731_, _09730_);
  and (_09732_, _24274_, _24237_);
  and (_09733_, _09732_, _24027_);
  not (_09734_, _09732_);
  and (_09735_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_27081_, _09735_, _09733_);
  and (_09736_, _09732_, _23900_);
  and (_09737_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_04068_, _09737_, _09736_);
  and (_09738_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and (_09739_, _09603_, _24053_);
  or (_04079_, _09739_, _09738_);
  and (_09740_, _24237_, _23905_);
  and (_09741_, _09740_, _23900_);
  not (_09742_, _09740_);
  and (_09743_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or (_04084_, _09743_, _09741_);
  and (_09744_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  and (_09745_, _09603_, _23693_);
  or (_04086_, _09745_, _09744_);
  or (_09746_, _05576_, _23413_);
  and (_09747_, _05646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_09748_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_09749_, _09748_, _09747_);
  or (_09750_, _09749_, _02473_);
  and (_09751_, _09750_, _22773_);
  and (_04088_, _09751_, _09746_);
  and (_09752_, _02829_, _23715_);
  and (_09753_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or (_27123_, _09753_, _09752_);
  and (_09754_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  and (_09755_, _09603_, _23715_);
  or (_04099_, _09755_, _09754_);
  and (_09756_, _05618_, _23247_);
  or (_09757_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_09758_, _05623_, _05616_);
  or (_09759_, _09758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand (_09760_, _05624_, _05616_);
  and (_09761_, _09760_, _09759_);
  or (_09762_, _09761_, _05656_);
  and (_09764_, _05659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_09765_, _09764_, _09762_);
  and (_09766_, _09765_, _09757_);
  and (_09767_, _09766_, _05619_);
  and (_09768_, _05617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_09769_, _09768_, _09767_);
  or (_09770_, _09769_, _09756_);
  and (_04101_, _09770_, _22773_);
  and (_09771_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_09772_, _09597_, _23983_);
  or (_04103_, _09772_, _09771_);
  and (_09773_, _24237_, _23924_);
  and (_09774_, _09773_, _23920_);
  not (_09775_, _09773_);
  and (_09776_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_04108_, _09776_, _09774_);
  and (_09778_, _09578_, _23930_);
  not (_09779_, _09778_);
  and (_09780_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_09782_, _09778_, _24053_);
  or (_26963_, _09782_, _09780_);
  and (_09783_, _09773_, _23715_);
  and (_09784_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or (_04112_, _09784_, _09783_);
  and (_09785_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_09786_, _09778_, _23693_);
  or (_04115_, _09786_, _09785_);
  and (_09787_, _09718_, _23983_);
  and (_09788_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_04119_, _09788_, _09787_);
  and (_09791_, _09773_, _24053_);
  and (_09792_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_04122_, _09792_, _09791_);
  and (_09793_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_09794_, _09778_, _23715_);
  or (_04126_, _09794_, _09793_);
  and (_09795_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_09796_, _09778_, _24027_);
  or (_04129_, _09796_, _09795_);
  or (_09797_, _05659_, _05656_);
  and (_09798_, _09797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_09799_, _05667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_09800_, _09799_, _05668_);
  and (_09801_, _09800_, _05674_);
  or (_09802_, _09801_, _05618_);
  or (_09803_, _09802_, _09798_);
  or (_09804_, _05682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_09805_, _09804_, _09803_);
  or (_09806_, _09805_, _05617_);
  nand (_09807_, _05617_, _24017_);
  and (_09809_, _09807_, _22773_);
  and (_04131_, _09809_, _09806_);
  and (_09810_, _08011_, _23693_);
  and (_09811_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or (_04132_, _09811_, _09810_);
  not (_09813_, _05713_);
  and (_09814_, _05705_, _24184_);
  or (_09815_, _09814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_09816_, _09815_, _09813_);
  nand (_09817_, _09814_, _23681_);
  and (_09818_, _09817_, _09816_);
  and (_09820_, _05713_, _23247_);
  or (_09821_, _09820_, _09818_);
  and (_04139_, _09821_, _22773_);
  and (_09822_, _09625_, _24053_);
  and (_09823_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  or (_04140_, _09823_, _09822_);
  and (_09824_, _09634_, _23920_);
  and (_09825_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  or (_04145_, _09825_, _09824_);
  and (_09827_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_09829_, _09778_, _23983_);
  or (_04148_, _09829_, _09827_);
  and (_09830_, _09578_, _23444_);
  not (_09831_, _09830_);
  and (_09832_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  and (_09833_, _09830_, _23751_);
  or (_26964_, _09833_, _09832_);
  and (_09835_, _09642_, _23983_);
  and (_09836_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_04153_, _09836_, _09835_);
  and (_09837_, _09642_, _24053_);
  and (_09838_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_27089_, _09838_, _09837_);
  and (_09839_, _09660_, _23920_);
  and (_09840_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_04157_, _09840_, _09839_);
  and (_09842_, _09676_, _23900_);
  and (_09843_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  or (_04161_, _09843_, _09842_);
  and (_09844_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and (_09845_, _09830_, _23693_);
  or (_04168_, _09845_, _09844_);
  and (_09847_, _09740_, _24027_);
  and (_09849_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or (_04181_, _09849_, _09847_);
  and (_09850_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  and (_09851_, _09830_, _23900_);
  or (_04184_, _09851_, _09850_);
  and (_09852_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  and (_09853_, _09830_, _24027_);
  or (_26966_, _09853_, _09852_);
  and (_09854_, _09740_, _24053_);
  and (_09855_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_27071_, _09855_, _09854_);
  and (_09856_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  and (_09857_, _09830_, _23983_);
  or (_04193_, _09857_, _09856_);
  and (_09858_, _08011_, _23920_);
  and (_09860_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or (_04199_, _09860_, _09858_);
  and (_09863_, _09625_, _23900_);
  and (_09865_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  or (_04212_, _09865_, _09863_);
  and (_09866_, _09578_, _23905_);
  not (_09867_, _09866_);
  and (_09868_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  and (_09869_, _09866_, _24053_);
  or (_04217_, _09869_, _09868_);
  and (_09870_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  and (_09871_, _09866_, _23715_);
  or (_04221_, _09871_, _09870_);
  and (_09872_, _07087_, _23920_);
  and (_09873_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_04226_, _09873_, _09872_);
  and (_09875_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  and (_09876_, _09866_, _23900_);
  or (_26967_, _09876_, _09875_);
  and (_09877_, _09732_, _23751_);
  and (_09878_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_04239_, _09878_, _09877_);
  nand (_09880_, _24192_, _23357_);
  nand (_09881_, _09685_, _09682_);
  and (_09882_, _09686_, _24975_);
  and (_09884_, _09882_, _09881_);
  or (_09886_, _09691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_09887_, _09692_);
  and (_09888_, _09887_, _24196_);
  and (_09889_, _09888_, _09886_);
  and (_09890_, _25012_, _24203_);
  and (_09891_, _09890_, _25000_);
  or (_09892_, _09891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_09893_, _09891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_09894_, _09893_, _25003_);
  and (_09896_, _09894_, _09892_);
  or (_09897_, _09896_, _09889_);
  or (_09898_, _09897_, _24192_);
  or (_09899_, _09898_, _09884_);
  and (_09900_, _09899_, _24188_);
  and (_09901_, _09900_, _09880_);
  and (_09903_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_09904_, _09903_, _09901_);
  and (_04241_, _09904_, _22773_);
  and (_09905_, _09773_, _23983_);
  and (_09906_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or (_04245_, _09906_, _09905_);
  and (_09907_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and (_09908_, _09866_, _24027_);
  or (_04248_, _09908_, _09907_);
  and (_09910_, _09578_, _24274_);
  not (_09912_, _09910_);
  and (_09913_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_09914_, _09910_, _23693_);
  or (_04276_, _09914_, _09913_);
  and (_09916_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_09918_, _09910_, _23900_);
  or (_04279_, _09918_, _09916_);
  and (_09921_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_09922_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_09924_, _23763_, _09922_);
  or (_09925_, _09924_, _09921_);
  and (_26854_[15], _09925_, _22773_);
  and (_09926_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_09927_, _09910_, _24027_);
  or (_26968_, _09927_, _09926_);
  and (_09929_, _06631_, _24027_);
  and (_09930_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or (_04290_, _09930_, _09929_);
  and (_09931_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  and (_09932_, _02842_, _23900_);
  or (_04294_, _09932_, _09931_);
  and (_09934_, _06631_, _23920_);
  and (_09936_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or (_04297_, _09936_, _09934_);
  and (_09937_, _09718_, _23920_);
  and (_09939_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_04299_, _09939_, _09937_);
  and (_09941_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_09942_, _09910_, _23983_);
  or (_04302_, _09942_, _09941_);
  and (_09944_, _09578_, _24145_);
  not (_09945_, _09944_);
  and (_09946_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_09947_, _09944_, _23751_);
  or (_04307_, _09947_, _09946_);
  and (_09948_, _09718_, _24027_);
  and (_09949_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_04309_, _09949_, _09948_);
  and (_09950_, _09773_, _23751_);
  and (_09952_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or (_04314_, _09952_, _09950_);
  and (_09953_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_09954_, _09944_, _23715_);
  or (_26969_, _09954_, _09953_);
  and (_09956_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_09957_, _02687_, _23751_);
  or (_27016_, _09957_, _09956_);
  and (_09959_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_09960_, _09944_, _23920_);
  or (_26970_, _09960_, _09959_);
  and (_09961_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_09963_, _09944_, _24027_);
  or (_26971_, _09963_, _09961_);
  and (_09965_, _09578_, _23924_);
  not (_09967_, _09965_);
  and (_09968_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  and (_09969_, _09965_, _23751_);
  or (_26973_, _09969_, _09968_);
  and (_09971_, _02688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_09972_, _02687_, _23920_);
  or (_27017_, _09972_, _09971_);
  and (_09973_, _09773_, _23693_);
  and (_09975_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or (_27085_, _09975_, _09973_);
  or (_09976_, _07311_, _23205_);
  and (_09977_, _24984_, _24202_);
  and (_09978_, _09977_, _25011_);
  or (_09980_, _09978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_09981_, _09890_);
  and (_09982_, _09981_, _25002_);
  and (_09983_, _09982_, _09980_);
  and (_09984_, _09977_, _25007_);
  nand (_09985_, _09984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_09986_, _09984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_09987_, _09986_, _24975_);
  and (_09988_, _09987_, _09985_);
  nand (_09989_, _09691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_09990_, _24202_, _24193_);
  and (_09991_, _09990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_09992_, _09991_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_09994_, _09992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_09995_, _09994_, _09989_);
  or (_09996_, _09995_, _09988_);
  or (_09997_, _09996_, _09983_);
  or (_09998_, _09997_, _24192_);
  and (_09999_, _09998_, _24188_);
  and (_10000_, _09999_, _09976_);
  and (_10001_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_10002_, _10001_, _10000_);
  and (_04357_, _10002_, _22773_);
  and (_10003_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and (_10004_, _09965_, _23693_);
  or (_26974_, _10004_, _10003_);
  and (_10005_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  and (_10006_, _09965_, _23900_);
  or (_26975_, _10006_, _10005_);
  and (_10007_, _09773_, _23900_);
  and (_10008_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or (_27086_, _10008_, _10007_);
  and (_10009_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  and (_10010_, _09965_, _24027_);
  or (_26976_, _10010_, _10009_);
  and (_10012_, _09773_, _24027_);
  and (_10013_, _09775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or (_27087_, _10013_, _10012_);
  and (_10015_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and (_10017_, _24275_, _23715_);
  or (_27019_, _10017_, _10015_);
  and (_10018_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and (_10019_, _24275_, _23693_);
  or (_27018_, _10019_, _10018_);
  and (_10020_, _04141_, _24027_);
  and (_10022_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or (_27069_, _10022_, _10020_);
  and (_10024_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_10025_, _02499_, _23751_);
  or (_26984_, _10025_, _10024_);
  and (_10026_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and (_10028_, _02662_, _23751_);
  or (_26981_, _10028_, _10026_);
  and (_10030_, _04141_, _23983_);
  and (_10031_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or (_27070_, _10031_, _10030_);
  and (_10032_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  and (_10033_, _02662_, _23693_);
  or (_26982_, _10033_, _10032_);
  and (_10035_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_10036_, _02499_, _23715_);
  or (_26985_, _10036_, _10035_);
  and (_10038_, _09740_, _23751_);
  and (_10040_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or (_27072_, _10040_, _10038_);
  and (_10042_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and (_10043_, _02662_, _23900_);
  or (_26983_, _10043_, _10042_);
  and (_10044_, _09740_, _23693_);
  and (_10045_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or (_27073_, _10045_, _10044_);
  and (_10046_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_10047_, _02409_, _23920_);
  or (_26990_, _10047_, _10046_);
  and (_10049_, _02410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_10051_, _02409_, _23715_);
  or (_26989_, _10051_, _10049_);
  and (_10052_, _09740_, _23715_);
  and (_10053_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or (_27074_, _10053_, _10052_);
  and (_10054_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and (_10055_, _02362_, _24053_);
  or (_26992_, _10055_, _10054_);
  and (_10057_, _09740_, _23920_);
  and (_10058_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_27075_, _10058_, _10057_);
  and (_10059_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_10060_, _09579_, _23715_);
  or (_26955_, _10060_, _10059_);
  and (_10061_, _02363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and (_10062_, _02362_, _23983_);
  or (_26994_, _10062_, _10061_);
  and (_10064_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_10065_, _09579_, _23693_);
  or (_26954_, _10065_, _10064_);
  and (_10067_, _09740_, _23983_);
  and (_10069_, _09742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or (_27076_, _10069_, _10067_);
  and (_10070_, _09732_, _24053_);
  and (_10071_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_27077_, _10071_, _10070_);
  and (_10074_, _02171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  and (_10075_, _02170_, _23920_);
  or (_26995_, _10075_, _10074_);
  and (_10077_, _09732_, _23693_);
  and (_10078_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_27078_, _10078_, _10077_);
  and (_10079_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_10080_, _01768_, _23693_);
  or (_26996_, _10080_, _10079_);
  and (_10081_, _09732_, _23715_);
  and (_10083_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_27079_, _10083_, _10081_);
  and (_10084_, _01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_10085_, _01768_, _24027_);
  or (_26999_, _10085_, _10084_);
  and (_10086_, _25491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_10088_, _25490_, _23900_);
  or (_27001_, _10088_, _10086_);
  and (_10090_, _09578_, _24097_);
  not (_10092_, _10090_);
  and (_10094_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_10096_, _10090_, _23900_);
  or (_26953_, _10096_, _10094_);
  and (_10099_, _09732_, _23920_);
  and (_10101_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_27080_, _10101_, _10099_);
  and (_10102_, _07484_, _24053_);
  and (_10103_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_27218_, _10103_, _10102_);
  and (_10106_, _09732_, _23983_);
  and (_10107_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_27082_, _10107_, _10106_);
  and (_10108_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_10109_, _10090_, _23715_);
  or (_04522_, _10109_, _10108_);
  and (_10110_, _09718_, _24053_);
  and (_10111_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_27083_, _10111_, _10110_);
  and (_10112_, _01927_, _23693_);
  and (_10113_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_04531_, _10113_, _10112_);
  and (_10115_, _09718_, _23751_);
  and (_10117_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_04540_, _10117_, _10115_);
  and (_10118_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_10120_, _10090_, _23693_);
  or (_04552_, _10120_, _10118_);
  and (_10122_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_10123_, _25153_, _23900_);
  or (_04559_, _10123_, _10122_);
  and (_10125_, _09718_, _23693_);
  and (_10127_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_04562_, _10127_, _10125_);
  and (_10128_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  and (_10129_, _24393_, _23900_);
  or (_04567_, _10129_, _10128_);
  and (_10130_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  and (_10131_, _24393_, _23751_);
  or (_04575_, _10131_, _10130_);
  and (_10132_, _24796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and (_10134_, _24795_, _23693_);
  or (_04580_, _10134_, _10132_);
  and (_10136_, _09718_, _23715_);
  and (_10137_, _09720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_27084_, _10137_, _10136_);
  and (_10138_, _24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and (_10139_, _24393_, _23983_);
  or (_04584_, _10139_, _10138_);
  and (_10140_, _24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  and (_10141_, _24275_, _23983_);
  or (_27021_, _10141_, _10140_);
  and (_10144_, _09676_, _24053_);
  and (_10145_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  or (_04597_, _10145_, _10144_);
  and (_10148_, _25364_, _23751_);
  and (_10150_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or (_04603_, _10150_, _10148_);
  and (_10152_, _24147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and (_10153_, _24146_, _23715_);
  or (_04613_, _10153_, _10152_);
  and (_10154_, _09676_, _23751_);
  and (_10155_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  or (_04620_, _10155_, _10154_);
  and (_10158_, _09676_, _23715_);
  and (_10160_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  or (_04626_, _10160_, _10158_);
  and (_10162_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_10164_, _10090_, _24027_);
  or (_04633_, _10164_, _10162_);
  and (_10166_, _09676_, _23920_);
  and (_10168_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  or (_04638_, _10168_, _10166_);
  and (_10170_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_10171_, _10090_, _23920_);
  or (_04659_, _10171_, _10170_);
  and (_10172_, _23939_, _23715_);
  and (_10173_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or (_27026_, _10173_, _10172_);
  and (_10175_, _09676_, _24027_);
  and (_10176_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  or (_04664_, _10176_, _10175_);
  and (_10177_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  and (_10178_, _02842_, _23715_);
  or (_27138_, _10178_, _10177_);
  and (_10180_, _09676_, _23983_);
  and (_10181_, _09678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  or (_04675_, _10181_, _10180_);
  or (_10183_, _23413_, _23253_);
  and (_10184_, _23270_, _23268_);
  nor (_10186_, _10184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_10187_, _10184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_10188_, _10187_, _10186_);
  nor (_10189_, _25045_, _23210_);
  and (_10190_, _10189_, _10188_);
  not (_10191_, _10189_);
  and (_10192_, _10191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_10193_, _24294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_10195_, _10193_, _23210_);
  or (_10196_, _10195_, _10192_);
  or (_10198_, _10196_, _10190_);
  or (_10199_, _10198_, _23252_);
  and (_10200_, _10199_, _22773_);
  and (_04679_, _10200_, _10183_);
  and (_10203_, _10189_, _23268_);
  nand (_10204_, _24284_, _23360_);
  or (_10205_, _10204_, _23210_);
  and (_10206_, _10205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_10207_, _10206_, _10203_);
  or (_10208_, _10203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_10209_, _10208_, _10207_);
  or (_10210_, _10209_, _23252_);
  nand (_10211_, _24047_, _23252_);
  and (_10213_, _10211_, _22773_);
  and (_04685_, _10213_, _10210_);
  and (_10214_, _09660_, _24053_);
  and (_10215_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_04687_, _10215_, _10214_);
  and (_10218_, _23272_, _23268_);
  and (_10219_, _10218_, _23373_);
  nor (_10220_, _10219_, _23277_);
  and (_10221_, _10220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_10222_, _10220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_10223_, _10222_, _10221_);
  nor (_10224_, _10223_, _23210_);
  and (_10225_, _24788_, _23210_);
  or (_10226_, _10225_, _23252_);
  or (_10227_, _10226_, _10224_);
  or (_10229_, _23253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_10230_, _10229_, _22773_);
  and (_04690_, _10230_, _10227_);
  and (_10233_, _01759_, _23920_);
  and (_10235_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or (_04693_, _10235_, _10233_);
  and (_10237_, _01701_, _24053_);
  and (_10238_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or (_04696_, _10238_, _10237_);
  and (_10239_, _09660_, _23693_);
  and (_10240_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_04701_, _10240_, _10239_);
  and (_10241_, _09660_, _23900_);
  and (_10242_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_04703_, _10242_, _10241_);
  or (_10243_, _07311_, _23413_);
  and (_10244_, _25012_, _24201_);
  and (_10245_, _10244_, _25000_);
  or (_10246_, _10245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_10247_, _10245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_10248_, _10247_, _25003_);
  and (_10249_, _10248_, _10246_);
  and (_10250_, _24201_, _24193_);
  or (_10251_, _10250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_10252_, _09990_);
  and (_10253_, _10252_, _24196_);
  and (_10255_, _10253_, _10251_);
  and (_10257_, _24989_, _24201_);
  or (_10259_, _10257_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_10260_, _09684_, _24975_);
  and (_10261_, _10260_, _10259_);
  or (_10263_, _10261_, _10255_);
  or (_10265_, _10263_, _10249_);
  or (_10267_, _10265_, _24192_);
  and (_10268_, _10267_, _24188_);
  and (_10270_, _10268_, _10243_);
  and (_10271_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_10272_, _10271_, _10270_);
  and (_04706_, _10272_, _22773_);
  and (_10273_, _23938_, _23891_);
  and (_10274_, _10273_, _23983_);
  not (_10275_, _10273_);
  and (_10276_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  or (_04713_, _10276_, _10274_);
  or (_10277_, _24188_, _23413_);
  or (_10278_, _07311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_10279_, _25011_, _25001_);
  and (_10280_, _10279_, _24984_);
  and (_10282_, _10280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_10283_, _24987_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  not (_10285_, _24988_);
  or (_10286_, _10285_, _24192_);
  and (_10288_, _10286_, _10283_);
  or (_10290_, _10288_, _10282_);
  and (_10291_, _10290_, _10278_);
  or (_10292_, _10291_, _24186_);
  and (_10293_, _10292_, _22773_);
  and (_04716_, _10293_, _10277_);
  and (_10294_, _09660_, _24027_);
  and (_10295_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_27088_, _10295_, _10294_);
  and (_10298_, _02403_, _24027_);
  and (_10300_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_04720_, _10300_, _10298_);
  and (_10303_, _09578_, _24068_);
  not (_10304_, _10303_);
  and (_10305_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  and (_10306_, _10303_, _24027_);
  or (_04723_, _10306_, _10305_);
  or (_10307_, _07311_, _23247_);
  and (_10308_, _07314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_10309_, _10308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  not (_10310_, _10244_);
  and (_10311_, _10310_, _25002_);
  and (_10312_, _10311_, _10309_);
  nand (_10314_, _07328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_10315_, _07328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_10316_, _10315_, _10314_);
  and (_10317_, _10316_, _24975_);
  nand (_10318_, _10250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_10319_, _07322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_10320_, _10319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_10322_, _10320_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_10323_, _10322_, _10318_);
  or (_10324_, _10323_, _10317_);
  or (_10326_, _10324_, _10312_);
  or (_10327_, _10326_, _24192_);
  and (_10328_, _10327_, _24188_);
  and (_10329_, _10328_, _10307_);
  and (_10330_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_10331_, _10330_, _10329_);
  and (_04726_, _10331_, _22773_);
  or (_10333_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_10334_, _10333_, _22773_);
  or (_10335_, _23247_, _22931_);
  and (_04729_, _10335_, _10334_);
  and (_10337_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and (_10338_, _10303_, _23920_);
  or (_04732_, _10338_, _10337_);
  and (_10341_, _25164_, _24274_);
  and (_10342_, _10341_, _24053_);
  not (_10343_, _10341_);
  and (_10345_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_04737_, _10345_, _10342_);
  and (_10347_, _09660_, _23983_);
  and (_10349_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_04739_, _10349_, _10347_);
  and (_10351_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and (_10352_, _10303_, _23900_);
  or (_04743_, _10352_, _10351_);
  and (_10353_, _01908_, _23920_);
  and (_10354_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or (_27032_, _10354_, _10353_);
  and (_10356_, _09642_, _23751_);
  and (_10358_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_04764_, _10358_, _10356_);
  and (_10360_, _09642_, _23715_);
  and (_10361_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_27090_, _10361_, _10360_);
  and (_10363_, _02509_, _23983_);
  and (_10364_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_27034_, _10364_, _10363_);
  and (_10365_, _09642_, _23900_);
  and (_10367_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_04776_, _10367_, _10365_);
  and (_10370_, _09642_, _24027_);
  and (_10372_, _09644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_04780_, _10372_, _10370_);
  and (_10375_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  and (_10376_, _02718_, _23920_);
  or (_04781_, _10376_, _10375_);
  and (_10378_, _02248_, _23900_);
  and (_10379_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or (_04784_, _10379_, _10378_);
  and (_10381_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  and (_10382_, _02718_, _23900_);
  or (_04789_, _10382_, _10381_);
  and (_10383_, _02248_, _23693_);
  and (_10384_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or (_04791_, _10384_, _10383_);
  and (_10385_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_10387_, _10090_, _24053_);
  or (_04798_, _10387_, _10385_);
  and (_10390_, _25364_, _23715_);
  and (_10392_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or (_04804_, _10392_, _10390_);
  and (_10395_, _25364_, _24053_);
  and (_10396_, _25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or (_27035_, _10396_, _10395_);
  and (_10398_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  and (_10399_, _02718_, _23715_);
  or (_04810_, _10399_, _10398_);
  and (_10400_, _09634_, _23751_);
  and (_10402_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  or (_27092_, _10402_, _10400_);
  and (_10403_, _09634_, _23693_);
  and (_10404_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  or (_04831_, _10404_, _10403_);
  and (_10405_, _09634_, _23900_);
  and (_10407_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  or (_27093_, _10407_, _10405_);
  and (_10409_, _09634_, _24027_);
  and (_10410_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  or (_04855_, _10410_, _10409_);
  and (_10411_, _24274_, _23719_);
  and (_10412_, _10411_, _23900_);
  not (_10413_, _10411_);
  and (_10414_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or (_04862_, _10414_, _10412_);
  and (_10415_, _09634_, _23983_);
  and (_10416_, _09636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  or (_04878_, _10416_, _10415_);
  and (_10417_, _10411_, _23983_);
  and (_10418_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or (_04882_, _10418_, _10417_);
  and (_10420_, _09625_, _23751_);
  and (_10421_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  or (_04885_, _10421_, _10420_);
  and (_10422_, _09625_, _23693_);
  and (_10424_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  or (_04894_, _10424_, _10422_);
  and (_10425_, _09625_, _23920_);
  and (_10426_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or (_04898_, _10426_, _10425_);
  and (_10427_, _24901_, _24027_);
  and (_10428_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_04903_, _10428_, _10427_);
  and (_10429_, _24901_, _23715_);
  and (_10430_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_04907_, _10430_, _10429_);
  and (_10431_, _09578_, _23700_);
  not (_10432_, _10431_);
  and (_10433_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and (_10434_, _10431_, _23983_);
  or (_26950_, _10434_, _10433_);
  and (_10436_, _24268_, _23900_);
  and (_10437_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or (_04909_, _10437_, _10436_);
  and (_10439_, _09625_, _24027_);
  and (_10440_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  or (_27094_, _10440_, _10439_);
  and (_10441_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  and (_10442_, _02718_, _23983_);
  or (_04910_, _10442_, _10441_);
  and (_10443_, _02719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  and (_10444_, _02718_, _24027_);
  or (_04930_, _10444_, _10443_);
  and (_10445_, _09625_, _23983_);
  and (_10446_, _09627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or (_04933_, _10446_, _10445_);
  and (_10447_, _24268_, _24027_);
  and (_10448_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or (_04936_, _10448_, _10447_);
  and (_10449_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and (_10450_, _10303_, _23751_);
  or (_04946_, _10450_, _10449_);
  and (_10452_, _08011_, _24027_);
  and (_10453_, _08013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or (_04956_, _10453_, _10452_);
  and (_10454_, _09608_, _24053_);
  and (_10455_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_04958_, _10455_, _10454_);
  and (_10456_, _24305_, _23920_);
  and (_10457_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_27049_, _10457_, _10456_);
  and (_10458_, _09608_, _23693_);
  and (_10459_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_27095_, _10459_, _10458_);
  and (_10461_, _09570_, _23715_);
  and (_10462_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_27053_, _10462_, _10461_);
  and (_10463_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and (_10464_, _10303_, _23693_);
  or (_04972_, _10464_, _10463_);
  and (_10466_, _05883_, _23751_);
  and (_10469_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_04974_, _10469_, _10466_);
  and (_10470_, _08005_, _24053_);
  and (_10471_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_04976_, _10471_, _10470_);
  and (_10472_, _09608_, _23715_);
  and (_10473_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_04978_, _10473_, _10472_);
  and (_10474_, _09608_, _23920_);
  and (_10475_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_04980_, _10475_, _10474_);
  and (_10476_, _24098_, _23715_);
  and (_10477_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or (_04984_, _10477_, _10476_);
  and (_10478_, _24238_, _24053_);
  and (_10479_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or (_04987_, _10479_, _10478_);
  and (_10480_, _09463_, _24027_);
  and (_10481_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_04990_, _10481_, _10480_);
  and (_10482_, _24238_, _24027_);
  and (_10483_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or (_27058_, _10483_, _10482_);
  and (_10485_, _09608_, _24027_);
  and (_10487_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_04997_, _10487_, _10485_);
  and (_10488_, _24238_, _23715_);
  and (_10489_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or (_27057_, _10489_, _10488_);
  and (_10490_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_10491_, _02722_, _23920_);
  or (_05000_, _10491_, _10490_);
  and (_10494_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_10495_, _02722_, _23900_);
  or (_05004_, _10495_, _10494_);
  and (_10496_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  and (_10497_, _10431_, _23693_);
  or (_05060_, _10497_, _10496_);
  and (_10498_, _05883_, _24053_);
  and (_10499_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_05066_, _10499_, _10498_);
  and (_10500_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  and (_10501_, _10431_, _23751_);
  or (_05078_, _10501_, _10500_);
  and (_10502_, _08005_, _23751_);
  and (_10503_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_05095_, _10503_, _10502_);
  and (_10504_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  and (_10505_, _10431_, _24053_);
  or (_05106_, _10505_, _10504_);
  and (_10507_, _08005_, _23900_);
  and (_10509_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_05121_, _10509_, _10507_);
  and (_10510_, _08005_, _24027_);
  and (_10511_, _08007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_05147_, _10511_, _10510_);
  and (_10512_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  and (_10513_, _10431_, _23900_);
  or (_05152_, _10513_, _10512_);
  and (_10514_, _25164_, _23924_);
  and (_10515_, _10514_, _23983_);
  not (_10516_, _10514_);
  and (_10517_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_05158_, _10517_, _10515_);
  and (_10519_, _10514_, _24027_);
  and (_10520_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_26980_, _10520_, _10519_);
  and (_10521_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_10522_, _02722_, _23983_);
  or (_05171_, _10522_, _10521_);
  and (_10523_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  and (_10524_, _10431_, _23920_);
  or (_05175_, _10524_, _10523_);
  and (_10525_, _23930_, _23891_);
  and (_10526_, _10525_, _23920_);
  not (_10527_, _10525_);
  and (_10528_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or (_05192_, _10528_, _10526_);
  and (_10531_, _07999_, _23751_);
  and (_10532_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_05195_, _10532_, _10531_);
  and (_10533_, _10525_, _23983_);
  and (_10534_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or (_05200_, _10534_, _10533_);
  and (_10536_, _24388_, _24097_);
  and (_10537_, _10536_, _23751_);
  not (_10538_, _10536_);
  and (_10539_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or (_05203_, _10539_, _10537_);
  and (_10541_, _10525_, _24027_);
  and (_10542_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or (_05211_, _10542_, _10541_);
  and (_10543_, _01936_, _23983_);
  and (_10544_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_05216_, _10544_, _10543_);
  and (_10545_, _10536_, _24053_);
  and (_10546_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or (_05237_, _10546_, _10545_);
  and (_10547_, _24388_, _23938_);
  and (_10548_, _10547_, _23751_);
  not (_10549_, _10547_);
  and (_10550_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or (_05244_, _10550_, _10548_);
  and (_10551_, _07999_, _23715_);
  and (_10552_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_27119_, _10552_, _10551_);
  and (_10553_, _10547_, _24053_);
  and (_10554_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or (_27008_, _10554_, _10553_);
  and (_10556_, _07999_, _23920_);
  and (_10558_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_05256_, _10558_, _10556_);
  and (_10561_, _09480_, _23920_);
  and (_10562_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or (_05259_, _10562_, _10561_);
  and (_10563_, _09578_, _23938_);
  not (_10564_, _10563_);
  and (_10565_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_10566_, _10563_, _23900_);
  or (_05268_, _10566_, _10565_);
  and (_10567_, _07999_, _23983_);
  and (_10568_, _08001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_05272_, _10568_, _10567_);
  and (_10569_, _25176_, _24053_);
  and (_10570_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or (_05279_, _10570_, _10569_);
  and (_10573_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_10574_, _10563_, _23715_);
  or (_05284_, _10574_, _10573_);
  and (_10575_, _09480_, _23900_);
  and (_10576_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or (_05290_, _10576_, _10575_);
  and (_10577_, _01932_, _23751_);
  and (_10579_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_05292_, _10579_, _10577_);
  and (_10580_, _10514_, _24053_);
  and (_10581_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_05297_, _10581_, _10580_);
  and (_10583_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_10584_, _10563_, _23693_);
  or (_05299_, _10584_, _10583_);
  and (_10585_, _09552_, _23751_);
  and (_10586_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_05302_, _10586_, _10585_);
  and (_10588_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_10590_, _02722_, _24053_);
  or (_05305_, _10590_, _10588_);
  and (_10591_, _09552_, _24053_);
  and (_10592_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_05331_, _10592_, _10591_);
  and (_10594_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_10595_, _02726_, _23983_);
  or (_05333_, _10595_, _10594_);
  and (_10597_, _10514_, _23693_);
  and (_10598_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_26978_, _10598_, _10597_);
  and (_10599_, _10514_, _23900_);
  and (_10600_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_05342_, _10600_, _10599_);
  and (_10601_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_10602_, _10563_, _23983_);
  or (_05348_, _10602_, _10601_);
  and (_10603_, _10514_, _23715_);
  and (_10604_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_26979_, _10604_, _10603_);
  and (_10605_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_10606_, _10563_, _24027_);
  or (_05353_, _10606_, _10605_);
  and (_10609_, _04091_, _23693_);
  and (_10610_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  or (_05360_, _10610_, _10609_);
  and (_10611_, _24238_, _23920_);
  and (_10612_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_05366_, _10612_, _10611_);
  and (_10615_, _04077_, _24027_);
  and (_10616_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or (_05370_, _10616_, _10615_);
  and (_10617_, _04095_, _23715_);
  and (_10619_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_05373_, _10619_, _10617_);
  and (_10620_, _04077_, _23693_);
  and (_10622_, _04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or (_05378_, _10622_, _10620_);
  and (_10624_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_10625_, _10563_, _23920_);
  or (_05379_, _10625_, _10624_);
  and (_10628_, _04073_, _23900_);
  and (_10629_, _04075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_05382_, _10629_, _10628_);
  and (_10631_, _24069_, _23900_);
  and (_10632_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or (_27195_, _10632_, _10631_);
  and (_10634_, _24238_, _23900_);
  and (_10636_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or (_05386_, _10636_, _10634_);
  and (_10637_, _02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_10639_, _02722_, _23693_);
  or (_05389_, _10639_, _10637_);
  and (_10641_, _04095_, _23900_);
  and (_10642_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_27097_, _10642_, _10641_);
  and (_10643_, _10536_, _23920_);
  and (_10644_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or (_05420_, _10644_, _10643_);
  and (_10646_, _10536_, _23693_);
  and (_10647_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or (_05427_, _10647_, _10646_);
  and (_10648_, _06631_, _23693_);
  and (_10649_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or (_05438_, _10649_, _10648_);
  and (_10650_, _10536_, _23715_);
  and (_10651_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or (_05440_, _10651_, _10650_);
  and (_10652_, _24164_, _24053_);
  and (_10654_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_05446_, _10654_, _10652_);
  and (_10655_, _04200_, _24027_);
  and (_10656_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_05461_, _10656_, _10655_);
  and (_10657_, _04095_, _23983_);
  and (_10658_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_05465_, _10658_, _10657_);
  or (_10661_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_10662_, _25591_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_10663_, _10662_, _22773_);
  and (_26875_[31], _10663_, _10661_);
  and (_10666_, _04091_, _24053_);
  and (_10667_, _04093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  or (_05469_, _10667_, _10666_);
  and (_10669_, _23986_, _24083_);
  and (_10670_, _10669_, _23924_);
  not (_10671_, _10670_);
  and (_10672_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_10673_, _10670_, _23919_);
  or (_26949_, _10673_, _10672_);
  and (_10674_, _25198_, _24053_);
  and (_10675_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or (_05472_, _10675_, _10674_);
  and (_10677_, _10536_, _24027_);
  and (_10678_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or (_05476_, _10678_, _10677_);
  and (_10681_, _10536_, _23983_);
  and (_10682_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or (_05483_, _10682_, _10681_);
  and (_05488_, _26508_, _22773_);
  and (_05490_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _22773_);
  and (_05493_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _22773_);
  and (_05495_, _26601_, _22773_);
  and (_10683_, _04095_, _24027_);
  and (_10684_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_05497_, _10684_, _10683_);
  and (_05503_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _22773_);
  and (_10685_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_10687_, _10670_, _23899_);
  or (_26948_, _10687_, _10685_);
  and (_10689_, _02423_, _23693_);
  and (_10690_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or (_05506_, _10690_, _10689_);
  and (_10692_, _04200_, _23693_);
  and (_10693_, _04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_27065_, _10693_, _10692_);
  and (_10695_, _24388_, _23700_);
  and (_10697_, _10695_, _23983_);
  not (_10698_, _10695_);
  and (_10699_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_05520_, _10699_, _10697_);
  and (_10702_, _04141_, _23900_);
  and (_10703_, _04143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or (_05522_, _10703_, _10702_);
  and (_10705_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_10706_, _10670_, _23714_);
  or (_05525_, _10706_, _10705_);
  and (_10708_, _10695_, _24027_);
  and (_10709_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_05528_, _10709_, _10708_);
  or (_10710_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_10711_, _04915_, rst);
  and (_05531_, _10711_, _10710_);
  nand (_10713_, _23976_, _23210_);
  not (_10714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_10716_, _23360_, _23268_);
  and (_10717_, _10716_, _23257_);
  not (_10718_, _25037_);
  and (_10719_, _23281_, _23279_);
  nor (_10720_, _10719_, _23257_);
  nor (_10721_, _10720_, _10718_);
  not (_10722_, _10721_);
  nor (_10723_, _10722_, _10717_);
  and (_10724_, _10723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_10726_, _10724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_10727_, _10726_, _10714_);
  and (_10728_, _10726_, _10714_);
  or (_10729_, _10728_, _10727_);
  or (_10730_, _10729_, _23210_);
  and (_10731_, _10730_, _23253_);
  and (_10733_, _10731_, _10713_);
  and (_10734_, _23252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_10736_, _10734_, _10733_);
  and (_05533_, _10736_, _22773_);
  and (_10738_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_10740_, _02726_, _23715_);
  or (_05539_, _10740_, _10738_);
  and (_05542_, _00060_, _22773_);
  and (_05545_, _00149_, _22773_);
  and (_05548_, _26605_, _22773_);
  and (_10742_, _24164_, _23900_);
  and (_10743_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_05551_, _10743_, _10742_);
  and (_10745_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_10746_, _10563_, _24053_);
  or (_05554_, _10746_, _10745_);
  and (_05558_, _00327_, _22773_);
  and (_10747_, _01936_, _23693_);
  and (_10749_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_05560_, _10749_, _10747_);
  and (_05562_, _00406_, _22773_);
  and (_05565_, _00235_, _22773_);
  and (_10751_, _10525_, _24053_);
  and (_10752_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or (_05568_, _10752_, _10751_);
  and (_05572_, _00527_, _22773_);
  and (_10754_, _01936_, _23751_);
  and (_10755_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_27040_, _10755_, _10754_);
  and (_10756_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  nor (_10757_, _10671_, _23982_);
  or (_05574_, _10757_, _10756_);
  and (_10758_, _24740_, _23693_);
  and (_10759_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_05581_, _10759_, _10758_);
  and (_10760_, _01936_, _24053_);
  and (_10761_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_05583_, _10761_, _10760_);
  and (_10764_, _25524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_10765_, _25591_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_10766_, _10765_, _10764_);
  and (_26874_[31], _10766_, _22773_);
  and (_10768_, _04095_, _23693_);
  and (_10770_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_05600_, _10770_, _10768_);
  and (_10771_, _08402_, _23983_);
  and (_10772_, _08405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_05603_, _10772_, _10771_);
  and (_10774_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_10775_, _02726_, _23693_);
  or (_05608_, _10775_, _10774_);
  and (_10776_, _04095_, _24053_);
  and (_10777_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_05612_, _10777_, _10776_);
  and (_10779_, _02350_, _24053_);
  and (_10780_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_05614_, _10780_, _10779_);
  and (_10781_, _04095_, _23751_);
  and (_10782_, _04097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_27096_, _10782_, _10781_);
  and (_10784_, _24740_, _23751_);
  and (_10785_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_26915_, _10785_, _10784_);
  and (_10787_, _10695_, _24053_);
  and (_10788_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_27028_, _10788_, _10787_);
  and (_10790_, _10547_, _23983_);
  and (_10792_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or (_05638_, _10792_, _10790_);
  and (_10793_, _24164_, _23751_);
  and (_10795_, _24166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_05640_, _10795_, _10793_);
  and (_10796_, _10547_, _24027_);
  and (_10797_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or (_05642_, _10797_, _10796_);
  and (_10799_, _10669_, _24145_);
  not (_10801_, _10799_);
  and (_10802_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  nor (_10803_, _10801_, _24026_);
  or (_05649_, _10803_, _10802_);
  and (_10805_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  and (_10807_, _10799_, _23919_);
  or (_05654_, _10807_, _10805_);
  or (_10808_, _01583_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_26873_[3], _10808_, _22773_);
  not (_10809_, _01577_);
  and (_10811_, _01580_, _10809_);
  and (_10812_, _26873_[3], _01586_);
  and (_26872_, _10812_, _10811_);
  and (_10813_, _10695_, _23693_);
  and (_10814_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_05666_, _10814_, _10813_);
  and (_10815_, _10695_, _23900_);
  and (_10817_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_27030_, _10817_, _10815_);
  and (_10819_, _10695_, _23715_);
  and (_10820_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_05669_, _10820_, _10819_);
  and (_10821_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_10822_, _02726_, _23920_);
  or (_05690_, _10822_, _10821_);
  and (_10823_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and (_10824_, _02662_, _23715_);
  or (_05695_, _10824_, _10823_);
  and (_10825_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and (_10827_, _02662_, _24053_);
  or (_05701_, _10827_, _10825_);
  and (_10828_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_10829_, _02726_, _23900_);
  or (_05703_, _10829_, _10828_);
  and (_10830_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  and (_10831_, _09965_, _23920_);
  or (_05707_, _10831_, _10830_);
  and (_10833_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  and (_10834_, _09965_, _23715_);
  or (_05712_, _10834_, _10833_);
  or (_10836_, _24188_, _23247_);
  nor (_10837_, _24986_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_10838_, _10837_, _24987_);
  and (_10840_, _10280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_10841_, _10840_, _10838_);
  nor (_10842_, _10841_, _24192_);
  and (_10843_, _24192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_10844_, _10843_, _10842_);
  or (_10846_, _10844_, _24186_);
  and (_10847_, _10846_, _22773_);
  and (_05715_, _10847_, _10836_);
  and (_10848_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and (_10849_, _10670_, _23750_);
  or (_05717_, _10849_, _10848_);
  and (_10850_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_10851_, _10670_, _24052_);
  or (_26947_, _10851_, _10850_);
  and (_10852_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_10853_, _09944_, _23983_);
  or (_05722_, _10853_, _10852_);
  and (_10856_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_10857_, _09944_, _23693_);
  or (_05729_, _10857_, _10856_);
  and (_10859_, _10547_, _23920_);
  and (_10860_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or (_27010_, _10860_, _10859_);
  and (_10862_, _10547_, _23900_);
  and (_10864_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or (_05735_, _10864_, _10862_);
  and (_10865_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_10866_, _09910_, _23715_);
  or (_05750_, _10866_, _10865_);
  and (_10868_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_10869_, _09910_, _24053_);
  or (_05753_, _10869_, _10868_);
  and (_10871_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and (_10872_, _09866_, _23983_);
  or (_05757_, _10872_, _10871_);
  and (_10874_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  and (_10876_, _09866_, _23920_);
  or (_05760_, _10876_, _10874_);
  nor (_10877_, _24985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_10879_, _10877_, _24986_);
  and (_10880_, _10280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_10881_, _10880_, _10879_);
  nor (_10882_, _10881_, _24192_);
  and (_10883_, _24192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_10884_, _10883_, _10882_);
  and (_10886_, _10884_, _24188_);
  and (_10887_, _24186_, _23744_);
  or (_10888_, _10887_, _10886_);
  and (_05762_, _10888_, _22773_);
  and (_10889_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and (_10891_, _09866_, _23751_);
  or (_05764_, _10891_, _10889_);
  and (_10892_, _02843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  and (_10894_, _02842_, _24053_);
  or (_05767_, _10894_, _10892_);
  and (_10896_, _10341_, _23715_);
  and (_10897_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_26943_, _10897_, _10896_);
  and (_10899_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  and (_10900_, _09830_, _23920_);
  or (_26965_, _10900_, _10899_);
  and (_10901_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  and (_10902_, _09830_, _23715_);
  or (_05774_, _10902_, _10901_);
  and (_10904_, _10341_, _23693_);
  and (_10905_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_05777_, _10905_, _10904_);
  and (_10906_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  and (_10907_, _03157_, _23920_);
  or (_05789_, _10907_, _10906_);
  nor (_10908_, _24984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_10909_, _10908_, _24985_);
  and (_10910_, _07313_, _10279_);
  or (_10911_, _10910_, _10909_);
  or (_10913_, _10911_, _24192_);
  or (_10914_, _07311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_10915_, _10914_, _10913_);
  or (_10916_, _10915_, _24186_);
  nand (_10918_, _24186_, _24047_);
  and (_10919_, _10918_, _22773_);
  and (_05792_, _10919_, _10916_);
  and (_10920_, _10341_, _23751_);
  and (_10921_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_05794_, _10921_, _10920_);
  and (_10922_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_10923_, _09778_, _23900_);
  or (_05800_, _10923_, _10922_);
  not (_10926_, _04868_);
  not (_10928_, _04832_);
  and (_10930_, _04823_, _04821_);
  and (_10931_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and (_10932_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_10933_, _10932_, _10931_);
  and (_10934_, _10933_, _10928_);
  and (_10936_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_10937_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_10939_, _10937_, _10936_);
  and (_10940_, _10939_, _04832_);
  or (_10942_, _10940_, _10934_);
  or (_10943_, _10942_, _10926_);
  not (_10945_, _04859_);
  and (_10946_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and (_10948_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_10950_, _10948_, _10946_);
  and (_10952_, _10950_, _10928_);
  and (_10953_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_10955_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_10957_, _10955_, _10953_);
  and (_10958_, _10957_, _04832_);
  or (_10959_, _10958_, _10952_);
  or (_10961_, _10959_, _04868_);
  and (_10962_, _10961_, _10945_);
  and (_10963_, _10962_, _10943_);
  or (_10964_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_10965_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_10966_, _10965_, _04832_);
  and (_10967_, _10966_, _10964_);
  or (_10969_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_10970_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and (_10972_, _10970_, _10928_);
  and (_10973_, _10972_, _10969_);
  or (_10974_, _10973_, _10967_);
  or (_10975_, _10974_, _10926_);
  or (_10976_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_10977_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_10978_, _10977_, _04832_);
  and (_10980_, _10978_, _10976_);
  or (_10982_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_10984_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_10985_, _10984_, _10928_);
  and (_10986_, _10985_, _10982_);
  or (_10987_, _10986_, _10980_);
  or (_10989_, _10987_, _04868_);
  and (_10990_, _10989_, _04859_);
  and (_10992_, _10990_, _10975_);
  or (_10994_, _10992_, _10963_);
  or (_10995_, _10994_, _04849_);
  not (_10996_, _04839_);
  not (_10997_, _04849_);
  and (_10999_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and (_11001_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_11003_, _11001_, _04832_);
  or (_11005_, _11003_, _10999_);
  and (_11006_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_11008_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_11010_, _11008_, _10928_);
  or (_11012_, _11010_, _11006_);
  and (_11013_, _11012_, _11005_);
  or (_11015_, _11013_, _10926_);
  and (_11016_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_11017_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_11019_, _11017_, _04832_);
  or (_11021_, _11019_, _11016_);
  and (_11023_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_11025_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_11026_, _11025_, _10928_);
  or (_11027_, _11026_, _11023_);
  and (_11029_, _11027_, _11021_);
  or (_11031_, _11029_, _04868_);
  and (_11033_, _11031_, _10945_);
  and (_11034_, _11033_, _11015_);
  or (_11035_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_11037_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and (_11038_, _11037_, _11035_);
  or (_11040_, _11038_, _10928_);
  or (_11041_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_11042_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_11044_, _11042_, _11041_);
  or (_11046_, _11044_, _04832_);
  and (_11047_, _11046_, _11040_);
  or (_11048_, _11047_, _10926_);
  or (_11049_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_11050_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_11051_, _11050_, _11049_);
  or (_11052_, _11051_, _10928_);
  or (_11053_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_11054_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and (_11055_, _11054_, _11053_);
  or (_11056_, _11055_, _04832_);
  and (_11057_, _11056_, _11052_);
  or (_11059_, _11057_, _04868_);
  and (_11060_, _11059_, _04859_);
  and (_11062_, _11060_, _11048_);
  or (_11063_, _11062_, _11034_);
  or (_11064_, _11063_, _10997_);
  and (_11066_, _11064_, _10996_);
  and (_11067_, _11066_, _10995_);
  and (_11068_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_11069_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_11070_, _11069_, _11068_);
  and (_11071_, _11070_, _04832_);
  and (_11072_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_11073_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_11074_, _11073_, _11072_);
  and (_11075_, _11074_, _10928_);
  or (_11077_, _11075_, _11071_);
  and (_11079_, _11077_, _04868_);
  and (_11080_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_11081_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_11082_, _11081_, _11080_);
  and (_11083_, _11082_, _04832_);
  and (_11084_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_11085_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_11087_, _11085_, _11084_);
  and (_11089_, _11087_, _10928_);
  or (_11091_, _11089_, _11083_);
  and (_11092_, _11091_, _10926_);
  or (_11093_, _11092_, _11079_);
  and (_11094_, _11093_, _10945_);
  or (_11096_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_11098_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_11100_, _11098_, _11096_);
  and (_11101_, _11100_, _04832_);
  or (_11102_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_11104_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_11105_, _11104_, _11102_);
  and (_11106_, _11105_, _10928_);
  or (_11108_, _11106_, _11101_);
  and (_11110_, _11108_, _04868_);
  or (_11112_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_11114_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_11115_, _11114_, _11112_);
  and (_11116_, _11115_, _04832_);
  or (_11117_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_11118_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_11119_, _11118_, _11117_);
  and (_11120_, _11119_, _10928_);
  or (_11122_, _11120_, _11116_);
  and (_11123_, _11122_, _10926_);
  or (_11125_, _11123_, _11110_);
  and (_11127_, _11125_, _04859_);
  or (_11128_, _11127_, _11094_);
  and (_11129_, _11128_, _10997_);
  and (_11131_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_11133_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_11135_, _11133_, _11131_);
  and (_11137_, _11135_, _04832_);
  and (_11139_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and (_11140_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_11142_, _11140_, _11139_);
  and (_11143_, _11142_, _10928_);
  or (_11144_, _11143_, _11137_);
  and (_11146_, _11144_, _04868_);
  and (_11147_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_11148_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_11150_, _11148_, _11147_);
  and (_11151_, _11150_, _04832_);
  and (_11152_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_11153_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_11155_, _11153_, _11152_);
  and (_11157_, _11155_, _10928_);
  or (_11158_, _11157_, _11151_);
  and (_11160_, _11158_, _10926_);
  or (_11161_, _11160_, _11146_);
  and (_11162_, _11161_, _10945_);
  or (_11164_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_11165_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_11167_, _11165_, _11164_);
  and (_11168_, _11167_, _04832_);
  or (_11169_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_11171_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_11172_, _11171_, _11169_);
  and (_11174_, _11172_, _10928_);
  or (_11175_, _11174_, _11168_);
  and (_11177_, _11175_, _04868_);
  or (_11179_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_11180_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_11181_, _11180_, _11179_);
  and (_11182_, _11181_, _04832_);
  or (_11184_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_11185_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_11186_, _11185_, _11184_);
  and (_11188_, _11186_, _10928_);
  or (_11189_, _11188_, _11182_);
  and (_11191_, _11189_, _10926_);
  or (_11193_, _11191_, _11177_);
  and (_11195_, _11193_, _04859_);
  or (_11196_, _11195_, _11162_);
  and (_11198_, _11196_, _04849_);
  or (_11200_, _11198_, _11129_);
  and (_11201_, _11200_, _04839_);
  or (_11202_, _11201_, _11067_);
  or (_11203_, _11202_, _04843_);
  not (_11204_, _04843_);
  and (_11205_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_11206_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_11207_, _11206_, _11205_);
  and (_11208_, _11207_, _04832_);
  and (_11209_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_11210_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_11211_, _11210_, _11209_);
  and (_11212_, _11211_, _10928_);
  or (_11213_, _11212_, _11208_);
  or (_11214_, _11213_, _10926_);
  and (_11215_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_11216_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_11217_, _11216_, _11215_);
  and (_11218_, _11217_, _04832_);
  and (_11219_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_11220_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_11221_, _11220_, _11219_);
  and (_11222_, _11221_, _10928_);
  or (_11223_, _11222_, _11218_);
  or (_11224_, _11223_, _04868_);
  and (_11225_, _11224_, _10945_);
  and (_11226_, _11225_, _11214_);
  or (_11228_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_11229_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and (_11230_, _11229_, _10928_);
  and (_11231_, _11230_, _11228_);
  or (_11232_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_11233_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_11234_, _11233_, _04832_);
  and (_11235_, _11234_, _11232_);
  or (_11236_, _11235_, _11231_);
  or (_11237_, _11236_, _10926_);
  or (_11238_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_11239_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_11240_, _11239_, _10928_);
  and (_11241_, _11240_, _11238_);
  or (_11242_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_11243_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_11244_, _11243_, _04832_);
  and (_11245_, _11244_, _11242_);
  or (_11246_, _11245_, _11241_);
  or (_11247_, _11246_, _04868_);
  and (_11249_, _11247_, _04859_);
  and (_11250_, _11249_, _11237_);
  or (_11251_, _11250_, _11226_);
  and (_11252_, _11251_, _10997_);
  and (_11253_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_11254_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_11255_, _11254_, _11253_);
  and (_11256_, _11255_, _04832_);
  and (_11257_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_11258_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_11259_, _11258_, _11257_);
  and (_11260_, _11259_, _10928_);
  or (_11261_, _11260_, _11256_);
  or (_11262_, _11261_, _10926_);
  and (_11263_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_11264_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_11265_, _11264_, _11263_);
  and (_11266_, _11265_, _04832_);
  and (_11267_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_11268_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_11270_, _11268_, _11267_);
  and (_11271_, _11270_, _10928_);
  or (_11272_, _11271_, _11266_);
  or (_11273_, _11272_, _04868_);
  and (_11274_, _11273_, _10945_);
  and (_11275_, _11274_, _11262_);
  or (_11276_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_11277_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_11278_, _11277_, _11276_);
  and (_11279_, _11278_, _04832_);
  or (_11280_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_11281_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_11282_, _11281_, _11280_);
  and (_11283_, _11282_, _10928_);
  or (_11284_, _11283_, _11279_);
  or (_11285_, _11284_, _10926_);
  or (_11286_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_11287_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_11288_, _11287_, _11286_);
  and (_11289_, _11288_, _04832_);
  or (_11291_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_11292_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_11293_, _11292_, _11291_);
  and (_11294_, _11293_, _10928_);
  or (_11295_, _11294_, _11289_);
  or (_11296_, _11295_, _04868_);
  and (_11297_, _11296_, _04859_);
  and (_11298_, _11297_, _11285_);
  or (_11299_, _11298_, _11275_);
  and (_11300_, _11299_, _04849_);
  or (_11301_, _11300_, _11252_);
  and (_11302_, _11301_, _10996_);
  or (_11303_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_11304_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_11305_, _11304_, _11303_);
  and (_11306_, _11305_, _04832_);
  or (_11307_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_11308_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_11309_, _11308_, _11307_);
  and (_11310_, _11309_, _10928_);
  or (_11311_, _11310_, _11306_);
  and (_11312_, _11311_, _10926_);
  or (_11313_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_11314_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_11315_, _11314_, _11313_);
  and (_11316_, _11315_, _04832_);
  or (_11317_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_11318_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_11319_, _11318_, _11317_);
  and (_11320_, _11319_, _10928_);
  or (_11321_, _11320_, _11316_);
  and (_11322_, _11321_, _04868_);
  or (_11323_, _11322_, _11312_);
  and (_11325_, _11323_, _04859_);
  and (_11326_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_11327_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_11328_, _11327_, _11326_);
  and (_11329_, _11328_, _04832_);
  and (_11330_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_11332_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_11333_, _11332_, _11330_);
  and (_11334_, _11333_, _10928_);
  or (_11335_, _11334_, _11329_);
  and (_11337_, _11335_, _10926_);
  and (_11338_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_11339_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_11340_, _11339_, _11338_);
  and (_11341_, _11340_, _04832_);
  and (_11342_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_11343_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_11344_, _11343_, _11342_);
  and (_11345_, _11344_, _10928_);
  or (_11346_, _11345_, _11341_);
  and (_11347_, _11346_, _04868_);
  or (_11348_, _11347_, _11337_);
  and (_11349_, _11348_, _10945_);
  or (_11350_, _11349_, _11325_);
  and (_11351_, _11350_, _04849_);
  or (_11352_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_11353_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and (_11354_, _11353_, _10928_);
  and (_11356_, _11354_, _11352_);
  or (_11358_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_11360_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and (_11361_, _11360_, _04832_);
  and (_11362_, _11361_, _11358_);
  or (_11364_, _11362_, _11356_);
  and (_11366_, _11364_, _10926_);
  or (_11367_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_11368_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and (_11369_, _11368_, _10928_);
  and (_11370_, _11369_, _11367_);
  or (_11371_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_11372_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and (_11374_, _11372_, _04832_);
  and (_11375_, _11374_, _11371_);
  or (_11376_, _11375_, _11370_);
  and (_11377_, _11376_, _04868_);
  or (_11378_, _11377_, _11366_);
  and (_11379_, _11378_, _04859_);
  and (_11380_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and (_11381_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_11382_, _11381_, _11380_);
  and (_11383_, _11382_, _04832_);
  and (_11384_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and (_11385_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_11386_, _11385_, _11384_);
  and (_11387_, _11386_, _10928_);
  or (_11388_, _11387_, _11383_);
  and (_11390_, _11388_, _10926_);
  and (_11391_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and (_11392_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_11393_, _11392_, _11391_);
  and (_11394_, _11393_, _04832_);
  and (_11395_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_11396_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_11397_, _11396_, _11395_);
  and (_11398_, _11397_, _10928_);
  or (_11399_, _11398_, _11394_);
  and (_11400_, _11399_, _04868_);
  or (_11401_, _11400_, _11390_);
  and (_11402_, _11401_, _10945_);
  or (_11403_, _11402_, _11379_);
  and (_11405_, _11403_, _10997_);
  or (_11407_, _11405_, _11351_);
  and (_11408_, _11407_, _04839_);
  or (_11409_, _11408_, _11302_);
  or (_11410_, _11409_, _11204_);
  and (_11411_, _11410_, _11203_);
  or (_11412_, _11411_, _26153_);
  and (_11413_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_11414_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_11416_, _11414_, _11413_);
  and (_11418_, _11416_, _04832_);
  and (_11419_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_11420_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_11421_, _11420_, _11419_);
  and (_11422_, _11421_, _10928_);
  or (_11424_, _11422_, _11418_);
  or (_11425_, _11424_, _10926_);
  and (_11426_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_11427_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_11428_, _11427_, _11426_);
  and (_11429_, _11428_, _04832_);
  and (_11431_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_11432_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_11433_, _11432_, _11431_);
  and (_11434_, _11433_, _10928_);
  or (_11435_, _11434_, _11429_);
  or (_11436_, _11435_, _04868_);
  and (_11437_, _11436_, _10945_);
  and (_11438_, _11437_, _11425_);
  or (_11439_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_11441_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_11442_, _11441_, _11439_);
  and (_11443_, _11442_, _04832_);
  or (_11445_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_11446_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_11447_, _11446_, _11445_);
  and (_11448_, _11447_, _10928_);
  or (_11449_, _11448_, _11443_);
  or (_11451_, _11449_, _10926_);
  or (_11452_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_11454_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_11455_, _11454_, _11452_);
  and (_11457_, _11455_, _04832_);
  or (_11458_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_11460_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_11461_, _11460_, _11458_);
  and (_11463_, _11461_, _10928_);
  or (_11464_, _11463_, _11457_);
  or (_11465_, _11464_, _04868_);
  and (_11466_, _11465_, _04859_);
  and (_11467_, _11466_, _11451_);
  or (_11468_, _11467_, _11438_);
  and (_11470_, _11468_, _04849_);
  and (_11471_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_11473_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_11474_, _11473_, _11471_);
  and (_11475_, _11474_, _04832_);
  and (_11476_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_11477_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_11478_, _11477_, _11476_);
  and (_11479_, _11478_, _10928_);
  or (_11481_, _11479_, _11475_);
  or (_11482_, _11481_, _10926_);
  and (_11483_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_11484_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_11485_, _11484_, _11483_);
  and (_11486_, _11485_, _04832_);
  and (_11487_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_11488_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_11489_, _11488_, _11487_);
  and (_11490_, _11489_, _10928_);
  or (_11491_, _11490_, _11486_);
  or (_11493_, _11491_, _04868_);
  and (_11494_, _11493_, _10945_);
  and (_11495_, _11494_, _11482_);
  or (_11496_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_11498_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_11501_, _11498_, _10928_);
  and (_11502_, _11501_, _11496_);
  or (_11503_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_11504_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_11505_, _11504_, _04832_);
  and (_11506_, _11505_, _11503_);
  or (_11507_, _11506_, _11502_);
  or (_11508_, _11507_, _10926_);
  or (_11509_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_11510_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_11511_, _11510_, _10928_);
  and (_11512_, _11511_, _11509_);
  or (_11513_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_11514_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_11515_, _11514_, _04832_);
  and (_11516_, _11515_, _11513_);
  or (_11517_, _11516_, _11512_);
  or (_11518_, _11517_, _04868_);
  and (_11519_, _11518_, _04859_);
  and (_11520_, _11519_, _11508_);
  or (_11521_, _11520_, _11495_);
  and (_11523_, _11521_, _10997_);
  or (_11524_, _11523_, _11470_);
  and (_11525_, _11524_, _10996_);
  and (_11526_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_11527_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_11528_, _11527_, _11526_);
  and (_11529_, _11528_, _04832_);
  and (_11530_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_11531_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_11532_, _11531_, _11530_);
  and (_11533_, _11532_, _10928_);
  or (_11534_, _11533_, _11529_);
  and (_11535_, _11534_, _04868_);
  and (_11536_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_11537_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_11539_, _11537_, _11536_);
  and (_11540_, _11539_, _04832_);
  and (_11542_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_11543_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_11544_, _11543_, _11542_);
  and (_11545_, _11544_, _10928_);
  or (_11546_, _11545_, _11540_);
  and (_11547_, _11546_, _10926_);
  or (_11548_, _11547_, _11535_);
  and (_11549_, _11548_, _10945_);
  or (_11550_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_11551_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_11553_, _11551_, _10928_);
  and (_11555_, _11553_, _11550_);
  or (_11556_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_11557_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_11558_, _11557_, _04832_);
  and (_11559_, _11558_, _11556_);
  or (_11560_, _11559_, _11555_);
  and (_11561_, _11560_, _04868_);
  or (_11562_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_11563_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_11564_, _11563_, _10928_);
  and (_11565_, _11564_, _11562_);
  or (_11567_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_11568_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_11569_, _11568_, _04832_);
  and (_11571_, _11569_, _11567_);
  or (_11573_, _11571_, _11565_);
  and (_11574_, _11573_, _10926_);
  or (_11575_, _11574_, _11561_);
  and (_11576_, _11575_, _04859_);
  or (_11577_, _11576_, _11549_);
  and (_11578_, _11577_, _10997_);
  and (_11579_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_11580_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_11581_, _11580_, _11579_);
  and (_11582_, _11581_, _04832_);
  and (_11583_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_11584_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_11585_, _11584_, _11583_);
  and (_11586_, _11585_, _10928_);
  or (_11587_, _11586_, _11582_);
  and (_11588_, _11587_, _04868_);
  and (_11589_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_11590_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_11592_, _11590_, _11589_);
  and (_11593_, _11592_, _04832_);
  and (_11594_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_11595_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_11596_, _11595_, _11594_);
  and (_11597_, _11596_, _10928_);
  or (_11598_, _11597_, _11593_);
  and (_11599_, _11598_, _10926_);
  or (_11600_, _11599_, _11588_);
  and (_11601_, _11600_, _10945_);
  or (_11602_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_11603_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_11604_, _11603_, _11602_);
  and (_11606_, _11604_, _04832_);
  or (_11608_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_11610_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_11612_, _11610_, _11608_);
  and (_11613_, _11612_, _10928_);
  or (_11614_, _11613_, _11606_);
  and (_11615_, _11614_, _04868_);
  or (_11616_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_11618_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_11620_, _11618_, _11616_);
  and (_11622_, _11620_, _04832_);
  or (_11623_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_11624_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_11625_, _11624_, _11623_);
  and (_11626_, _11625_, _10928_);
  or (_11628_, _11626_, _11622_);
  and (_11629_, _11628_, _10926_);
  or (_11630_, _11629_, _11615_);
  and (_11631_, _11630_, _04859_);
  or (_11632_, _11631_, _11601_);
  and (_11634_, _11632_, _04849_);
  or (_11635_, _11634_, _11578_);
  and (_11636_, _11635_, _04839_);
  or (_11638_, _11636_, _11525_);
  or (_11640_, _11638_, _04843_);
  and (_11642_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_11644_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_11646_, _11644_, _11642_);
  and (_11648_, _11646_, _04832_);
  and (_11650_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_11652_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_11654_, _11652_, _11650_);
  and (_11656_, _11654_, _10928_);
  or (_11658_, _11656_, _11648_);
  or (_11660_, _11658_, _10926_);
  and (_11662_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_11664_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_11666_, _11664_, _11662_);
  and (_11668_, _11666_, _04832_);
  and (_11669_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_11671_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_11672_, _11671_, _11669_);
  and (_11673_, _11672_, _10928_);
  or (_11675_, _11673_, _11668_);
  or (_11676_, _11675_, _04868_);
  and (_11677_, _11676_, _10945_);
  and (_11679_, _11677_, _11660_);
  or (_11681_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_11682_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_11683_, _11682_, _10928_);
  and (_11684_, _11683_, _11681_);
  or (_11686_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_11687_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_11688_, _11687_, _04832_);
  and (_11690_, _11688_, _11686_);
  or (_11691_, _11690_, _11684_);
  or (_11693_, _11691_, _10926_);
  or (_11694_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_11695_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_11696_, _11695_, _10928_);
  and (_11697_, _11696_, _11694_);
  or (_11698_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_11699_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_11700_, _11699_, _04832_);
  and (_11701_, _11700_, _11698_);
  or (_11702_, _11701_, _11697_);
  or (_11703_, _11702_, _04868_);
  and (_11704_, _11703_, _04859_);
  and (_11705_, _11704_, _11693_);
  or (_11706_, _11705_, _11679_);
  and (_11707_, _11706_, _10997_);
  and (_11708_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_11709_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_11710_, _11709_, _11708_);
  and (_11711_, _11710_, _04832_);
  and (_11712_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_11713_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_11714_, _11713_, _11712_);
  and (_11715_, _11714_, _10928_);
  or (_11717_, _11715_, _11711_);
  or (_11718_, _11717_, _10926_);
  and (_11719_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_11720_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_11722_, _11720_, _11719_);
  and (_11723_, _11722_, _04832_);
  and (_11725_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_11726_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_11728_, _11726_, _11725_);
  and (_11729_, _11728_, _10928_);
  or (_11730_, _11729_, _11723_);
  or (_11731_, _11730_, _04868_);
  and (_11732_, _11731_, _10945_);
  and (_11733_, _11732_, _11718_);
  or (_11734_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_11735_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_11737_, _11735_, _11734_);
  and (_11738_, _11737_, _04832_);
  or (_11739_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_11740_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_11741_, _11740_, _11739_);
  and (_11742_, _11741_, _10928_);
  or (_11743_, _11742_, _11738_);
  or (_11744_, _11743_, _10926_);
  or (_11745_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_11746_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_11747_, _11746_, _11745_);
  and (_11748_, _11747_, _04832_);
  or (_11749_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_11750_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_11751_, _11750_, _11749_);
  and (_11752_, _11751_, _10928_);
  or (_11753_, _11752_, _11748_);
  or (_11754_, _11753_, _04868_);
  and (_11755_, _11754_, _04859_);
  and (_11756_, _11755_, _11744_);
  or (_11757_, _11756_, _11733_);
  and (_11758_, _11757_, _04849_);
  or (_11759_, _11758_, _11707_);
  and (_11760_, _11759_, _10996_);
  or (_11761_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_11762_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_11763_, _11762_, _11761_);
  and (_11764_, _11763_, _04832_);
  or (_11765_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_11766_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_11767_, _11766_, _11765_);
  and (_11768_, _11767_, _10928_);
  or (_11769_, _11768_, _11764_);
  and (_11770_, _11769_, _10926_);
  or (_11771_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_11772_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_11773_, _11772_, _11771_);
  and (_11774_, _11773_, _04832_);
  or (_11775_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_11776_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_11777_, _11776_, _11775_);
  and (_11778_, _11777_, _10928_);
  or (_11779_, _11778_, _11774_);
  and (_11780_, _11779_, _04868_);
  or (_11781_, _11780_, _11770_);
  and (_11782_, _11781_, _04859_);
  and (_11783_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_11784_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_11785_, _11784_, _11783_);
  and (_11786_, _11785_, _04832_);
  and (_11787_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_11788_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_11789_, _11788_, _11787_);
  and (_11790_, _11789_, _10928_);
  or (_11791_, _11790_, _11786_);
  and (_11792_, _11791_, _10926_);
  and (_11793_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_11794_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_11795_, _11794_, _11793_);
  and (_11796_, _11795_, _04832_);
  and (_11797_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_11798_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_11799_, _11798_, _11797_);
  and (_11800_, _11799_, _10928_);
  or (_11801_, _11800_, _11796_);
  and (_11802_, _11801_, _04868_);
  or (_11803_, _11802_, _11792_);
  and (_11804_, _11803_, _10945_);
  or (_11805_, _11804_, _11782_);
  and (_11806_, _11805_, _04849_);
  or (_11807_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_11808_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and (_11809_, _11808_, _10928_);
  and (_11810_, _11809_, _11807_);
  or (_11811_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_11812_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and (_11813_, _11812_, _04832_);
  and (_11814_, _11813_, _11811_);
  or (_11815_, _11814_, _11810_);
  and (_11816_, _11815_, _10926_);
  or (_11817_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_11818_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_11819_, _11818_, _10928_);
  and (_11820_, _11819_, _11817_);
  or (_11821_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_11822_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and (_11823_, _11822_, _04832_);
  and (_11824_, _11823_, _11821_);
  or (_11825_, _11824_, _11820_);
  and (_11826_, _11825_, _04868_);
  or (_11827_, _11826_, _11816_);
  and (_11828_, _11827_, _04859_);
  and (_11830_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and (_11831_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_11832_, _11831_, _11830_);
  and (_11834_, _11832_, _04832_);
  and (_11835_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and (_11837_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_11838_, _11837_, _11835_);
  and (_11839_, _11838_, _10928_);
  or (_11841_, _11839_, _11834_);
  and (_11843_, _11841_, _10926_);
  and (_11844_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_11846_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_11847_, _11846_, _11844_);
  and (_11848_, _11847_, _04832_);
  and (_11850_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and (_11852_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_11854_, _11852_, _11850_);
  and (_11856_, _11854_, _10928_);
  or (_11857_, _11856_, _11848_);
  and (_11858_, _11857_, _04868_);
  or (_11859_, _11858_, _11843_);
  and (_11860_, _11859_, _10945_);
  or (_11862_, _11860_, _11828_);
  and (_11863_, _11862_, _10997_);
  or (_11865_, _11863_, _11806_);
  and (_11867_, _11865_, _04839_);
  or (_11869_, _11867_, _11760_);
  or (_11870_, _11869_, _11204_);
  and (_11873_, _11870_, _11640_);
  or (_11874_, _11873_, _03196_);
  and (_11876_, _11874_, _11412_);
  or (_11877_, _11876_, _04876_);
  not (_11878_, _04876_);
  or (_11879_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_11880_, _11879_, _22773_);
  and (_05818_, _11880_, _11877_);
  and (_11881_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_11882_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_11883_, _11882_, _11881_);
  and (_11884_, _11883_, _04832_);
  and (_11885_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_11886_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_11887_, _11886_, _11885_);
  and (_11888_, _11887_, _10928_);
  or (_11889_, _11888_, _11884_);
  or (_11890_, _11889_, _10926_);
  and (_11891_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_11892_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_11893_, _11892_, _11891_);
  and (_11894_, _11893_, _04832_);
  and (_11895_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and (_11896_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_11897_, _11896_, _11895_);
  and (_11898_, _11897_, _10928_);
  or (_11899_, _11898_, _11894_);
  or (_11900_, _11899_, _04868_);
  and (_11901_, _11900_, _10945_);
  and (_11902_, _11901_, _11890_);
  or (_11903_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_11904_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_11905_, _11904_, _11903_);
  and (_11906_, _11905_, _04832_);
  or (_11907_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_11908_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_11909_, _11908_, _11907_);
  and (_11910_, _11909_, _10928_);
  or (_11911_, _11910_, _11906_);
  or (_11912_, _11911_, _10926_);
  or (_11913_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_11914_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and (_11915_, _11914_, _11913_);
  and (_11916_, _11915_, _04832_);
  or (_11917_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_11918_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_11919_, _11918_, _11917_);
  and (_11920_, _11919_, _10928_);
  or (_11921_, _11920_, _11916_);
  or (_11922_, _11921_, _04868_);
  and (_11923_, _11922_, _04859_);
  and (_11924_, _11923_, _11912_);
  or (_11925_, _11924_, _11902_);
  or (_11926_, _11925_, _10997_);
  and (_11927_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_11928_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_11929_, _11928_, _11927_);
  and (_11930_, _11929_, _04832_);
  and (_11931_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_11932_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_11933_, _11932_, _11931_);
  and (_11934_, _11933_, _10928_);
  or (_11935_, _11934_, _11930_);
  or (_11936_, _11935_, _10926_);
  and (_11937_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and (_11938_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_11939_, _11938_, _11937_);
  and (_11940_, _11939_, _04832_);
  and (_11941_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_11942_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_11943_, _11942_, _11941_);
  and (_11944_, _11943_, _10928_);
  or (_11945_, _11944_, _11940_);
  or (_11946_, _11945_, _04868_);
  and (_11947_, _11946_, _10945_);
  and (_11948_, _11947_, _11936_);
  or (_11949_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_11950_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and (_11951_, _11950_, _10928_);
  and (_11952_, _11951_, _11949_);
  or (_11953_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_11954_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_11955_, _11954_, _04832_);
  and (_11956_, _11955_, _11953_);
  or (_11957_, _11956_, _11952_);
  or (_11958_, _11957_, _10926_);
  or (_11959_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_11960_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and (_11961_, _11960_, _10928_);
  and (_11962_, _11961_, _11959_);
  or (_11963_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_11964_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_11965_, _11964_, _04832_);
  and (_11966_, _11965_, _11963_);
  or (_11967_, _11966_, _11962_);
  or (_11968_, _11967_, _04868_);
  and (_11969_, _11968_, _04859_);
  and (_11970_, _11969_, _11958_);
  or (_11971_, _11970_, _11948_);
  or (_11972_, _11971_, _04849_);
  and (_11973_, _11972_, _10996_);
  and (_11974_, _11973_, _11926_);
  and (_11975_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_11976_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_11977_, _11976_, _11975_);
  and (_11978_, _11977_, _04832_);
  and (_11979_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_11980_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_11981_, _11980_, _11979_);
  and (_11982_, _11981_, _10928_);
  or (_11984_, _11982_, _11978_);
  and (_11985_, _11984_, _04868_);
  and (_11986_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_11987_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_11988_, _11987_, _11986_);
  and (_11989_, _11988_, _04832_);
  and (_11990_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_11991_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_11992_, _11991_, _11990_);
  and (_11993_, _11992_, _10928_);
  or (_11994_, _11993_, _11989_);
  and (_11995_, _11994_, _10926_);
  or (_11996_, _11995_, _04859_);
  or (_11997_, _11996_, _11985_);
  or (_11998_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_11999_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_12000_, _11999_, _10928_);
  and (_12001_, _12000_, _11998_);
  or (_12002_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_12003_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_12005_, _12003_, _04832_);
  and (_12006_, _12005_, _12002_);
  or (_12007_, _12006_, _12001_);
  and (_12008_, _12007_, _04868_);
  or (_12009_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_12010_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_12011_, _12010_, _10928_);
  and (_12012_, _12011_, _12009_);
  or (_12013_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_12014_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_12015_, _12014_, _04832_);
  and (_12016_, _12015_, _12013_);
  or (_12017_, _12016_, _12012_);
  and (_12018_, _12017_, _10926_);
  or (_12019_, _12018_, _10945_);
  or (_12020_, _12019_, _12008_);
  and (_12021_, _12020_, _11997_);
  or (_12022_, _12021_, _04849_);
  and (_12023_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and (_12024_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_12025_, _12024_, _12023_);
  and (_12026_, _12025_, _04832_);
  and (_12027_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_12028_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_12029_, _12028_, _12027_);
  and (_12030_, _12029_, _10928_);
  or (_12031_, _12030_, _12026_);
  and (_12032_, _12031_, _04868_);
  and (_12033_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_12034_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_12035_, _12034_, _12033_);
  and (_12036_, _12035_, _04832_);
  and (_12037_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_12038_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_12039_, _12038_, _12037_);
  and (_12040_, _12039_, _10928_);
  or (_12041_, _12040_, _12036_);
  and (_12042_, _12041_, _10926_);
  or (_12043_, _12042_, _04859_);
  or (_12044_, _12043_, _12032_);
  or (_12045_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_12046_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and (_12047_, _12046_, _12045_);
  and (_12048_, _12047_, _04832_);
  or (_12049_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_12050_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_12051_, _12050_, _12049_);
  and (_12052_, _12051_, _10928_);
  or (_12053_, _12052_, _12048_);
  and (_12054_, _12053_, _04868_);
  or (_12055_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_12056_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_12057_, _12056_, _12055_);
  and (_12058_, _12057_, _04832_);
  or (_12059_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_12060_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_12061_, _12060_, _12059_);
  and (_12062_, _12061_, _10928_);
  or (_12063_, _12062_, _12058_);
  and (_12064_, _12063_, _10926_);
  or (_12065_, _12064_, _10945_);
  or (_12066_, _12065_, _12054_);
  and (_12067_, _12066_, _12044_);
  or (_12068_, _12067_, _10997_);
  and (_12069_, _12068_, _04839_);
  and (_12070_, _12069_, _12022_);
  or (_12071_, _12070_, _11974_);
  or (_12072_, _12071_, _04843_);
  and (_12073_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and (_12074_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_12075_, _12074_, _12073_);
  and (_12077_, _12075_, _04832_);
  and (_12079_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and (_12080_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_12081_, _12080_, _12079_);
  and (_12083_, _12081_, _10928_);
  or (_12084_, _12083_, _12077_);
  and (_12085_, _12084_, _04868_);
  and (_12087_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  and (_12089_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_12091_, _12089_, _12087_);
  and (_12093_, _12091_, _04832_);
  and (_12095_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and (_12096_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_12097_, _12096_, _12095_);
  and (_12098_, _12097_, _10928_);
  or (_12099_, _12098_, _12093_);
  and (_12100_, _12099_, _10926_);
  or (_12101_, _12100_, _04859_);
  or (_12102_, _12101_, _12085_);
  or (_12103_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_12104_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and (_12106_, _12104_, _12103_);
  and (_12107_, _12106_, _04832_);
  or (_12108_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_12109_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  and (_12110_, _12109_, _12108_);
  and (_12111_, _12110_, _10928_);
  or (_12112_, _12111_, _12107_);
  and (_12113_, _12112_, _04868_);
  or (_12114_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_12115_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  and (_12116_, _12115_, _12114_);
  and (_12117_, _12116_, _04832_);
  or (_12118_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_12119_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and (_12120_, _12119_, _12118_);
  and (_12121_, _12120_, _10928_);
  or (_12122_, _12121_, _12117_);
  and (_12123_, _12122_, _10926_);
  or (_12124_, _12123_, _10945_);
  or (_12125_, _12124_, _12113_);
  and (_12126_, _12125_, _12102_);
  or (_12127_, _12126_, _04849_);
  and (_12128_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_12129_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_12130_, _12129_, _12128_);
  and (_12131_, _12130_, _04832_);
  and (_12132_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and (_12133_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_12134_, _12133_, _12132_);
  and (_12135_, _12134_, _10928_);
  or (_12136_, _12135_, _12131_);
  and (_12137_, _12136_, _04868_);
  and (_12138_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_12139_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_12140_, _12139_, _12138_);
  and (_12141_, _12140_, _04832_);
  and (_12143_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and (_12144_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_12145_, _12144_, _12143_);
  and (_12146_, _12145_, _10928_);
  or (_12147_, _12146_, _12141_);
  and (_12149_, _12147_, _10926_);
  or (_12150_, _12149_, _04859_);
  or (_12151_, _12150_, _12137_);
  or (_12152_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_12153_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_12154_, _12153_, _12152_);
  and (_12155_, _12154_, _04832_);
  or (_12156_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_12157_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and (_12158_, _12157_, _12156_);
  and (_12159_, _12158_, _10928_);
  or (_12160_, _12159_, _12155_);
  and (_12161_, _12160_, _04868_);
  or (_12162_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_12163_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_12164_, _12163_, _12162_);
  and (_12165_, _12164_, _04832_);
  or (_12166_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_12167_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and (_12168_, _12167_, _12166_);
  and (_12169_, _12168_, _10928_);
  or (_12170_, _12169_, _12165_);
  and (_12171_, _12170_, _10926_);
  or (_12172_, _12171_, _10945_);
  or (_12173_, _12172_, _12161_);
  and (_12174_, _12173_, _12151_);
  or (_12175_, _12174_, _10997_);
  and (_12176_, _12175_, _04839_);
  and (_12177_, _12176_, _12127_);
  and (_12178_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_12179_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_12180_, _12179_, _12178_);
  and (_12181_, _12180_, _10928_);
  and (_12182_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and (_12183_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_12184_, _12183_, _12182_);
  and (_12185_, _12184_, _04832_);
  or (_12186_, _12185_, _12181_);
  or (_12187_, _12186_, _10926_);
  and (_12188_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_12189_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_12190_, _12189_, _12188_);
  and (_12191_, _12190_, _10928_);
  and (_12192_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and (_12193_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_12194_, _12193_, _12192_);
  and (_12195_, _12194_, _04832_);
  or (_12196_, _12195_, _12191_);
  or (_12197_, _12196_, _04868_);
  and (_12198_, _12197_, _10945_);
  and (_12199_, _12198_, _12187_);
  or (_12200_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_12202_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_12204_, _12202_, _04832_);
  and (_12205_, _12204_, _12200_);
  or (_12206_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_12207_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_12208_, _12207_, _10928_);
  and (_12209_, _12208_, _12206_);
  or (_12210_, _12209_, _12205_);
  or (_12211_, _12210_, _10926_);
  or (_12212_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_12213_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and (_12214_, _12213_, _04832_);
  and (_12215_, _12214_, _12212_);
  or (_12217_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_12218_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_12221_, _12218_, _10928_);
  and (_12222_, _12221_, _12217_);
  or (_12223_, _12222_, _12215_);
  or (_12224_, _12223_, _04868_);
  and (_12225_, _12224_, _04859_);
  and (_12226_, _12225_, _12211_);
  or (_12227_, _12226_, _12199_);
  and (_12228_, _12227_, _10997_);
  and (_12229_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_12230_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_12231_, _12230_, _04832_);
  or (_12232_, _12231_, _12229_);
  and (_12233_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_12234_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_12235_, _12234_, _10928_);
  or (_12236_, _12235_, _12233_);
  and (_12237_, _12236_, _12232_);
  or (_12238_, _12237_, _10926_);
  and (_12239_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_12240_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_12241_, _12240_, _04832_);
  or (_12242_, _12241_, _12239_);
  and (_12243_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_12244_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_12245_, _12244_, _10928_);
  or (_12246_, _12245_, _12243_);
  and (_12247_, _12246_, _12242_);
  or (_12248_, _12247_, _04868_);
  and (_12249_, _12248_, _10945_);
  and (_12250_, _12249_, _12238_);
  or (_12251_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_12252_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_12253_, _12252_, _12251_);
  or (_12254_, _12253_, _10928_);
  or (_12255_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_12256_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_12257_, _12256_, _12255_);
  or (_12258_, _12257_, _04832_);
  and (_12260_, _12258_, _12254_);
  or (_12262_, _12260_, _10926_);
  or (_12263_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_12264_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_12265_, _12264_, _12263_);
  or (_12266_, _12265_, _10928_);
  or (_12267_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_12268_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_12270_, _12268_, _12267_);
  or (_12271_, _12270_, _04832_);
  and (_12272_, _12271_, _12266_);
  or (_12274_, _12272_, _04868_);
  and (_12275_, _12274_, _04859_);
  and (_12276_, _12275_, _12262_);
  or (_12277_, _12276_, _12250_);
  and (_12279_, _12277_, _04849_);
  or (_12280_, _12279_, _12228_);
  and (_12281_, _12280_, _10996_);
  or (_12282_, _12281_, _12177_);
  or (_12283_, _12282_, _11204_);
  and (_12284_, _12283_, _12072_);
  or (_12286_, _12284_, _26153_);
  and (_12287_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_12288_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_12289_, _12288_, _12287_);
  and (_12290_, _12289_, _10928_);
  and (_12291_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_12292_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_12293_, _12292_, _12291_);
  and (_12294_, _12293_, _04832_);
  or (_12295_, _12294_, _12290_);
  or (_12296_, _12295_, _10926_);
  and (_12298_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_12300_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_12301_, _12300_, _12298_);
  and (_12302_, _12301_, _10928_);
  and (_12303_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_12304_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_12305_, _12304_, _12303_);
  and (_12306_, _12305_, _04832_);
  or (_12307_, _12306_, _12302_);
  or (_12308_, _12307_, _04868_);
  and (_12310_, _12308_, _10945_);
  and (_12311_, _12310_, _12296_);
  or (_12312_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_12314_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_12315_, _12314_, _04832_);
  and (_12316_, _12315_, _12312_);
  or (_12317_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_12318_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_12320_, _12318_, _10928_);
  and (_12321_, _12320_, _12317_);
  or (_12322_, _12321_, _12316_);
  or (_12323_, _12322_, _10926_);
  or (_12324_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_12325_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_12327_, _12325_, _04832_);
  and (_12328_, _12327_, _12324_);
  or (_12329_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_12330_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_12331_, _12330_, _10928_);
  and (_12332_, _12331_, _12329_);
  or (_12334_, _12332_, _12328_);
  or (_12335_, _12334_, _04868_);
  and (_12336_, _12335_, _04859_);
  and (_12337_, _12336_, _12323_);
  or (_12339_, _12337_, _12311_);
  and (_12341_, _12339_, _10997_);
  and (_12343_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_12344_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_12345_, _12344_, _04832_);
  or (_12347_, _12345_, _12343_);
  and (_12348_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_12349_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_12350_, _12349_, _10928_);
  or (_12351_, _12350_, _12348_);
  and (_12352_, _12351_, _12347_);
  or (_12353_, _12352_, _10926_);
  and (_12354_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_12355_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_12356_, _12355_, _04832_);
  or (_12357_, _12356_, _12354_);
  and (_12359_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_12360_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_12361_, _12360_, _10928_);
  or (_12362_, _12361_, _12359_);
  and (_12363_, _12362_, _12357_);
  or (_12364_, _12363_, _04868_);
  and (_12365_, _12364_, _10945_);
  and (_12366_, _12365_, _12353_);
  or (_12367_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_12368_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_12369_, _12368_, _12367_);
  or (_12370_, _12369_, _10928_);
  or (_12371_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_12372_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_12373_, _12372_, _12371_);
  or (_12374_, _12373_, _04832_);
  and (_12375_, _12374_, _12370_);
  or (_12376_, _12375_, _10926_);
  or (_12377_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_12378_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_12379_, _12378_, _12377_);
  or (_12380_, _12379_, _10928_);
  or (_12381_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_12382_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_12383_, _12382_, _12381_);
  or (_12384_, _12383_, _04832_);
  and (_12385_, _12384_, _12380_);
  or (_12386_, _12385_, _04868_);
  and (_12387_, _12386_, _04859_);
  and (_12388_, _12387_, _12376_);
  or (_12389_, _12388_, _12366_);
  and (_12390_, _12389_, _04849_);
  or (_12391_, _12390_, _12341_);
  and (_12392_, _12391_, _10996_);
  and (_12393_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and (_12394_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or (_12395_, _12394_, _12393_);
  and (_12396_, _12395_, _04832_);
  and (_12397_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  and (_12398_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or (_12400_, _12398_, _12397_);
  and (_12401_, _12400_, _10928_);
  or (_12402_, _12401_, _12396_);
  and (_12403_, _12402_, _04868_);
  and (_12404_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and (_12405_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or (_12406_, _12405_, _12404_);
  and (_12407_, _12406_, _04832_);
  and (_12408_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and (_12409_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or (_12410_, _12409_, _12408_);
  and (_12411_, _12410_, _10928_);
  or (_12412_, _12411_, _12407_);
  and (_12413_, _12412_, _10926_);
  or (_12414_, _12413_, _12403_);
  and (_12415_, _12414_, _10945_);
  or (_12416_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or (_12417_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  and (_12418_, _12417_, _12416_);
  and (_12419_, _12418_, _04832_);
  or (_12421_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or (_12422_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and (_12423_, _12422_, _12421_);
  and (_12424_, _12423_, _10928_);
  or (_12425_, _12424_, _12419_);
  and (_12426_, _12425_, _04868_);
  or (_12427_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or (_12428_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and (_12429_, _12428_, _12427_);
  and (_12430_, _12429_, _04832_);
  or (_12431_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or (_12432_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and (_12433_, _12432_, _12431_);
  and (_12434_, _12433_, _10928_);
  or (_12435_, _12434_, _12430_);
  and (_12436_, _12435_, _10926_);
  or (_12437_, _12436_, _12426_);
  and (_12438_, _12437_, _04859_);
  or (_12439_, _12438_, _12415_);
  and (_12440_, _12439_, _10997_);
  and (_12441_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_12442_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_12443_, _12442_, _12441_);
  and (_12444_, _12443_, _04832_);
  and (_12445_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_12446_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_12447_, _12446_, _12445_);
  and (_12448_, _12447_, _10928_);
  or (_12449_, _12448_, _12444_);
  and (_12450_, _12449_, _04868_);
  and (_12451_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_12452_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_12453_, _12452_, _12451_);
  and (_12454_, _12453_, _04832_);
  and (_12455_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_12456_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_12457_, _12456_, _12455_);
  and (_12458_, _12457_, _10928_);
  or (_12459_, _12458_, _12454_);
  and (_12460_, _12459_, _10926_);
  or (_12461_, _12460_, _12450_);
  and (_12462_, _12461_, _10945_);
  or (_12463_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_12464_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_12465_, _12464_, _12463_);
  and (_12466_, _12465_, _04832_);
  or (_12467_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_12468_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_12469_, _12468_, _12467_);
  and (_12470_, _12469_, _10928_);
  or (_12471_, _12470_, _12466_);
  and (_12472_, _12471_, _04868_);
  or (_12473_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_12474_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_12475_, _12474_, _12473_);
  and (_12476_, _12475_, _04832_);
  or (_12477_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_12478_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_12479_, _12478_, _12477_);
  and (_12480_, _12479_, _10928_);
  or (_12481_, _12480_, _12476_);
  and (_12482_, _12481_, _10926_);
  or (_12483_, _12482_, _12472_);
  and (_12484_, _12483_, _04859_);
  or (_12485_, _12484_, _12462_);
  and (_12486_, _12485_, _04849_);
  or (_12487_, _12486_, _12440_);
  and (_12488_, _12487_, _04839_);
  or (_12489_, _12488_, _12392_);
  or (_12490_, _12489_, _04843_);
  and (_12491_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_12492_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_12493_, _12492_, _12491_);
  and (_12494_, _12493_, _04832_);
  and (_12495_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_12496_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_12497_, _12496_, _12495_);
  and (_12498_, _12497_, _10928_);
  or (_12499_, _12498_, _12494_);
  or (_12500_, _12499_, _10926_);
  and (_12501_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_12502_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_12503_, _12502_, _12501_);
  and (_12504_, _12503_, _04832_);
  and (_12505_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_12506_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_12507_, _12506_, _12505_);
  and (_12508_, _12507_, _10928_);
  or (_12509_, _12508_, _12504_);
  or (_12510_, _12509_, _04868_);
  and (_12511_, _12510_, _10945_);
  and (_12512_, _12511_, _12500_);
  or (_12513_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_12514_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_12515_, _12514_, _10928_);
  and (_12516_, _12515_, _12513_);
  or (_12517_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_12518_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_12519_, _12518_, _04832_);
  and (_12520_, _12519_, _12517_);
  or (_12521_, _12520_, _12516_);
  or (_12522_, _12521_, _10926_);
  or (_12523_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_12524_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_12525_, _12524_, _10928_);
  and (_12526_, _12525_, _12523_);
  or (_12527_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_12528_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_12529_, _12528_, _04832_);
  and (_12530_, _12529_, _12527_);
  or (_12531_, _12530_, _12526_);
  or (_12532_, _12531_, _04868_);
  and (_12533_, _12532_, _04859_);
  and (_12534_, _12533_, _12522_);
  or (_12535_, _12534_, _12512_);
  and (_12536_, _12535_, _10997_);
  and (_12537_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_12538_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_12539_, _12538_, _12537_);
  and (_12540_, _12539_, _04832_);
  and (_12541_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_12542_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_12543_, _12542_, _12541_);
  and (_12544_, _12543_, _10928_);
  or (_12545_, _12544_, _12540_);
  or (_12546_, _12545_, _10926_);
  and (_12547_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_12548_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_12549_, _12548_, _12547_);
  and (_12550_, _12549_, _04832_);
  and (_12551_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_12552_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_12553_, _12552_, _12551_);
  and (_12554_, _12553_, _10928_);
  or (_12555_, _12554_, _12550_);
  or (_12556_, _12555_, _04868_);
  and (_12557_, _12556_, _10945_);
  and (_12558_, _12557_, _12546_);
  or (_12559_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_12560_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_12561_, _12560_, _12559_);
  and (_12562_, _12561_, _04832_);
  or (_12563_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_12564_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_12565_, _12564_, _12563_);
  and (_12566_, _12565_, _10928_);
  or (_12567_, _12566_, _12562_);
  or (_12568_, _12567_, _10926_);
  or (_12569_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_12570_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_12571_, _12570_, _12569_);
  and (_12572_, _12571_, _04832_);
  or (_12573_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_12574_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_12575_, _12574_, _12573_);
  and (_12576_, _12575_, _10928_);
  or (_12577_, _12576_, _12572_);
  or (_12578_, _12577_, _04868_);
  and (_12579_, _12578_, _04859_);
  and (_12580_, _12579_, _12568_);
  or (_12581_, _12580_, _12558_);
  and (_12582_, _12581_, _04849_);
  or (_12583_, _12582_, _12536_);
  and (_12584_, _12583_, _10996_);
  or (_12585_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_12586_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_12587_, _12586_, _12585_);
  and (_12588_, _12587_, _04832_);
  or (_12589_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_12590_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_12591_, _12590_, _12589_);
  and (_12592_, _12591_, _10928_);
  or (_12593_, _12592_, _12588_);
  and (_12594_, _12593_, _10926_);
  or (_12595_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_12596_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_12597_, _12596_, _12595_);
  and (_12598_, _12597_, _04832_);
  or (_12599_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_12600_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_12601_, _12600_, _12599_);
  and (_12602_, _12601_, _10928_);
  or (_12603_, _12602_, _12598_);
  and (_12604_, _12603_, _04868_);
  or (_12605_, _12604_, _12594_);
  and (_12606_, _12605_, _04859_);
  and (_12607_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_12608_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_12609_, _12608_, _12607_);
  and (_12610_, _12609_, _04832_);
  and (_12611_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_12612_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_12613_, _12612_, _12611_);
  and (_12614_, _12613_, _10928_);
  or (_12615_, _12614_, _12610_);
  and (_12616_, _12615_, _10926_);
  and (_12617_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_12618_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_12619_, _12618_, _12617_);
  and (_12620_, _12619_, _04832_);
  and (_12622_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_12623_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_12624_, _12623_, _12622_);
  and (_12625_, _12624_, _10928_);
  or (_12626_, _12625_, _12620_);
  and (_12627_, _12626_, _04868_);
  or (_12628_, _12627_, _12616_);
  and (_12629_, _12628_, _10945_);
  or (_12630_, _12629_, _12606_);
  and (_12631_, _12630_, _04849_);
  or (_12632_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_12633_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_12634_, _12633_, _10928_);
  and (_12635_, _12634_, _12632_);
  or (_12636_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_12637_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_12638_, _12637_, _04832_);
  and (_12639_, _12638_, _12636_);
  or (_12640_, _12639_, _12635_);
  and (_12641_, _12640_, _10926_);
  or (_12642_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_12643_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_12644_, _12643_, _10928_);
  and (_12645_, _12644_, _12642_);
  or (_12646_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_12647_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_12648_, _12647_, _04832_);
  and (_12649_, _12648_, _12646_);
  or (_12650_, _12649_, _12645_);
  and (_12651_, _12650_, _04868_);
  or (_12652_, _12651_, _12641_);
  and (_12653_, _12652_, _04859_);
  and (_12654_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_12655_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_12656_, _12655_, _12654_);
  and (_12657_, _12656_, _04832_);
  and (_12658_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_12659_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_12660_, _12659_, _12658_);
  and (_12661_, _12660_, _10928_);
  or (_12662_, _12661_, _12657_);
  and (_12663_, _12662_, _10926_);
  and (_12664_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_12665_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_12666_, _12665_, _12664_);
  and (_12667_, _12666_, _04832_);
  and (_12668_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_12669_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_12670_, _12669_, _12668_);
  and (_12671_, _12670_, _10928_);
  or (_12672_, _12671_, _12667_);
  and (_12673_, _12672_, _04868_);
  or (_12674_, _12673_, _12663_);
  and (_12675_, _12674_, _10945_);
  or (_12676_, _12675_, _12653_);
  and (_12677_, _12676_, _10997_);
  or (_12678_, _12677_, _12631_);
  and (_12679_, _12678_, _04839_);
  or (_12680_, _12679_, _12584_);
  or (_12681_, _12680_, _11204_);
  and (_12682_, _12681_, _12490_);
  or (_12683_, _12682_, _03196_);
  and (_12684_, _12683_, _12286_);
  or (_12685_, _12684_, _04876_);
  or (_12686_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_12687_, _12686_, _22773_);
  and (_27321_[1], _12687_, _12685_);
  and (_12688_, _10669_, _24274_);
  not (_12689_, _12688_);
  and (_12690_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nor (_12691_, _12689_, _24026_);
  or (_05829_, _12691_, _12690_);
  and (_12692_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  nor (_12693_, _12689_, _23982_);
  or (_26945_, _12693_, _12692_);
  and (_12694_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  and (_12695_, _03157_, _23900_);
  or (_27159_, _12695_, _12694_);
  and (_12696_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  and (_12697_, _09603_, _23900_);
  or (_05839_, _12697_, _12696_);
  and (_12698_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  and (_12699_, _03157_, _23715_);
  or (_05843_, _12699_, _12698_);
  and (_12700_, _10341_, _24027_);
  and (_12701_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_05845_, _12701_, _12700_);
  and (_12702_, _24061_, _23706_);
  and (_12703_, _12702_, _23920_);
  not (_12704_, _12702_);
  and (_12705_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or (_05848_, _12705_, _12703_);
  and (_12706_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  and (_12707_, _03157_, _23693_);
  or (_05852_, _12707_, _12706_);
  and (_12708_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_12709_, _09722_, _23920_);
  or (_05855_, _12709_, _12708_);
  and (_12710_, _10341_, _23920_);
  and (_12711_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_05857_, _12711_, _12710_);
  and (_12712_, _10341_, _23900_);
  and (_12713_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_05861_, _12713_, _12712_);
  and (_12714_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_12715_, _09722_, _24053_);
  or (_05865_, _12715_, _12714_);
  and (_12716_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  and (_12717_, _09647_, _24027_);
  or (_26958_, _12717_, _12716_);
  and (_12718_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  and (_12719_, _10799_, _24052_);
  or (_05875_, _12719_, _12718_);
  and (_12720_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  and (_12721_, _09647_, _23751_);
  or (_05879_, _12721_, _12720_);
  and (_12722_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  and (_12723_, _09620_, _23983_);
  or (_05884_, _12723_, _12722_);
  and (_12724_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and (_12725_, _10799_, _23692_);
  or (_05892_, _12725_, _12724_);
  and (_12726_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  and (_12727_, _09620_, _23693_);
  or (_05899_, _12727_, _12726_);
  and (_12728_, _25165_, _23920_);
  and (_12729_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_05901_, _12729_, _12728_);
  and (_12730_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and (_12731_, _10799_, _23750_);
  or (_05903_, _12731_, _12730_);
  and (_12732_, _02727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_12733_, _02726_, _24053_);
  or (_05905_, _12733_, _12732_);
  and (_12734_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_12735_, _09597_, _23715_);
  or (_26961_, _12735_, _12734_);
  and (_12736_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_12737_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_12738_, _12737_, _12736_);
  and (_12739_, _12738_, _04832_);
  and (_12740_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_12741_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_12742_, _12741_, _12740_);
  and (_12743_, _12742_, _10928_);
  or (_12744_, _12743_, _12739_);
  or (_12745_, _12744_, _10926_);
  and (_12746_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_12747_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_12748_, _12747_, _12746_);
  and (_12749_, _12748_, _04832_);
  and (_12750_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and (_12751_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_12752_, _12751_, _12750_);
  and (_12753_, _12752_, _10928_);
  or (_12754_, _12753_, _12749_);
  or (_12755_, _12754_, _04868_);
  and (_12756_, _12755_, _10945_);
  and (_12757_, _12756_, _12745_);
  or (_12758_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_12760_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_12761_, _12760_, _12758_);
  and (_12762_, _12761_, _04832_);
  or (_12763_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_12764_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and (_12765_, _12764_, _12763_);
  and (_12766_, _12765_, _10928_);
  or (_12767_, _12766_, _12762_);
  or (_12768_, _12767_, _10926_);
  or (_12769_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_12770_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_12771_, _12770_, _12769_);
  and (_12772_, _12771_, _04832_);
  or (_12773_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_12774_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_12775_, _12774_, _12773_);
  and (_12776_, _12775_, _10928_);
  or (_12777_, _12776_, _12772_);
  or (_12778_, _12777_, _04868_);
  and (_12779_, _12778_, _04859_);
  and (_12780_, _12779_, _12768_);
  or (_12781_, _12780_, _12757_);
  and (_12782_, _12781_, _04849_);
  and (_12783_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_12784_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_12785_, _12784_, _12783_);
  and (_12786_, _12785_, _04832_);
  and (_12787_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and (_12788_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_12789_, _12788_, _12787_);
  and (_12790_, _12789_, _10928_);
  or (_12791_, _12790_, _12786_);
  or (_12792_, _12791_, _10926_);
  and (_12793_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_12794_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_12795_, _12794_, _12793_);
  and (_12796_, _12795_, _04832_);
  and (_12797_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_12798_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_12799_, _12798_, _12797_);
  and (_12800_, _12799_, _10928_);
  or (_12801_, _12800_, _12796_);
  or (_12802_, _12801_, _04868_);
  and (_12803_, _12802_, _10945_);
  and (_12804_, _12803_, _12792_);
  or (_12805_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_12806_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_12807_, _12806_, _10928_);
  and (_12808_, _12807_, _12805_);
  or (_12809_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_12810_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_12811_, _12810_, _04832_);
  and (_12812_, _12811_, _12809_);
  or (_12813_, _12812_, _12808_);
  or (_12814_, _12813_, _10926_);
  or (_12815_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_12816_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_12817_, _12816_, _10928_);
  and (_12818_, _12817_, _12815_);
  or (_12819_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_12820_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and (_12821_, _12820_, _04832_);
  and (_12822_, _12821_, _12819_);
  or (_12823_, _12822_, _12818_);
  or (_12824_, _12823_, _04868_);
  and (_12825_, _12824_, _04859_);
  and (_12826_, _12825_, _12814_);
  or (_12827_, _12826_, _12804_);
  and (_12828_, _12827_, _10997_);
  or (_12829_, _12828_, _12782_);
  and (_12830_, _12829_, _10996_);
  and (_12831_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_12832_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_12833_, _12832_, _12831_);
  and (_12834_, _12833_, _04832_);
  and (_12835_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_12836_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_12837_, _12836_, _12835_);
  and (_12838_, _12837_, _10928_);
  or (_12839_, _12838_, _12834_);
  and (_12840_, _12839_, _04868_);
  and (_12841_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_12842_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_12843_, _12842_, _12841_);
  and (_12844_, _12843_, _04832_);
  and (_12845_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_12846_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_12847_, _12846_, _12845_);
  and (_12848_, _12847_, _10928_);
  or (_12849_, _12848_, _12844_);
  and (_12850_, _12849_, _10926_);
  or (_12851_, _12850_, _12840_);
  and (_12852_, _12851_, _10945_);
  or (_12853_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_12854_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_12855_, _12854_, _10928_);
  and (_12856_, _12855_, _12853_);
  or (_12857_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_12858_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_12859_, _12858_, _04832_);
  and (_12860_, _12859_, _12857_);
  or (_12861_, _12860_, _12856_);
  and (_12862_, _12861_, _04868_);
  or (_12863_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_12864_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_12865_, _12864_, _10928_);
  and (_12866_, _12865_, _12863_);
  or (_12867_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_12868_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_12869_, _12868_, _04832_);
  and (_12870_, _12869_, _12867_);
  or (_12871_, _12870_, _12866_);
  and (_12872_, _12871_, _10926_);
  or (_12873_, _12872_, _12862_);
  and (_12874_, _12873_, _04859_);
  or (_12875_, _12874_, _12852_);
  and (_12876_, _12875_, _10997_);
  and (_12877_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_12878_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_12879_, _12878_, _12877_);
  and (_12880_, _12879_, _04832_);
  and (_12881_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_12882_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_12883_, _12882_, _12881_);
  and (_12884_, _12883_, _10928_);
  or (_12885_, _12884_, _12880_);
  and (_12886_, _12885_, _04868_);
  and (_12887_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_12888_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_12889_, _12888_, _12887_);
  and (_12890_, _12889_, _04832_);
  and (_12891_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_12892_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_12893_, _12892_, _12891_);
  and (_12894_, _12893_, _10928_);
  or (_12895_, _12894_, _12890_);
  and (_12896_, _12895_, _10926_);
  or (_12897_, _12896_, _12886_);
  and (_12898_, _12897_, _10945_);
  or (_12899_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_12900_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_12901_, _12900_, _12899_);
  and (_12902_, _12901_, _04832_);
  or (_12903_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_12904_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_12905_, _12904_, _12903_);
  and (_12906_, _12905_, _10928_);
  or (_12907_, _12906_, _12902_);
  and (_12908_, _12907_, _04868_);
  or (_12909_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_12911_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_12912_, _12911_, _12909_);
  and (_12913_, _12912_, _04832_);
  or (_12914_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_12915_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_12916_, _12915_, _12914_);
  and (_12917_, _12916_, _10928_);
  or (_12918_, _12917_, _12913_);
  and (_12919_, _12918_, _10926_);
  or (_12920_, _12919_, _12908_);
  and (_12921_, _12920_, _04859_);
  or (_12922_, _12921_, _12898_);
  and (_12923_, _12922_, _04849_);
  or (_12924_, _12923_, _12876_);
  and (_12925_, _12924_, _04839_);
  or (_12926_, _12925_, _12830_);
  or (_12927_, _12926_, _04843_);
  and (_12928_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and (_12929_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_12930_, _12929_, _12928_);
  and (_12931_, _12930_, _04832_);
  and (_12932_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_12933_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_12934_, _12933_, _12932_);
  and (_12935_, _12934_, _10928_);
  or (_12936_, _12935_, _12931_);
  or (_12937_, _12936_, _10926_);
  and (_12938_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_12939_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_12940_, _12939_, _12938_);
  and (_12941_, _12940_, _04832_);
  and (_12942_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_12943_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_12944_, _12943_, _12942_);
  and (_12945_, _12944_, _10928_);
  or (_12946_, _12945_, _12941_);
  or (_12947_, _12946_, _04868_);
  and (_12948_, _12947_, _10945_);
  and (_12949_, _12948_, _12937_);
  or (_12950_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_12951_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_12952_, _12951_, _10928_);
  and (_12953_, _12952_, _12950_);
  or (_12954_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_12955_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_12956_, _12955_, _04832_);
  and (_12957_, _12956_, _12954_);
  or (_12958_, _12957_, _12953_);
  or (_12959_, _12958_, _10926_);
  or (_12960_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_12961_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_12962_, _12961_, _10928_);
  and (_12963_, _12962_, _12960_);
  or (_12964_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_12965_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and (_12966_, _12965_, _04832_);
  and (_12967_, _12966_, _12964_);
  or (_12968_, _12967_, _12963_);
  or (_12969_, _12968_, _04868_);
  and (_12970_, _12969_, _04859_);
  and (_12971_, _12970_, _12959_);
  or (_12972_, _12971_, _12949_);
  and (_12973_, _12972_, _10997_);
  and (_12974_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_12975_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_12976_, _12975_, _12974_);
  and (_12977_, _12976_, _04832_);
  and (_12978_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_12979_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_12980_, _12979_, _12978_);
  and (_12981_, _12980_, _10928_);
  or (_12982_, _12981_, _12977_);
  or (_12983_, _12982_, _10926_);
  and (_12984_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_12985_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_12986_, _12985_, _12984_);
  and (_12987_, _12986_, _04832_);
  and (_12988_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_12989_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_12990_, _12989_, _12988_);
  and (_12991_, _12990_, _10928_);
  or (_12992_, _12991_, _12987_);
  or (_12993_, _12992_, _04868_);
  and (_12994_, _12993_, _10945_);
  and (_12995_, _12994_, _12983_);
  or (_12996_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_12997_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_12998_, _12997_, _12996_);
  and (_12999_, _12998_, _04832_);
  or (_13000_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_13001_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_13002_, _13001_, _13000_);
  and (_13003_, _13002_, _10928_);
  or (_13004_, _13003_, _12999_);
  or (_13005_, _13004_, _10926_);
  or (_13006_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_13007_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_13008_, _13007_, _13006_);
  and (_13009_, _13008_, _04832_);
  or (_13010_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_13011_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_13012_, _13011_, _13010_);
  and (_13013_, _13012_, _10928_);
  or (_13014_, _13013_, _13009_);
  or (_13015_, _13014_, _04868_);
  and (_13016_, _13015_, _04859_);
  and (_13017_, _13016_, _13005_);
  or (_13018_, _13017_, _12995_);
  and (_13019_, _13018_, _04849_);
  or (_13020_, _13019_, _12973_);
  and (_13021_, _13020_, _10996_);
  or (_13022_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_13023_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and (_13024_, _13023_, _13022_);
  and (_13025_, _13024_, _04832_);
  or (_13026_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_13027_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_13028_, _13027_, _13026_);
  and (_13029_, _13028_, _10928_);
  or (_13030_, _13029_, _13025_);
  and (_13031_, _13030_, _10926_);
  or (_13032_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_13033_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_13034_, _13033_, _13032_);
  and (_13035_, _13034_, _04832_);
  or (_13036_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_13037_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and (_13038_, _13037_, _13036_);
  and (_13039_, _13038_, _10928_);
  or (_13040_, _13039_, _13035_);
  and (_13041_, _13040_, _04868_);
  or (_13042_, _13041_, _13031_);
  and (_13043_, _13042_, _04859_);
  and (_13044_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_13045_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_13046_, _13045_, _13044_);
  and (_13047_, _13046_, _04832_);
  and (_13048_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_13049_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_13050_, _13049_, _13048_);
  and (_13051_, _13050_, _10928_);
  or (_13052_, _13051_, _13047_);
  and (_13053_, _13052_, _10926_);
  and (_13054_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_13055_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_13056_, _13055_, _13054_);
  and (_13057_, _13056_, _04832_);
  and (_13058_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_13059_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_13060_, _13059_, _13058_);
  and (_13061_, _13060_, _10928_);
  or (_13062_, _13061_, _13057_);
  and (_13063_, _13062_, _04868_);
  or (_13064_, _13063_, _13053_);
  and (_13065_, _13064_, _10945_);
  or (_13066_, _13065_, _13043_);
  and (_13067_, _13066_, _04849_);
  or (_13068_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_13069_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and (_13070_, _13069_, _10928_);
  and (_13071_, _13070_, _13068_);
  or (_13072_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_13073_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and (_13074_, _13073_, _04832_);
  and (_13075_, _13074_, _13072_);
  or (_13076_, _13075_, _13071_);
  and (_13077_, _13076_, _10926_);
  or (_13078_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_13079_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and (_13080_, _13079_, _10928_);
  and (_13081_, _13080_, _13078_);
  or (_13082_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_13083_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and (_13084_, _13083_, _04832_);
  and (_13085_, _13084_, _13082_);
  or (_13086_, _13085_, _13081_);
  and (_13087_, _13086_, _04868_);
  or (_13088_, _13087_, _13077_);
  and (_13089_, _13088_, _04859_);
  and (_13090_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and (_13091_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_13092_, _13091_, _13090_);
  and (_13093_, _13092_, _04832_);
  and (_13094_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and (_13095_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_13096_, _13095_, _13094_);
  and (_13097_, _13096_, _10928_);
  or (_13098_, _13097_, _13093_);
  and (_13099_, _13098_, _10926_);
  and (_13100_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and (_13101_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_13102_, _13101_, _13100_);
  and (_13103_, _13102_, _04832_);
  and (_13104_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and (_13105_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_13106_, _13105_, _13104_);
  and (_13107_, _13106_, _10928_);
  or (_13108_, _13107_, _13103_);
  and (_13109_, _13108_, _04868_);
  or (_13110_, _13109_, _13099_);
  and (_13111_, _13110_, _10945_);
  or (_13112_, _13111_, _13089_);
  and (_13113_, _13112_, _10997_);
  or (_13114_, _13113_, _13067_);
  and (_13115_, _13114_, _04839_);
  or (_13116_, _13115_, _13021_);
  or (_13117_, _13116_, _11204_);
  and (_13118_, _13117_, _12927_);
  or (_13119_, _13118_, _26153_);
  and (_13120_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_13121_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_13122_, _13121_, _13120_);
  and (_13123_, _13122_, _04832_);
  and (_13124_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_13125_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_13126_, _13125_, _13124_);
  and (_13127_, _13126_, _10928_);
  or (_13128_, _13127_, _13123_);
  or (_13129_, _13128_, _10926_);
  and (_13130_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_13131_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_13132_, _13131_, _13130_);
  and (_13133_, _13132_, _04832_);
  and (_13134_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_13135_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_13136_, _13135_, _13134_);
  and (_13137_, _13136_, _10928_);
  or (_13138_, _13137_, _13133_);
  or (_13139_, _13138_, _04868_);
  and (_13140_, _13139_, _10945_);
  and (_13141_, _13140_, _13129_);
  or (_13142_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_13143_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_13144_, _13143_, _13142_);
  and (_13145_, _13144_, _04832_);
  or (_13146_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_13147_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_13148_, _13147_, _13146_);
  and (_13149_, _13148_, _10928_);
  or (_13150_, _13149_, _13145_);
  or (_13151_, _13150_, _10926_);
  or (_13152_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_13153_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_13154_, _13153_, _13152_);
  and (_13155_, _13154_, _04832_);
  or (_13156_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_13157_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_13158_, _13157_, _13156_);
  and (_13159_, _13158_, _10928_);
  or (_13160_, _13159_, _13155_);
  or (_13161_, _13160_, _04868_);
  and (_13162_, _13161_, _04859_);
  and (_13163_, _13162_, _13151_);
  or (_13164_, _13163_, _13141_);
  and (_13165_, _13164_, _04849_);
  and (_13166_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_13167_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_13168_, _13167_, _13166_);
  and (_13169_, _13168_, _04832_);
  and (_13170_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_13171_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_13172_, _13171_, _13170_);
  and (_13173_, _13172_, _10928_);
  or (_13174_, _13173_, _13169_);
  or (_13175_, _13174_, _10926_);
  and (_13176_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_13177_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_13178_, _13177_, _13176_);
  and (_13179_, _13178_, _04832_);
  and (_13180_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_13181_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_13182_, _13181_, _13180_);
  and (_13183_, _13182_, _10928_);
  or (_13184_, _13183_, _13179_);
  or (_13185_, _13184_, _04868_);
  and (_13186_, _13185_, _10945_);
  and (_13187_, _13186_, _13175_);
  or (_13188_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_13189_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_13190_, _13189_, _10928_);
  and (_13191_, _13190_, _13188_);
  or (_13192_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_13193_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_13194_, _13193_, _04832_);
  and (_13195_, _13194_, _13192_);
  or (_13196_, _13195_, _13191_);
  or (_13197_, _13196_, _10926_);
  or (_13198_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_13199_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_13200_, _13199_, _10928_);
  and (_13201_, _13200_, _13198_);
  or (_13202_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_13203_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_13204_, _13203_, _04832_);
  and (_13205_, _13204_, _13202_);
  or (_13206_, _13205_, _13201_);
  or (_13207_, _13206_, _04868_);
  and (_13208_, _13207_, _04859_);
  and (_13209_, _13208_, _13197_);
  or (_13210_, _13209_, _13187_);
  and (_13211_, _13210_, _10997_);
  or (_13212_, _13211_, _13165_);
  and (_13213_, _13212_, _10996_);
  and (_13214_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_13215_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_13216_, _13215_, _13214_);
  and (_13217_, _13216_, _04832_);
  and (_13218_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_13219_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_13220_, _13219_, _13218_);
  and (_13222_, _13220_, _10928_);
  or (_13223_, _13222_, _13217_);
  and (_13224_, _13223_, _04868_);
  and (_13225_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_13226_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_13227_, _13226_, _13225_);
  and (_13228_, _13227_, _04832_);
  and (_13229_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_13230_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_13231_, _13230_, _13229_);
  and (_13232_, _13231_, _10928_);
  or (_13233_, _13232_, _13228_);
  and (_13234_, _13233_, _10926_);
  or (_13235_, _13234_, _13224_);
  and (_13236_, _13235_, _10945_);
  or (_13237_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_13238_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_13239_, _13238_, _10928_);
  and (_13240_, _13239_, _13237_);
  or (_13241_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_13242_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_13243_, _13242_, _04832_);
  and (_13244_, _13243_, _13241_);
  or (_13245_, _13244_, _13240_);
  and (_13246_, _13245_, _04868_);
  or (_13247_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_13248_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_13249_, _13248_, _10928_);
  and (_13250_, _13249_, _13247_);
  or (_13251_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_13252_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_13253_, _13252_, _04832_);
  and (_13254_, _13253_, _13251_);
  or (_13255_, _13254_, _13250_);
  and (_13256_, _13255_, _10926_);
  or (_13257_, _13256_, _13246_);
  and (_13258_, _13257_, _04859_);
  or (_13259_, _13258_, _13236_);
  and (_13260_, _13259_, _10997_);
  and (_13261_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_13262_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_13263_, _13262_, _13261_);
  and (_13264_, _13263_, _04832_);
  and (_13265_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_13266_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_13267_, _13266_, _13265_);
  and (_13268_, _13267_, _10928_);
  or (_13269_, _13268_, _13264_);
  and (_13270_, _13269_, _04868_);
  and (_13271_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_13272_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_13273_, _13272_, _13271_);
  and (_13274_, _13273_, _04832_);
  and (_13275_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_13276_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_13277_, _13276_, _13275_);
  and (_13278_, _13277_, _10928_);
  or (_13279_, _13278_, _13274_);
  and (_13280_, _13279_, _10926_);
  or (_13281_, _13280_, _13270_);
  and (_13282_, _13281_, _10945_);
  or (_13283_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_13284_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_13285_, _13284_, _13283_);
  and (_13286_, _13285_, _04832_);
  or (_13287_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_13288_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_13289_, _13288_, _13287_);
  and (_13290_, _13289_, _10928_);
  or (_13291_, _13290_, _13286_);
  and (_13292_, _13291_, _04868_);
  or (_13293_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_13294_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_13295_, _13294_, _13293_);
  and (_13296_, _13295_, _04832_);
  or (_13297_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_13298_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_13299_, _13298_, _13297_);
  and (_13300_, _13299_, _10928_);
  or (_13301_, _13300_, _13296_);
  and (_13302_, _13301_, _10926_);
  or (_13303_, _13302_, _13292_);
  and (_13304_, _13303_, _04859_);
  or (_13305_, _13304_, _13282_);
  and (_13306_, _13305_, _04849_);
  or (_13307_, _13306_, _13260_);
  and (_13308_, _13307_, _04839_);
  or (_13309_, _13308_, _13213_);
  or (_13310_, _13309_, _04843_);
  and (_13311_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_13312_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_13313_, _13312_, _13311_);
  and (_13314_, _13313_, _04832_);
  and (_13315_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_13316_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_13317_, _13316_, _13315_);
  and (_13318_, _13317_, _10928_);
  or (_13319_, _13318_, _13314_);
  or (_13320_, _13319_, _10926_);
  and (_13321_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_13322_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_13323_, _13322_, _13321_);
  and (_13324_, _13323_, _04832_);
  and (_13325_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_13326_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_13327_, _13326_, _13325_);
  and (_13328_, _13327_, _10928_);
  or (_13329_, _13328_, _13324_);
  or (_13330_, _13329_, _04868_);
  and (_13331_, _13330_, _10945_);
  and (_13332_, _13331_, _13320_);
  or (_13333_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_13334_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_13335_, _13334_, _10928_);
  and (_13336_, _13335_, _13333_);
  or (_13337_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_13338_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_13339_, _13338_, _04832_);
  and (_13340_, _13339_, _13337_);
  or (_13341_, _13340_, _13336_);
  or (_13342_, _13341_, _10926_);
  or (_13343_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_13344_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_13345_, _13344_, _10928_);
  and (_13346_, _13345_, _13343_);
  or (_13347_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_13348_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_13349_, _13348_, _04832_);
  and (_13350_, _13349_, _13347_);
  or (_13351_, _13350_, _13346_);
  or (_13352_, _13351_, _04868_);
  and (_13353_, _13352_, _04859_);
  and (_13354_, _13353_, _13342_);
  or (_13355_, _13354_, _13332_);
  and (_13356_, _13355_, _10997_);
  and (_13357_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_13358_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_13359_, _13358_, _13357_);
  and (_13360_, _13359_, _04832_);
  and (_13361_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_13362_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_13363_, _13362_, _13361_);
  and (_13364_, _13363_, _10928_);
  or (_13365_, _13364_, _13360_);
  or (_13366_, _13365_, _10926_);
  and (_13367_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_13368_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_13369_, _13368_, _13367_);
  and (_13370_, _13369_, _04832_);
  and (_13371_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_13372_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_13373_, _13372_, _13371_);
  and (_13374_, _13373_, _10928_);
  or (_13375_, _13374_, _13370_);
  or (_13376_, _13375_, _04868_);
  and (_13377_, _13376_, _10945_);
  and (_13378_, _13377_, _13366_);
  or (_13379_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_13380_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_13381_, _13380_, _13379_);
  and (_13382_, _13381_, _04832_);
  or (_13383_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_13384_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_13385_, _13384_, _13383_);
  and (_13386_, _13385_, _10928_);
  or (_13387_, _13386_, _13382_);
  or (_13388_, _13387_, _10926_);
  or (_13389_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_13390_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_13391_, _13390_, _13389_);
  and (_13392_, _13391_, _04832_);
  or (_13393_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_13394_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_13395_, _13394_, _13393_);
  and (_13396_, _13395_, _10928_);
  or (_13397_, _13396_, _13392_);
  or (_13398_, _13397_, _04868_);
  and (_13399_, _13398_, _04859_);
  and (_13400_, _13399_, _13388_);
  or (_13401_, _13400_, _13378_);
  and (_13402_, _13401_, _04849_);
  or (_13403_, _13402_, _13356_);
  and (_13404_, _13403_, _10996_);
  or (_13405_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_13406_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_13407_, _13406_, _13405_);
  and (_13408_, _13407_, _04832_);
  or (_13409_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_13410_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_13411_, _13410_, _13409_);
  and (_13412_, _13411_, _10928_);
  or (_13413_, _13412_, _13408_);
  and (_13414_, _13413_, _10926_);
  or (_13415_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_13416_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_13417_, _13416_, _13415_);
  and (_13418_, _13417_, _04832_);
  or (_13419_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_13420_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_13421_, _13420_, _13419_);
  and (_13422_, _13421_, _10928_);
  or (_13423_, _13422_, _13418_);
  and (_13424_, _13423_, _04868_);
  or (_13425_, _13424_, _13414_);
  and (_13426_, _13425_, _04859_);
  and (_13427_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_13428_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_13429_, _13428_, _13427_);
  and (_13430_, _13429_, _04832_);
  and (_13431_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_13432_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_13433_, _13432_, _13431_);
  and (_13434_, _13433_, _10928_);
  or (_13435_, _13434_, _13430_);
  and (_13436_, _13435_, _10926_);
  and (_13437_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_13438_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_13439_, _13438_, _13437_);
  and (_13440_, _13439_, _04832_);
  and (_13441_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_13442_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_13443_, _13442_, _13441_);
  and (_13444_, _13443_, _10928_);
  or (_13445_, _13444_, _13440_);
  and (_13446_, _13445_, _04868_);
  or (_13447_, _13446_, _13436_);
  and (_13448_, _13447_, _10945_);
  or (_13449_, _13448_, _13426_);
  and (_13450_, _13449_, _04849_);
  or (_13451_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_13452_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_13453_, _13452_, _10928_);
  and (_13454_, _13453_, _13451_);
  or (_13455_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_13456_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_13457_, _13456_, _04832_);
  and (_13458_, _13457_, _13455_);
  or (_13459_, _13458_, _13454_);
  and (_13460_, _13459_, _10926_);
  or (_13461_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_13462_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_13463_, _13462_, _10928_);
  and (_13464_, _13463_, _13461_);
  or (_13465_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_13466_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_13467_, _13466_, _04832_);
  and (_13468_, _13467_, _13465_);
  or (_13469_, _13468_, _13464_);
  and (_13470_, _13469_, _04868_);
  or (_13471_, _13470_, _13460_);
  and (_13472_, _13471_, _04859_);
  and (_13473_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_13474_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_13475_, _13474_, _13473_);
  and (_13476_, _13475_, _04832_);
  and (_13477_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_13478_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_13479_, _13478_, _13477_);
  and (_13480_, _13479_, _10928_);
  or (_13481_, _13480_, _13476_);
  and (_13482_, _13481_, _10926_);
  and (_13483_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_13484_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_13485_, _13484_, _13483_);
  and (_13486_, _13485_, _04832_);
  and (_13487_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_13488_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_13489_, _13488_, _13487_);
  and (_13490_, _13489_, _10928_);
  or (_13491_, _13490_, _13486_);
  and (_13492_, _13491_, _04868_);
  or (_13493_, _13492_, _13482_);
  and (_13494_, _13493_, _10945_);
  or (_13495_, _13494_, _13472_);
  and (_13496_, _13495_, _10997_);
  or (_13497_, _13496_, _13450_);
  and (_13498_, _13497_, _04839_);
  or (_13499_, _13498_, _13404_);
  or (_13500_, _13499_, _11204_);
  and (_13501_, _13500_, _13310_);
  or (_13502_, _13501_, _03196_);
  and (_13503_, _13502_, _13119_);
  or (_13504_, _13503_, _04876_);
  or (_13505_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_13506_, _13505_, _22773_);
  and (_05907_, _13506_, _13504_);
  and (_13507_, _09463_, _23920_);
  and (_13508_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_27055_, _13508_, _13507_);
  and (_13509_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_13510_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_13511_, _13510_, _13509_);
  and (_13512_, _13511_, _10928_);
  and (_13513_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_13514_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_13515_, _13514_, _13513_);
  and (_13516_, _13515_, _04832_);
  or (_13517_, _13516_, _13512_);
  or (_13518_, _13517_, _10926_);
  and (_13519_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_13521_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_13522_, _13521_, _13519_);
  and (_13523_, _13522_, _10928_);
  and (_13524_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_13525_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_13526_, _13525_, _13524_);
  and (_13527_, _13526_, _04832_);
  or (_13528_, _13527_, _13523_);
  or (_13529_, _13528_, _04868_);
  and (_13530_, _13529_, _10945_);
  and (_13531_, _13530_, _13518_);
  or (_13532_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_13533_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_13534_, _13533_, _04832_);
  and (_13535_, _13534_, _13532_);
  or (_13536_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_13537_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and (_13538_, _13537_, _10928_);
  and (_13539_, _13538_, _13536_);
  or (_13540_, _13539_, _13535_);
  or (_13541_, _13540_, _10926_);
  or (_13542_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_13543_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_13544_, _13543_, _04832_);
  and (_13545_, _13544_, _13542_);
  or (_13546_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_13547_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and (_13548_, _13547_, _10928_);
  and (_13549_, _13548_, _13546_);
  or (_13550_, _13549_, _13545_);
  or (_13551_, _13550_, _04868_);
  and (_13552_, _13551_, _04859_);
  and (_13553_, _13552_, _13541_);
  or (_13554_, _13553_, _13531_);
  or (_13555_, _13554_, _04849_);
  and (_13556_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_13557_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_13558_, _13557_, _04832_);
  or (_13559_, _13558_, _13556_);
  and (_13560_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_13561_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_13562_, _13561_, _10928_);
  or (_13563_, _13562_, _13560_);
  and (_13564_, _13563_, _13559_);
  or (_13565_, _13564_, _10926_);
  and (_13566_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and (_13567_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_13568_, _13567_, _04832_);
  or (_13569_, _13568_, _13566_);
  and (_13570_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_13571_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_13572_, _13571_, _10928_);
  or (_13573_, _13572_, _13570_);
  and (_13574_, _13573_, _13569_);
  or (_13575_, _13574_, _04868_);
  and (_13576_, _13575_, _10945_);
  and (_13577_, _13576_, _13565_);
  or (_13578_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_13579_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_13580_, _13579_, _13578_);
  or (_13581_, _13580_, _10928_);
  or (_13582_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_13583_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_13584_, _13583_, _13582_);
  or (_13585_, _13584_, _04832_);
  and (_13586_, _13585_, _13581_);
  or (_13587_, _13586_, _10926_);
  or (_13588_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_13589_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_13590_, _13589_, _13588_);
  or (_13591_, _13590_, _10928_);
  or (_13592_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_13593_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_13594_, _13593_, _13592_);
  or (_13595_, _13594_, _04832_);
  and (_13596_, _13595_, _13591_);
  or (_13597_, _13596_, _04868_);
  and (_13598_, _13597_, _04859_);
  and (_13599_, _13598_, _13587_);
  or (_13600_, _13599_, _13577_);
  or (_13602_, _13600_, _10997_);
  and (_13603_, _13602_, _10996_);
  and (_13604_, _13603_, _13555_);
  and (_13605_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_13606_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_13607_, _13606_, _13605_);
  and (_13608_, _13607_, _04832_);
  and (_13609_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_13610_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_13611_, _13610_, _13609_);
  and (_13612_, _13611_, _10928_);
  or (_13613_, _13612_, _13608_);
  and (_13614_, _13613_, _04868_);
  and (_13615_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_13616_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_13617_, _13616_, _13615_);
  and (_13618_, _13617_, _04832_);
  and (_13619_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_13620_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_13621_, _13620_, _13619_);
  and (_13622_, _13621_, _10928_);
  or (_13623_, _13622_, _13618_);
  and (_13624_, _13623_, _10926_);
  or (_13625_, _13624_, _13614_);
  and (_13626_, _13625_, _10945_);
  or (_13627_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_13628_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_13629_, _13628_, _13627_);
  and (_13630_, _13629_, _04832_);
  or (_13631_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_13632_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_13633_, _13632_, _13631_);
  and (_13634_, _13633_, _10928_);
  or (_13635_, _13634_, _13630_);
  and (_13636_, _13635_, _04868_);
  or (_13637_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_13638_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_13639_, _13638_, _13637_);
  and (_13640_, _13639_, _04832_);
  or (_13641_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_13642_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_13643_, _13642_, _13641_);
  and (_13644_, _13643_, _10928_);
  or (_13645_, _13644_, _13640_);
  and (_13646_, _13645_, _10926_);
  or (_13647_, _13646_, _13636_);
  and (_13648_, _13647_, _04859_);
  or (_13649_, _13648_, _13626_);
  and (_13650_, _13649_, _10997_);
  and (_13651_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_13652_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_13653_, _13652_, _13651_);
  and (_13654_, _13653_, _04832_);
  and (_13655_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_13656_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_13657_, _13656_, _13655_);
  and (_13658_, _13657_, _10928_);
  or (_13659_, _13658_, _13654_);
  and (_13660_, _13659_, _04868_);
  and (_13661_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_13662_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_13663_, _13662_, _13661_);
  and (_13664_, _13663_, _04832_);
  and (_13665_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and (_13666_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_13667_, _13666_, _13665_);
  and (_13668_, _13667_, _10928_);
  or (_13669_, _13668_, _13664_);
  and (_13670_, _13669_, _10926_);
  or (_13671_, _13670_, _13660_);
  and (_13672_, _13671_, _10945_);
  or (_13673_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_13674_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and (_13675_, _13674_, _13673_);
  and (_13676_, _13675_, _04832_);
  or (_13677_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_13678_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_13679_, _13678_, _13677_);
  and (_13680_, _13679_, _10928_);
  or (_13681_, _13680_, _13676_);
  and (_13682_, _13681_, _04868_);
  or (_13683_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_13684_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and (_13685_, _13684_, _13683_);
  and (_13686_, _13685_, _04832_);
  or (_13687_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_13688_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_13689_, _13688_, _13687_);
  and (_13690_, _13689_, _10928_);
  or (_13691_, _13690_, _13686_);
  and (_13692_, _13691_, _10926_);
  or (_13693_, _13692_, _13682_);
  and (_13694_, _13693_, _04859_);
  or (_13695_, _13694_, _13672_);
  and (_13696_, _13695_, _04849_);
  or (_13697_, _13696_, _13650_);
  and (_13698_, _13697_, _04839_);
  or (_13699_, _13698_, _13604_);
  or (_13700_, _13699_, _04843_);
  and (_13701_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_13702_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_13703_, _13702_, _13701_);
  and (_13704_, _13703_, _04832_);
  and (_13705_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_13706_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_13707_, _13706_, _13705_);
  and (_13708_, _13707_, _10928_);
  or (_13709_, _13708_, _13704_);
  or (_13710_, _13709_, _10926_);
  and (_13711_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_13712_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_13713_, _13712_, _13711_);
  and (_13714_, _13713_, _04832_);
  and (_13715_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_13716_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_13717_, _13716_, _13715_);
  and (_13718_, _13717_, _10928_);
  or (_13719_, _13718_, _13714_);
  or (_13720_, _13719_, _04868_);
  and (_13721_, _13720_, _10945_);
  and (_13722_, _13721_, _13710_);
  or (_13723_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_13724_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_13725_, _13724_, _10928_);
  and (_13726_, _13725_, _13723_);
  or (_13727_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_13728_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_13729_, _13728_, _04832_);
  and (_13730_, _13729_, _13727_);
  or (_13731_, _13730_, _13726_);
  or (_13732_, _13731_, _10926_);
  or (_13733_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_13734_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and (_13735_, _13734_, _10928_);
  and (_13736_, _13735_, _13733_);
  or (_13737_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_13738_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and (_13739_, _13738_, _04832_);
  and (_13740_, _13739_, _13737_);
  or (_13741_, _13740_, _13736_);
  or (_13742_, _13741_, _04868_);
  and (_13743_, _13742_, _04859_);
  and (_13744_, _13743_, _13732_);
  or (_13745_, _13744_, _13722_);
  and (_13746_, _13745_, _10997_);
  and (_13747_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_13748_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_13749_, _13748_, _13747_);
  and (_13750_, _13749_, _04832_);
  and (_13751_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_13752_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_13753_, _13752_, _13751_);
  and (_13754_, _13753_, _10928_);
  or (_13755_, _13754_, _13750_);
  or (_13756_, _13755_, _10926_);
  and (_13757_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_13758_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_13759_, _13758_, _13757_);
  and (_13760_, _13759_, _04832_);
  and (_13761_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_13762_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_13763_, _13762_, _13761_);
  and (_13764_, _13763_, _10928_);
  or (_13765_, _13764_, _13760_);
  or (_13766_, _13765_, _04868_);
  and (_13767_, _13766_, _10945_);
  and (_13768_, _13767_, _13756_);
  or (_13769_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_13770_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_13771_, _13770_, _13769_);
  and (_13772_, _13771_, _04832_);
  or (_13773_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_13774_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_13775_, _13774_, _13773_);
  and (_13776_, _13775_, _10928_);
  or (_13777_, _13776_, _13772_);
  or (_13778_, _13777_, _10926_);
  or (_13779_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_13780_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_13781_, _13780_, _13779_);
  and (_13782_, _13781_, _04832_);
  or (_13783_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_13784_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_13785_, _13784_, _13783_);
  and (_13786_, _13785_, _10928_);
  or (_13787_, _13786_, _13782_);
  or (_13788_, _13787_, _04868_);
  and (_13789_, _13788_, _04859_);
  and (_13790_, _13789_, _13778_);
  or (_13791_, _13790_, _13768_);
  and (_13793_, _13791_, _04849_);
  or (_13794_, _13793_, _13746_);
  and (_13795_, _13794_, _10996_);
  or (_13796_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_13797_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and (_13798_, _13797_, _13796_);
  and (_13799_, _13798_, _04832_);
  or (_13800_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_13801_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_13802_, _13801_, _13800_);
  and (_13803_, _13802_, _10928_);
  or (_13804_, _13803_, _13799_);
  and (_13805_, _13804_, _10926_);
  or (_13806_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_13807_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_13808_, _13807_, _13806_);
  and (_13809_, _13808_, _04832_);
  or (_13810_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_13811_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_13812_, _13811_, _13810_);
  and (_13814_, _13812_, _10928_);
  or (_13815_, _13814_, _13809_);
  and (_13816_, _13815_, _04868_);
  or (_13817_, _13816_, _13805_);
  and (_13818_, _13817_, _04859_);
  and (_13819_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and (_13820_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_13821_, _13820_, _13819_);
  and (_13822_, _13821_, _04832_);
  and (_13823_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and (_13824_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_13825_, _13824_, _13823_);
  and (_13826_, _13825_, _10928_);
  or (_13827_, _13826_, _13822_);
  and (_13828_, _13827_, _10926_);
  and (_13829_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and (_13830_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_13831_, _13830_, _13829_);
  and (_13832_, _13831_, _04832_);
  and (_13833_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_13834_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_13835_, _13834_, _13833_);
  and (_13836_, _13835_, _10928_);
  or (_13837_, _13836_, _13832_);
  and (_13838_, _13837_, _04868_);
  or (_13839_, _13838_, _13828_);
  and (_13840_, _13839_, _10945_);
  or (_13841_, _13840_, _13818_);
  and (_13842_, _13841_, _04849_);
  or (_13843_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_13844_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_13845_, _13844_, _10928_);
  and (_13846_, _13845_, _13843_);
  or (_13847_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_13848_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_13849_, _13848_, _04832_);
  and (_13850_, _13849_, _13847_);
  or (_13851_, _13850_, _13846_);
  and (_13852_, _13851_, _10926_);
  or (_13853_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_13854_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_13855_, _13854_, _10928_);
  and (_13856_, _13855_, _13853_);
  or (_13857_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_13858_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and (_13859_, _13858_, _04832_);
  and (_13860_, _13859_, _13857_);
  or (_13861_, _13860_, _13856_);
  and (_13862_, _13861_, _04868_);
  or (_13863_, _13862_, _13852_);
  and (_13865_, _13863_, _04859_);
  and (_13866_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and (_13867_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_13868_, _13867_, _13866_);
  and (_13869_, _13868_, _04832_);
  and (_13870_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_13871_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_13872_, _13871_, _13870_);
  and (_13873_, _13872_, _10928_);
  or (_13874_, _13873_, _13869_);
  and (_13875_, _13874_, _10926_);
  and (_13876_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_13877_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_13878_, _13877_, _13876_);
  and (_13879_, _13878_, _04832_);
  and (_13880_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_13881_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_13882_, _13881_, _13880_);
  and (_13883_, _13882_, _10928_);
  or (_13884_, _13883_, _13879_);
  and (_13886_, _13884_, _04868_);
  or (_13887_, _13886_, _13875_);
  and (_13888_, _13887_, _10945_);
  or (_13889_, _13888_, _13865_);
  and (_13890_, _13889_, _10997_);
  or (_13891_, _13890_, _13842_);
  and (_13892_, _13891_, _04839_);
  or (_13893_, _13892_, _13795_);
  or (_13894_, _13893_, _11204_);
  and (_13895_, _13894_, _13700_);
  or (_13896_, _13895_, _26153_);
  and (_13897_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_13898_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_13899_, _13898_, _13897_);
  and (_13900_, _13899_, _04832_);
  and (_13901_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_13902_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_13903_, _13902_, _13901_);
  and (_13904_, _13903_, _10928_);
  or (_13905_, _13904_, _13900_);
  and (_13906_, _13905_, _04868_);
  and (_13907_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_13908_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_13909_, _13908_, _13907_);
  and (_13910_, _13909_, _04832_);
  and (_13911_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_13912_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_13913_, _13912_, _13911_);
  and (_13914_, _13913_, _10928_);
  or (_13915_, _13914_, _13910_);
  and (_13916_, _13915_, _10926_);
  or (_13917_, _13916_, _13906_);
  and (_13918_, _13917_, _10945_);
  or (_13919_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_13920_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_13921_, _13920_, _10928_);
  and (_13922_, _13921_, _13919_);
  or (_13923_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_13924_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_13925_, _13924_, _04832_);
  and (_13926_, _13925_, _13923_);
  or (_13927_, _13926_, _13922_);
  and (_13928_, _13927_, _04868_);
  or (_13929_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_13930_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_13931_, _13930_, _10928_);
  and (_13932_, _13931_, _13929_);
  or (_13933_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_13934_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_13935_, _13934_, _04832_);
  and (_13936_, _13935_, _13933_);
  or (_13937_, _13936_, _13932_);
  and (_13938_, _13937_, _10926_);
  or (_13939_, _13938_, _13928_);
  and (_13940_, _13939_, _04859_);
  or (_13941_, _13940_, _13918_);
  and (_13942_, _13941_, _10997_);
  and (_13943_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_13944_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_13945_, _13944_, _13943_);
  and (_13946_, _13945_, _04832_);
  and (_13947_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_13948_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_13949_, _13948_, _13947_);
  and (_13950_, _13949_, _10928_);
  or (_13951_, _13950_, _13946_);
  and (_13952_, _13951_, _04868_);
  and (_13953_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_13954_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_13955_, _13954_, _13953_);
  and (_13956_, _13955_, _04832_);
  and (_13957_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_13958_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_13959_, _13958_, _13957_);
  and (_13960_, _13959_, _10928_);
  or (_13961_, _13960_, _13956_);
  and (_13962_, _13961_, _10926_);
  or (_13963_, _13962_, _13952_);
  and (_13964_, _13963_, _10945_);
  or (_13965_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_13966_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_13967_, _13966_, _13965_);
  and (_13968_, _13967_, _04832_);
  or (_13969_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_13970_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_13971_, _13970_, _13969_);
  and (_13972_, _13971_, _10928_);
  or (_13973_, _13972_, _13968_);
  and (_13974_, _13973_, _04868_);
  or (_13975_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_13977_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_13978_, _13977_, _13975_);
  and (_13979_, _13978_, _04832_);
  or (_13980_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_13981_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_13982_, _13981_, _13980_);
  and (_13983_, _13982_, _10928_);
  or (_13984_, _13983_, _13979_);
  and (_13985_, _13984_, _10926_);
  or (_13986_, _13985_, _13974_);
  and (_13987_, _13986_, _04859_);
  or (_13988_, _13987_, _13964_);
  and (_13989_, _13988_, _04849_);
  or (_13990_, _13989_, _13942_);
  and (_13991_, _13990_, _04839_);
  and (_13992_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_13993_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_13994_, _13993_, _13992_);
  and (_13995_, _13994_, _04832_);
  and (_13996_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_13997_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_13998_, _13997_, _13996_);
  and (_13999_, _13998_, _10928_);
  or (_14000_, _13999_, _13995_);
  or (_14001_, _14000_, _10926_);
  and (_14002_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_14003_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_14004_, _14003_, _14002_);
  and (_14005_, _14004_, _04832_);
  and (_14006_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_14007_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_14008_, _14007_, _14006_);
  and (_14009_, _14008_, _10928_);
  or (_14010_, _14009_, _14005_);
  or (_14011_, _14010_, _04868_);
  and (_14012_, _14011_, _10945_);
  and (_14013_, _14012_, _14001_);
  or (_14014_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_14015_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_14016_, _14015_, _14014_);
  and (_14017_, _14016_, _04832_);
  or (_14018_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_14019_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_14020_, _14019_, _14018_);
  and (_14021_, _14020_, _10928_);
  or (_14022_, _14021_, _14017_);
  or (_14023_, _14022_, _10926_);
  or (_14024_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_14025_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_14026_, _14025_, _14024_);
  and (_14027_, _14026_, _04832_);
  or (_14028_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_14029_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_14030_, _14029_, _14028_);
  and (_14031_, _14030_, _10928_);
  or (_14032_, _14031_, _14027_);
  or (_14033_, _14032_, _04868_);
  and (_14034_, _14033_, _04859_);
  and (_14035_, _14034_, _14023_);
  or (_14036_, _14035_, _14013_);
  and (_14037_, _14036_, _04849_);
  and (_14038_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_14039_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_14040_, _14039_, _14038_);
  and (_14041_, _14040_, _04832_);
  and (_14042_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_14043_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_14044_, _14043_, _14042_);
  and (_14045_, _14044_, _10928_);
  or (_14046_, _14045_, _14041_);
  or (_14047_, _14046_, _10926_);
  and (_14048_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_14049_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_14050_, _14049_, _14048_);
  and (_14051_, _14050_, _04832_);
  and (_14052_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_14053_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_14054_, _14053_, _14052_);
  and (_14055_, _14054_, _10928_);
  or (_14056_, _14055_, _14051_);
  or (_14058_, _14056_, _04868_);
  and (_14059_, _14058_, _10945_);
  and (_14060_, _14059_, _14047_);
  or (_14061_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_14062_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_14063_, _14062_, _10928_);
  and (_14064_, _14063_, _14061_);
  or (_14065_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_14066_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_14067_, _14066_, _04832_);
  and (_14068_, _14067_, _14065_);
  or (_14069_, _14068_, _14064_);
  or (_14070_, _14069_, _10926_);
  or (_14071_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_14072_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_14073_, _14072_, _10928_);
  and (_14074_, _14073_, _14071_);
  or (_14075_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_14076_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_14077_, _14076_, _04832_);
  and (_14078_, _14077_, _14075_);
  or (_14079_, _14078_, _14074_);
  or (_14080_, _14079_, _04868_);
  and (_14081_, _14080_, _04859_);
  and (_14082_, _14081_, _14070_);
  or (_14083_, _14082_, _14060_);
  and (_14084_, _14083_, _10997_);
  or (_14085_, _14084_, _14037_);
  and (_14086_, _14085_, _10996_);
  or (_14087_, _14086_, _13991_);
  or (_14088_, _14087_, _04843_);
  and (_14089_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_14090_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_14091_, _14090_, _14089_);
  and (_14092_, _14091_, _10928_);
  and (_14093_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_14094_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_14095_, _14094_, _14093_);
  and (_14096_, _14095_, _04832_);
  or (_14097_, _14096_, _14092_);
  or (_14098_, _14097_, _10926_);
  and (_14099_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_14100_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_14101_, _14100_, _14099_);
  and (_14102_, _14101_, _10928_);
  and (_14103_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_14104_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_14105_, _14104_, _14103_);
  and (_14106_, _14105_, _04832_);
  or (_14107_, _14106_, _14102_);
  or (_14108_, _14107_, _04868_);
  and (_14109_, _14108_, _10945_);
  and (_14110_, _14109_, _14098_);
  or (_14111_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_14112_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_14113_, _14112_, _04832_);
  and (_14114_, _14113_, _14111_);
  or (_14115_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_14116_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_14117_, _14116_, _10928_);
  and (_14119_, _14117_, _14115_);
  or (_14120_, _14119_, _14114_);
  or (_14121_, _14120_, _10926_);
  or (_14122_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_14123_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_14124_, _14123_, _04832_);
  and (_14125_, _14124_, _14122_);
  or (_14126_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_14127_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_14128_, _14127_, _10928_);
  and (_14129_, _14128_, _14126_);
  or (_14130_, _14129_, _14125_);
  or (_14131_, _14130_, _04868_);
  and (_14132_, _14131_, _04859_);
  and (_14133_, _14132_, _14121_);
  or (_14134_, _14133_, _14110_);
  and (_14135_, _14134_, _10997_);
  and (_14136_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_14137_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_14138_, _14137_, _04832_);
  or (_14139_, _14138_, _14136_);
  and (_14140_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_14141_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_14142_, _14141_, _10928_);
  or (_14143_, _14142_, _14140_);
  and (_14144_, _14143_, _14139_);
  or (_14145_, _14144_, _10926_);
  and (_14146_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_14147_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_14148_, _14147_, _04832_);
  or (_14149_, _14148_, _14146_);
  and (_14150_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_14151_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_14152_, _14151_, _10928_);
  or (_14153_, _14152_, _14150_);
  and (_14154_, _14153_, _14149_);
  or (_14155_, _14154_, _04868_);
  and (_14156_, _14155_, _10945_);
  and (_14157_, _14156_, _14145_);
  or (_14158_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_14159_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_14160_, _14159_, _14158_);
  or (_14161_, _14160_, _10928_);
  or (_14162_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_14163_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_14164_, _14163_, _14162_);
  or (_14165_, _14164_, _04832_);
  and (_14166_, _14165_, _14161_);
  or (_14167_, _14166_, _10926_);
  or (_14168_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_14169_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_14170_, _14169_, _14168_);
  or (_14171_, _14170_, _10928_);
  or (_14172_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_14173_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_14174_, _14173_, _14172_);
  or (_14175_, _14174_, _04832_);
  and (_14176_, _14175_, _14171_);
  or (_14177_, _14176_, _04868_);
  and (_14178_, _14177_, _04859_);
  and (_14179_, _14178_, _14167_);
  or (_14180_, _14179_, _14157_);
  and (_14181_, _14180_, _04849_);
  or (_14182_, _14181_, _14135_);
  and (_14183_, _14182_, _10996_);
  and (_14184_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_14185_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_14186_, _14185_, _14184_);
  and (_14187_, _14186_, _04832_);
  and (_14188_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_14189_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_14190_, _14189_, _14188_);
  and (_14191_, _14190_, _10928_);
  or (_14192_, _14191_, _14187_);
  and (_14193_, _14192_, _04868_);
  and (_14194_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_14195_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_14196_, _14195_, _14194_);
  and (_14197_, _14196_, _04832_);
  and (_14198_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_14199_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_14200_, _14199_, _14198_);
  and (_14201_, _14200_, _10928_);
  or (_14202_, _14201_, _14197_);
  and (_14203_, _14202_, _10926_);
  or (_14204_, _14203_, _14193_);
  and (_14205_, _14204_, _10945_);
  or (_14206_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_14207_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_14208_, _14207_, _14206_);
  and (_14210_, _14208_, _04832_);
  or (_14211_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_14212_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_14213_, _14212_, _14211_);
  and (_14214_, _14213_, _10928_);
  or (_14215_, _14214_, _14210_);
  and (_14216_, _14215_, _04868_);
  or (_14217_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_14218_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_14219_, _14218_, _14217_);
  and (_14220_, _14219_, _04832_);
  or (_14221_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_14222_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_14223_, _14222_, _14221_);
  and (_14224_, _14223_, _10928_);
  or (_14225_, _14224_, _14220_);
  and (_14226_, _14225_, _10926_);
  or (_14227_, _14226_, _14216_);
  and (_14228_, _14227_, _04859_);
  or (_14229_, _14228_, _14205_);
  and (_14230_, _14229_, _04849_);
  and (_14231_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  and (_14232_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_14233_, _14232_, _14231_);
  and (_14234_, _14233_, _04832_);
  and (_14235_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  and (_14236_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_14237_, _14236_, _14235_);
  and (_14238_, _14237_, _10928_);
  or (_14239_, _14238_, _14234_);
  and (_14240_, _14239_, _04868_);
  and (_14241_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  and (_14242_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_14243_, _14242_, _14241_);
  and (_14244_, _14243_, _04832_);
  and (_14245_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  and (_14246_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_14247_, _14246_, _14245_);
  and (_14248_, _14247_, _10928_);
  or (_14249_, _14248_, _14244_);
  and (_14250_, _14249_, _10926_);
  or (_14251_, _14250_, _14240_);
  and (_14252_, _14251_, _10945_);
  or (_14253_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_14254_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and (_14255_, _14254_, _14253_);
  and (_14256_, _14255_, _04832_);
  or (_14257_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_14258_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  and (_14259_, _14258_, _14257_);
  and (_14260_, _14259_, _10928_);
  or (_14261_, _14260_, _14256_);
  and (_14262_, _14261_, _04868_);
  or (_14263_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_14264_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  and (_14265_, _14264_, _14263_);
  and (_14266_, _14265_, _04832_);
  or (_14267_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_14268_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  and (_14269_, _14268_, _14267_);
  and (_14270_, _14269_, _10928_);
  or (_14271_, _14270_, _14266_);
  and (_14272_, _14271_, _10926_);
  or (_14273_, _14272_, _14262_);
  and (_14274_, _14273_, _04859_);
  or (_14275_, _14274_, _14252_);
  and (_14276_, _14275_, _10997_);
  or (_14277_, _14276_, _14230_);
  and (_14278_, _14277_, _04839_);
  or (_14279_, _14278_, _14183_);
  or (_14280_, _14279_, _11204_);
  and (_14281_, _14280_, _14088_);
  or (_14282_, _14281_, _03196_);
  and (_14283_, _14282_, _13896_);
  or (_14284_, _14283_, _04876_);
  or (_14285_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_14286_, _14285_, _22773_);
  and (_05911_, _14286_, _14284_);
  and (_14287_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_14288_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_14289_, _14288_, _14287_);
  and (_14290_, _14289_, _04832_);
  and (_14291_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_14292_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_14293_, _14292_, _14291_);
  and (_14294_, _14293_, _10928_);
  or (_14295_, _14294_, _14290_);
  or (_14296_, _14295_, _10926_);
  and (_14297_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_14298_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_14299_, _14298_, _14297_);
  and (_14300_, _14299_, _04832_);
  and (_14301_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_14302_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_14303_, _14302_, _14301_);
  and (_14304_, _14303_, _10928_);
  or (_14305_, _14304_, _14300_);
  or (_14306_, _14305_, _04868_);
  and (_14307_, _14306_, _10945_);
  and (_14308_, _14307_, _14296_);
  or (_14309_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_14310_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_14311_, _14310_, _14309_);
  and (_14312_, _14311_, _04832_);
  or (_14313_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_14314_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_14315_, _14314_, _14313_);
  and (_14316_, _14315_, _10928_);
  or (_14317_, _14316_, _14312_);
  or (_14318_, _14317_, _10926_);
  or (_14319_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_14320_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and (_14321_, _14320_, _14319_);
  and (_14322_, _14321_, _04832_);
  or (_14323_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_14324_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_14325_, _14324_, _14323_);
  and (_14326_, _14325_, _10928_);
  or (_14327_, _14326_, _14322_);
  or (_14328_, _14327_, _04868_);
  and (_14329_, _14328_, _04859_);
  and (_14330_, _14329_, _14318_);
  or (_14331_, _14330_, _14308_);
  or (_14332_, _14331_, _10997_);
  and (_14333_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_14334_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_14335_, _14334_, _14333_);
  and (_14336_, _14335_, _04832_);
  and (_14337_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_14338_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_14339_, _14338_, _14337_);
  and (_14340_, _14339_, _10928_);
  or (_14341_, _14340_, _14336_);
  or (_14342_, _14341_, _10926_);
  and (_14343_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_14344_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_14345_, _14344_, _14343_);
  and (_14346_, _14345_, _04832_);
  and (_14347_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_14348_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_14349_, _14348_, _14347_);
  and (_14350_, _14349_, _10928_);
  or (_14351_, _14350_, _14346_);
  or (_14352_, _14351_, _04868_);
  and (_14353_, _14352_, _10945_);
  and (_14354_, _14353_, _14342_);
  or (_14355_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_14356_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_14357_, _14356_, _10928_);
  and (_14358_, _14357_, _14355_);
  or (_14359_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_14360_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_14361_, _14360_, _04832_);
  and (_14362_, _14361_, _14359_);
  or (_14363_, _14362_, _14358_);
  or (_14364_, _14363_, _10926_);
  or (_14365_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_14366_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_14367_, _14366_, _10928_);
  and (_14368_, _14367_, _14365_);
  or (_14369_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_14370_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_14371_, _14370_, _04832_);
  and (_14372_, _14371_, _14369_);
  or (_14373_, _14372_, _14368_);
  or (_14374_, _14373_, _04868_);
  and (_14375_, _14374_, _04859_);
  and (_14376_, _14375_, _14364_);
  or (_14377_, _14376_, _14354_);
  or (_14378_, _14377_, _04849_);
  and (_14379_, _14378_, _10996_);
  and (_14380_, _14379_, _14332_);
  and (_14381_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_14382_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_14383_, _14382_, _14381_);
  and (_14384_, _14383_, _04832_);
  and (_14385_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_14386_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_14387_, _14386_, _14385_);
  and (_14388_, _14387_, _10928_);
  or (_14389_, _14388_, _14384_);
  and (_14390_, _14389_, _04868_);
  and (_14391_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_14392_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_14393_, _14392_, _14391_);
  and (_14394_, _14393_, _04832_);
  and (_14395_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_14396_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_14397_, _14396_, _14395_);
  and (_14398_, _14397_, _10928_);
  or (_14399_, _14398_, _14394_);
  and (_14400_, _14399_, _10926_);
  or (_14401_, _14400_, _04859_);
  or (_14402_, _14401_, _14390_);
  or (_14403_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_14404_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_14405_, _14404_, _10928_);
  and (_14406_, _14405_, _14403_);
  or (_14407_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_14408_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_14409_, _14408_, _04832_);
  and (_14410_, _14409_, _14407_);
  or (_14411_, _14410_, _14406_);
  and (_14412_, _14411_, _04868_);
  or (_14413_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_14414_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_14415_, _14414_, _10928_);
  and (_14416_, _14415_, _14413_);
  or (_14417_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_14418_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_14419_, _14418_, _04832_);
  and (_14420_, _14419_, _14417_);
  or (_14421_, _14420_, _14416_);
  and (_14422_, _14421_, _10926_);
  or (_14423_, _14422_, _10945_);
  or (_14424_, _14423_, _14412_);
  and (_14425_, _14424_, _14402_);
  or (_14426_, _14425_, _04849_);
  and (_14427_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and (_14428_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_14429_, _14428_, _14427_);
  and (_14430_, _14429_, _04832_);
  and (_14431_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_14432_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_14433_, _14432_, _14431_);
  and (_14434_, _14433_, _10928_);
  or (_14435_, _14434_, _14430_);
  and (_14436_, _14435_, _04868_);
  and (_14437_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and (_14438_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_14439_, _14438_, _14437_);
  and (_14440_, _14439_, _04832_);
  and (_14441_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and (_14442_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_14443_, _14442_, _14441_);
  and (_14444_, _14443_, _10928_);
  or (_14445_, _14444_, _14440_);
  and (_14446_, _14445_, _10926_);
  or (_14447_, _14446_, _04859_);
  or (_14448_, _14447_, _14436_);
  or (_14449_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_14450_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and (_14451_, _14450_, _14449_);
  and (_14452_, _14451_, _04832_);
  or (_14453_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_14454_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_14455_, _14454_, _14453_);
  and (_14456_, _14455_, _10928_);
  or (_14457_, _14456_, _14452_);
  and (_14458_, _14457_, _04868_);
  or (_14459_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_14460_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and (_14461_, _14460_, _14459_);
  and (_14462_, _14461_, _04832_);
  or (_14463_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_14464_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_14465_, _14464_, _14463_);
  and (_14466_, _14465_, _10928_);
  or (_14467_, _14466_, _14462_);
  and (_14468_, _14467_, _10926_);
  or (_14470_, _14468_, _10945_);
  or (_14471_, _14470_, _14458_);
  and (_14472_, _14471_, _14448_);
  or (_14473_, _14472_, _10997_);
  and (_14474_, _14473_, _04839_);
  and (_14475_, _14474_, _14426_);
  or (_14476_, _14475_, _14380_);
  or (_14477_, _14476_, _04843_);
  and (_14478_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  and (_14479_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or (_14480_, _14479_, _14478_);
  and (_14481_, _14480_, _04832_);
  and (_14482_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  and (_14483_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or (_14484_, _14483_, _14482_);
  and (_14485_, _14484_, _10928_);
  or (_14486_, _14485_, _14481_);
  and (_14487_, _14486_, _04868_);
  and (_14488_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  and (_14489_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or (_14490_, _14489_, _14488_);
  and (_14491_, _14490_, _04832_);
  and (_14492_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  and (_14493_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or (_14494_, _14493_, _14492_);
  and (_14495_, _14494_, _10928_);
  or (_14496_, _14495_, _14491_);
  and (_14497_, _14496_, _10926_);
  or (_14498_, _14497_, _04859_);
  or (_14499_, _14498_, _14487_);
  or (_14500_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or (_14501_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  and (_14502_, _14501_, _14500_);
  and (_14503_, _14502_, _04832_);
  or (_14504_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or (_14505_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  and (_14506_, _14505_, _14504_);
  and (_14507_, _14506_, _10928_);
  or (_14508_, _14507_, _14503_);
  and (_14509_, _14508_, _04868_);
  or (_14510_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or (_14511_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  and (_14512_, _14511_, _14510_);
  and (_14513_, _14512_, _04832_);
  or (_14514_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or (_14515_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  and (_14516_, _14515_, _14514_);
  and (_14517_, _14516_, _10928_);
  or (_14518_, _14517_, _14513_);
  and (_14519_, _14518_, _10926_);
  or (_14521_, _14519_, _10945_);
  or (_14522_, _14521_, _14509_);
  and (_14523_, _14522_, _14499_);
  or (_14524_, _14523_, _04849_);
  and (_14525_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_14526_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_14527_, _14526_, _14525_);
  and (_14528_, _14527_, _04832_);
  and (_14529_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and (_14530_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_14531_, _14530_, _14529_);
  and (_14532_, _14531_, _10928_);
  or (_14533_, _14532_, _14528_);
  and (_14534_, _14533_, _04868_);
  and (_14535_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_14536_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_14537_, _14536_, _14535_);
  and (_14538_, _14537_, _04832_);
  and (_14539_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_14540_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_14541_, _14540_, _14539_);
  and (_14542_, _14541_, _10928_);
  or (_14543_, _14542_, _14538_);
  and (_14544_, _14543_, _10926_);
  or (_14545_, _14544_, _04859_);
  or (_14546_, _14545_, _14534_);
  or (_14547_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_14548_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_14549_, _14548_, _14547_);
  and (_14550_, _14549_, _04832_);
  or (_14551_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_14552_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_14553_, _14552_, _14551_);
  and (_14554_, _14553_, _10928_);
  or (_14555_, _14554_, _14550_);
  and (_14556_, _14555_, _04868_);
  or (_14557_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_14558_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_14559_, _14558_, _14557_);
  and (_14560_, _14559_, _04832_);
  or (_14561_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_14562_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and (_14563_, _14562_, _14561_);
  and (_14564_, _14563_, _10928_);
  or (_14565_, _14564_, _14560_);
  and (_14566_, _14565_, _10926_);
  or (_14567_, _14566_, _10945_);
  or (_14568_, _14567_, _14556_);
  and (_14569_, _14568_, _14546_);
  or (_14570_, _14569_, _10997_);
  and (_14571_, _14570_, _04839_);
  and (_14572_, _14571_, _14524_);
  and (_14573_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_14574_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_14575_, _14574_, _14573_);
  and (_14576_, _14575_, _10928_);
  and (_14577_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and (_14578_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_14579_, _14578_, _14577_);
  and (_14580_, _14579_, _04832_);
  or (_14581_, _14580_, _14576_);
  or (_14582_, _14581_, _10926_);
  and (_14583_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and (_14584_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_14585_, _14584_, _14583_);
  and (_14586_, _14585_, _10928_);
  and (_14587_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_14588_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_14589_, _14588_, _14587_);
  and (_14590_, _14589_, _04832_);
  or (_14592_, _14590_, _14586_);
  or (_14593_, _14592_, _04868_);
  and (_14594_, _14593_, _10945_);
  and (_14595_, _14594_, _14582_);
  or (_14596_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_14597_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_14598_, _14597_, _04832_);
  and (_14599_, _14598_, _14596_);
  or (_14600_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_14601_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_14602_, _14601_, _10928_);
  and (_14603_, _14602_, _14600_);
  or (_14604_, _14603_, _14599_);
  or (_14605_, _14604_, _10926_);
  or (_14606_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_14607_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_14608_, _14607_, _04832_);
  and (_14609_, _14608_, _14606_);
  or (_14610_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_14611_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_14612_, _14611_, _10928_);
  and (_14613_, _14612_, _14610_);
  or (_14614_, _14613_, _14609_);
  or (_14615_, _14614_, _04868_);
  and (_14616_, _14615_, _04859_);
  and (_14617_, _14616_, _14605_);
  or (_14618_, _14617_, _14595_);
  and (_14619_, _14618_, _10997_);
  and (_14620_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_14621_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_14622_, _14621_, _04832_);
  or (_14623_, _14622_, _14620_);
  and (_14624_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_14625_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_14626_, _14625_, _10928_);
  or (_14627_, _14626_, _14624_);
  and (_14628_, _14627_, _14623_);
  or (_14629_, _14628_, _10926_);
  and (_14630_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_14631_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_14632_, _14631_, _04832_);
  or (_14633_, _14632_, _14630_);
  and (_14634_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_14635_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_14636_, _14635_, _10928_);
  or (_14637_, _14636_, _14634_);
  and (_14638_, _14637_, _14633_);
  or (_14639_, _14638_, _04868_);
  and (_14640_, _14639_, _10945_);
  and (_14641_, _14640_, _14629_);
  or (_14642_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_14643_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_14644_, _14643_, _14642_);
  or (_14645_, _14644_, _10928_);
  or (_14646_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_14647_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_14648_, _14647_, _14646_);
  or (_14649_, _14648_, _04832_);
  and (_14650_, _14649_, _14645_);
  or (_14651_, _14650_, _10926_);
  or (_14653_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_14654_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_14655_, _14654_, _14653_);
  or (_14656_, _14655_, _10928_);
  or (_14657_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_14658_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_14659_, _14658_, _14657_);
  or (_14660_, _14659_, _04832_);
  and (_14661_, _14660_, _14656_);
  or (_14662_, _14661_, _04868_);
  and (_14663_, _14662_, _04859_);
  and (_14664_, _14663_, _14651_);
  or (_14665_, _14664_, _14641_);
  and (_14666_, _14665_, _04849_);
  or (_14667_, _14666_, _14619_);
  and (_14668_, _14667_, _10996_);
  or (_14669_, _14668_, _14572_);
  or (_14670_, _14669_, _11204_);
  and (_14671_, _14670_, _14477_);
  or (_14672_, _14671_, _26153_);
  and (_14673_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_14674_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_14675_, _14674_, _14673_);
  and (_14676_, _14675_, _04832_);
  and (_14677_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_14678_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_14679_, _14678_, _14677_);
  and (_14680_, _14679_, _10928_);
  or (_14681_, _14680_, _14676_);
  or (_14682_, _14681_, _10926_);
  and (_14683_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_14684_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_14685_, _14684_, _14683_);
  and (_14686_, _14685_, _04832_);
  and (_14687_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_14688_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_14689_, _14688_, _14687_);
  and (_14690_, _14689_, _10928_);
  or (_14691_, _14690_, _14686_);
  or (_14692_, _14691_, _04868_);
  and (_14693_, _14692_, _10945_);
  and (_14694_, _14693_, _14682_);
  or (_14695_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_14696_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_14697_, _14696_, _14695_);
  and (_14698_, _14697_, _04832_);
  or (_14699_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_14700_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_14701_, _14700_, _14699_);
  and (_14702_, _14701_, _10928_);
  or (_14703_, _14702_, _14698_);
  or (_14704_, _14703_, _10926_);
  or (_14705_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_14706_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_14707_, _14706_, _14705_);
  and (_14708_, _14707_, _04832_);
  or (_14709_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_14710_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_14711_, _14710_, _14709_);
  and (_14712_, _14711_, _10928_);
  or (_14713_, _14712_, _14708_);
  or (_14714_, _14713_, _04868_);
  and (_14715_, _14714_, _04859_);
  and (_14716_, _14715_, _14704_);
  or (_14717_, _14716_, _14694_);
  and (_14718_, _14717_, _04849_);
  and (_14719_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_14720_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_14721_, _14720_, _14719_);
  and (_14722_, _14721_, _04832_);
  and (_14723_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_14724_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_14725_, _14724_, _14723_);
  and (_14726_, _14725_, _10928_);
  or (_14727_, _14726_, _14722_);
  or (_14728_, _14727_, _10926_);
  and (_14729_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_14730_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_14731_, _14730_, _14729_);
  and (_14732_, _14731_, _04832_);
  and (_14733_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_14734_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_14735_, _14734_, _14733_);
  and (_14736_, _14735_, _10928_);
  or (_14737_, _14736_, _14732_);
  or (_14738_, _14737_, _04868_);
  and (_14739_, _14738_, _10945_);
  and (_14740_, _14739_, _14728_);
  or (_14741_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_14742_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_14744_, _14742_, _10928_);
  and (_14745_, _14744_, _14741_);
  or (_14746_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_14747_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_14748_, _14747_, _04832_);
  and (_14749_, _14748_, _14746_);
  or (_14750_, _14749_, _14745_);
  or (_14751_, _14750_, _10926_);
  or (_14752_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_14753_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_14754_, _14753_, _10928_);
  and (_14755_, _14754_, _14752_);
  or (_14756_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_14757_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_14758_, _14757_, _04832_);
  and (_14759_, _14758_, _14756_);
  or (_14760_, _14759_, _14755_);
  or (_14761_, _14760_, _04868_);
  and (_14762_, _14761_, _04859_);
  and (_14763_, _14762_, _14751_);
  or (_14764_, _14763_, _14740_);
  and (_14765_, _14764_, _10997_);
  or (_14766_, _14765_, _14718_);
  and (_14767_, _14766_, _10996_);
  and (_14768_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_14769_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_14770_, _14769_, _14768_);
  and (_14771_, _14770_, _04832_);
  and (_14772_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_14773_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_14774_, _14773_, _14772_);
  and (_14775_, _14774_, _10928_);
  or (_14776_, _14775_, _14771_);
  and (_14777_, _14776_, _04868_);
  and (_14778_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_14779_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_14780_, _14779_, _14778_);
  and (_14781_, _14780_, _04832_);
  and (_14782_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_14783_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_14784_, _14783_, _14782_);
  and (_14785_, _14784_, _10928_);
  or (_14786_, _14785_, _14781_);
  and (_14787_, _14786_, _10926_);
  or (_14788_, _14787_, _14777_);
  and (_14789_, _14788_, _10945_);
  or (_14790_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_14791_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_14792_, _14791_, _10928_);
  and (_14793_, _14792_, _14790_);
  or (_14794_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_14795_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and (_14796_, _14795_, _04832_);
  and (_14797_, _14796_, _14794_);
  or (_14798_, _14797_, _14793_);
  and (_14799_, _14798_, _04868_);
  or (_14800_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_14801_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and (_14802_, _14801_, _10928_);
  and (_14803_, _14802_, _14800_);
  or (_14804_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_14805_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_14806_, _14805_, _04832_);
  and (_14807_, _14806_, _14804_);
  or (_14808_, _14807_, _14803_);
  and (_14809_, _14808_, _10926_);
  or (_14810_, _14809_, _14799_);
  and (_14811_, _14810_, _04859_);
  or (_14812_, _14811_, _14789_);
  and (_14813_, _14812_, _10997_);
  and (_14814_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_14815_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_14816_, _14815_, _14814_);
  and (_14817_, _14816_, _04832_);
  and (_14818_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_14819_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_14820_, _14819_, _14818_);
  and (_14821_, _14820_, _10928_);
  or (_14822_, _14821_, _14817_);
  and (_14823_, _14822_, _04868_);
  and (_14824_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_14825_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_14826_, _14825_, _14824_);
  and (_14827_, _14826_, _04832_);
  and (_14828_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_14829_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_14830_, _14829_, _14828_);
  and (_14831_, _14830_, _10928_);
  or (_14832_, _14831_, _14827_);
  and (_14833_, _14832_, _10926_);
  or (_14834_, _14833_, _14823_);
  and (_14835_, _14834_, _10945_);
  or (_14836_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_14837_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_14838_, _14837_, _14836_);
  and (_14839_, _14838_, _04832_);
  or (_14840_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_14841_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_14842_, _14841_, _14840_);
  and (_14843_, _14842_, _10928_);
  or (_14844_, _14843_, _14839_);
  and (_14845_, _14844_, _04868_);
  or (_14846_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_14847_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_14848_, _14847_, _14846_);
  and (_14849_, _14848_, _04832_);
  or (_14850_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_14851_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_14852_, _14851_, _14850_);
  and (_14853_, _14852_, _10928_);
  or (_14854_, _14853_, _14849_);
  and (_14855_, _14854_, _10926_);
  or (_14856_, _14855_, _14845_);
  and (_14857_, _14856_, _04859_);
  or (_14858_, _14857_, _14835_);
  and (_14859_, _14858_, _04849_);
  or (_14860_, _14859_, _14813_);
  and (_14861_, _14860_, _04839_);
  or (_14862_, _14861_, _14767_);
  or (_14863_, _14862_, _04843_);
  and (_14864_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_14865_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_14866_, _14865_, _14864_);
  and (_14867_, _14866_, _04832_);
  and (_14868_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_14869_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_14870_, _14869_, _14868_);
  and (_14871_, _14870_, _10928_);
  or (_14872_, _14871_, _14867_);
  or (_14873_, _14872_, _10926_);
  and (_14874_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_14875_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_14876_, _14875_, _14874_);
  and (_14877_, _14876_, _04832_);
  and (_14878_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_14879_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_14880_, _14879_, _14878_);
  and (_14881_, _14880_, _10928_);
  or (_14882_, _14881_, _14877_);
  or (_14883_, _14882_, _04868_);
  and (_14884_, _14883_, _10945_);
  and (_14885_, _14884_, _14873_);
  or (_14886_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_14887_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_14888_, _14887_, _10928_);
  and (_14889_, _14888_, _14886_);
  or (_14890_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_14891_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_14892_, _14891_, _04832_);
  and (_14893_, _14892_, _14890_);
  or (_14894_, _14893_, _14889_);
  or (_14895_, _14894_, _10926_);
  or (_14896_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_14897_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_14898_, _14897_, _10928_);
  and (_14899_, _14898_, _14896_);
  or (_14900_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_14901_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_14902_, _14901_, _04832_);
  and (_14903_, _14902_, _14900_);
  or (_14904_, _14903_, _14899_);
  or (_14905_, _14904_, _04868_);
  and (_14906_, _14905_, _04859_);
  and (_14907_, _14906_, _14895_);
  or (_14908_, _14907_, _14885_);
  and (_14909_, _14908_, _10997_);
  and (_14910_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_14911_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_14912_, _14911_, _14910_);
  and (_14913_, _14912_, _04832_);
  and (_14914_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_14915_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_14916_, _14915_, _14914_);
  and (_14917_, _14916_, _10928_);
  or (_14918_, _14917_, _14913_);
  or (_14919_, _14918_, _10926_);
  and (_14920_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_14921_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_14922_, _14921_, _14920_);
  and (_14923_, _14922_, _04832_);
  and (_14924_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_14925_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_14926_, _14925_, _14924_);
  and (_14927_, _14926_, _10928_);
  or (_14928_, _14927_, _14923_);
  or (_14929_, _14928_, _04868_);
  and (_14930_, _14929_, _10945_);
  and (_14931_, _14930_, _14919_);
  or (_14932_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_14933_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_14934_, _14933_, _14932_);
  and (_14935_, _14934_, _04832_);
  or (_14936_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_14937_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_14938_, _14937_, _14936_);
  and (_14939_, _14938_, _10928_);
  or (_14940_, _14939_, _14935_);
  or (_14941_, _14940_, _10926_);
  or (_14942_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_14943_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_14944_, _14943_, _14942_);
  and (_14945_, _14944_, _04832_);
  or (_14946_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_14947_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_14948_, _14947_, _14946_);
  and (_14949_, _14948_, _10928_);
  or (_14950_, _14949_, _14945_);
  or (_14951_, _14950_, _04868_);
  and (_14952_, _14951_, _04859_);
  and (_14953_, _14952_, _14941_);
  or (_14954_, _14953_, _14931_);
  and (_14955_, _14954_, _04849_);
  or (_14956_, _14955_, _14909_);
  and (_14957_, _14956_, _10996_);
  or (_14958_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_14959_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_14960_, _14959_, _14958_);
  and (_14961_, _14960_, _04832_);
  or (_14962_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_14963_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_14964_, _14963_, _14962_);
  and (_14965_, _14964_, _10928_);
  or (_14966_, _14965_, _14961_);
  and (_14967_, _14966_, _10926_);
  or (_14968_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_14969_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_14970_, _14969_, _14968_);
  and (_14971_, _14970_, _04832_);
  or (_14972_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_14973_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_14975_, _14973_, _14972_);
  and (_14976_, _14975_, _10928_);
  or (_14977_, _14976_, _14971_);
  and (_14978_, _14977_, _04868_);
  or (_14979_, _14978_, _14967_);
  and (_14980_, _14979_, _04859_);
  and (_14981_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_14982_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_14983_, _14982_, _14981_);
  and (_14984_, _14983_, _04832_);
  and (_14985_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_14986_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_14987_, _14986_, _14985_);
  and (_14988_, _14987_, _10928_);
  or (_14989_, _14988_, _14984_);
  and (_14990_, _14989_, _10926_);
  and (_14991_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_14992_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_14993_, _14992_, _14991_);
  and (_14994_, _14993_, _04832_);
  and (_14996_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_14997_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_14998_, _14997_, _14996_);
  and (_14999_, _14998_, _10928_);
  or (_15000_, _14999_, _14994_);
  and (_15001_, _15000_, _04868_);
  or (_15002_, _15001_, _14990_);
  and (_15003_, _15002_, _10945_);
  or (_15004_, _15003_, _14980_);
  and (_15005_, _15004_, _04849_);
  or (_15006_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_15007_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_15008_, _15007_, _10928_);
  and (_15009_, _15008_, _15006_);
  or (_15010_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_15011_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_15012_, _15011_, _04832_);
  and (_15013_, _15012_, _15010_);
  or (_15014_, _15013_, _15009_);
  and (_15015_, _15014_, _10926_);
  or (_15016_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_15017_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_15018_, _15017_, _10928_);
  and (_15019_, _15018_, _15016_);
  or (_15020_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_15021_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_15022_, _15021_, _04832_);
  and (_15023_, _15022_, _15020_);
  or (_15024_, _15023_, _15019_);
  and (_15025_, _15024_, _04868_);
  or (_15026_, _15025_, _15015_);
  and (_15027_, _15026_, _04859_);
  and (_15028_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_15029_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_15030_, _15029_, _15028_);
  and (_15031_, _15030_, _04832_);
  and (_15032_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_15033_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_15034_, _15033_, _15032_);
  and (_15035_, _15034_, _10928_);
  or (_15036_, _15035_, _15031_);
  and (_15037_, _15036_, _10926_);
  and (_15038_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_15039_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_15040_, _15039_, _15038_);
  and (_15041_, _15040_, _04832_);
  and (_15042_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_15043_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_15044_, _15043_, _15042_);
  and (_15045_, _15044_, _10928_);
  or (_15047_, _15045_, _15041_);
  and (_15048_, _15047_, _04868_);
  or (_15049_, _15048_, _15037_);
  and (_15050_, _15049_, _10945_);
  or (_15051_, _15050_, _15027_);
  and (_15052_, _15051_, _10997_);
  or (_15053_, _15052_, _15005_);
  and (_15054_, _15053_, _04839_);
  or (_15055_, _15054_, _14957_);
  or (_15056_, _15055_, _11204_);
  and (_15057_, _15056_, _14863_);
  or (_15058_, _15057_, _03196_);
  and (_15059_, _15058_, _14672_);
  or (_15060_, _15059_, _04876_);
  or (_15061_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_15062_, _15061_, _22773_);
  and (_27321_[6], _15062_, _15060_);
  and (_15063_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_15064_, _09597_, _24053_);
  or (_05928_, _15064_, _15063_);
  and (_15065_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  and (_15066_, _09603_, _23983_);
  or (_05931_, _15066_, _15065_);
  and (_15067_, _02663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  and (_15068_, _02662_, _23920_);
  or (_05940_, _15068_, _15067_);
  and (_15069_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  and (_15070_, _03157_, _23983_);
  or (_05942_, _15070_, _15069_);
  and (_15071_, _03158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  and (_15072_, _03157_, _24027_);
  or (_05945_, _15072_, _15071_);
  and (_15073_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  and (_15074_, _09965_, _23983_);
  or (_05954_, _15074_, _15073_);
  and (_15075_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_15076_, _09944_, _23900_);
  or (_05964_, _15076_, _15075_);
  and (_15077_, _25165_, _23983_);
  and (_15078_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_26937_, _15078_, _15077_);
  and (_15079_, _10669_, _23905_);
  not (_15080_, _15079_);
  and (_15081_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nor (_15082_, _15080_, _23982_);
  or (_26944_, _15082_, _15081_);
  and (_05970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _22773_);
  and (_15083_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and (_15084_, _12688_, _23750_);
  or (_05972_, _15084_, _15083_);
  and (_15085_, _09945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_15086_, _09944_, _24053_);
  or (_05975_, _15086_, _15085_);
  and (_15087_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_15088_, _09910_, _23920_);
  or (_05981_, _15088_, _15087_);
  and (_15089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _22773_);
  and (_05984_, _15089_, _24855_);
  and (_15090_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  and (_15091_, _12688_, _24052_);
  or (_05986_, _15091_, _15090_);
  and (_15093_, _09831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and (_15094_, _09830_, _24053_);
  or (_06002_, _15094_, _15093_);
  and (_15095_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_15096_, _09778_, _23751_);
  or (_06009_, _15096_, _15095_);
  and (_15097_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  and (_15098_, _02748_, _23920_);
  or (_06038_, _15098_, _15097_);
  and (_15099_, _01927_, _23751_);
  and (_15100_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_06040_, _15100_, _15099_);
  and (_15101_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and (_15102_, _09603_, _23751_);
  or (_26960_, _15102_, _15101_);
  and (_15103_, _01927_, _24053_);
  and (_15104_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_26957_, _15104_, _15103_);
  and (_15105_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_15107_, _09722_, _23693_);
  or (_26959_, _15107_, _15105_);
  and (_15108_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and (_15109_, _02748_, _23900_);
  or (_06046_, _15109_, _15108_);
  and (_15110_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and (_15111_, _12688_, _23692_);
  or (_06050_, _15111_, _15110_);
  and (_15112_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and (_15113_, _09647_, _23715_);
  or (_06056_, _15113_, _15112_);
  and (_15114_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and (_15115_, _12688_, _23899_);
  or (_06062_, _15115_, _15114_);
  and (_15116_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and (_15117_, _02748_, _23715_);
  or (_06064_, _15117_, _15116_);
  and (_15118_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and (_15119_, _09620_, _23900_);
  or (_06067_, _15119_, _15118_);
  and (_15121_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  and (_15122_, _12688_, _23714_);
  or (_06075_, _15122_, _15121_);
  and (_15123_, _25169_, _23900_);
  and (_15124_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_06078_, _15124_, _15123_);
  and (_15125_, _01927_, _23900_);
  and (_15126_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_06083_, _15126_, _15125_);
  and (_15127_, _25190_, _23900_);
  and (_15128_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_06089_, _15128_, _15127_);
  and (_15129_, _01927_, _23715_);
  and (_15130_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_06092_, _15130_, _15129_);
  and (_15131_, _09480_, _23715_);
  and (_15132_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or (_27041_, _15132_, _15131_);
  and (_15133_, _09912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_15134_, _09910_, _23751_);
  or (_06099_, _15134_, _15133_);
  and (_15136_, _09867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  and (_15137_, _09866_, _23693_);
  or (_06101_, _15137_, _15136_);
  and (_15138_, _09779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_15139_, _09778_, _23920_);
  or (_06110_, _15139_, _15138_);
  and (_15140_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  and (_15141_, _09603_, _23920_);
  or (_06114_, _15141_, _15140_);
  and (_15142_, _09723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_15143_, _09722_, _24027_);
  or (_06119_, _15143_, _15142_);
  and (_15144_, _09648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and (_15145_, _09647_, _23983_);
  or (_06125_, _15145_, _15144_);
  and (_15146_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_15147_, _15079_, _24052_);
  or (_06127_, _15147_, _15146_);
  and (_15148_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  and (_15149_, _02748_, _24027_);
  or (_06129_, _15149_, _15148_);
  and (_15150_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_15151_, _15079_, _23692_);
  or (_06153_, _15151_, _15150_);
  and (_15152_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_15153_, _09597_, _23900_);
  or (_26962_, _15153_, _15152_);
  and (_15154_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_15155_, _15079_, _23750_);
  or (_06161_, _15155_, _15154_);
  and (_15156_, _09967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and (_15157_, _09965_, _24053_);
  or (_26972_, _15157_, _15156_);
  and (_15158_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  and (_15159_, _02748_, _23983_);
  or (_06166_, _15159_, _15158_);
  or (_15160_, _24188_, _23205_);
  nand (_15161_, _10280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_15162_, _10285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_15163_, _15162_, _15161_);
  nor (_15164_, _15163_, _24192_);
  nand (_15165_, _24989_, _07311_);
  and (_15166_, _15165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_15167_, _15166_, _15164_);
  or (_15168_, _15167_, _24186_);
  and (_15169_, _15168_, _22773_);
  and (_06170_, _15169_, _15160_);
  and (_15170_, _09598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_15171_, _09597_, _24027_);
  or (_06176_, _15171_, _15170_);
  and (_15172_, _24053_, _23925_);
  and (_15173_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_06185_, _15173_, _15172_);
  and (_15174_, _25169_, _23983_);
  and (_15175_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_06193_, _15175_, _15174_);
  and (_15176_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  and (_15177_, _10431_, _24027_);
  or (_06211_, _15177_, _15176_);
  and (_15178_, _10564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_15179_, _10563_, _23751_);
  or (_06218_, _15179_, _15178_);
  and (_15180_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and (_15181_, _10799_, _23714_);
  or (_26946_, _15181_, _15180_);
  and (_15182_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nor (_15183_, _15080_, _24026_);
  or (_06248_, _15183_, _15182_);
  and (_15184_, _10669_, _23444_);
  not (_15185_, _15184_);
  and (_15186_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_15187_, _15184_, _23750_);
  or (_26942_, _15187_, _15186_);
  and (_15188_, _10669_, _24108_);
  not (_15189_, _15188_);
  and (_15190_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_15191_, _15188_, _23750_);
  or (_06267_, _15191_, _15190_);
  and (_15192_, _25440_, _23751_);
  and (_15193_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or (_06270_, _15193_, _15192_);
  or (_15194_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_15195_, _15194_, _24330_);
  and (_15196_, _25226_, _24405_);
  nand (_15197_, _15196_, _23681_);
  and (_15198_, _15197_, _15195_);
  nand (_15199_, _25236_, _24047_);
  and (_15200_, _15194_, _22915_);
  and (_15201_, _15200_, _15199_);
  nor (_15202_, _22914_, _03773_);
  or (_15203_, _15202_, rst);
  or (_15204_, _15203_, _15201_);
  or (_06272_, _15204_, _15198_);
  and (_15205_, _10669_, _24235_);
  not (_15206_, _15205_);
  and (_15207_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  nor (_15208_, _15206_, _24026_);
  or (_06277_, _15208_, _15207_);
  and (_15209_, _10669_, _23890_);
  not (_15210_, _15209_);
  and (_15211_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nor (_15212_, _15210_, _24026_);
  or (_06280_, _15212_, _15211_);
  and (_15213_, _25316_, _22895_);
  nand (_15214_, _15213_, _23681_);
  or (_15215_, _15213_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_15216_, _15215_, _24330_);
  and (_15217_, _15216_, _15214_);
  or (_15218_, _02521_, _23744_);
  or (_15219_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_15220_, _15219_, _22915_);
  and (_15221_, _15220_, _15218_);
  nor (_15222_, _22914_, _03749_);
  or (_15223_, _15222_, rst);
  or (_15224_, _15223_, _15221_);
  or (_06283_, _15224_, _15217_);
  and (_15225_, _23924_, _23706_);
  and (_15226_, _15225_, _23900_);
  not (_15227_, _15225_);
  and (_15228_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_06293_, _15228_, _15226_);
  and (_15229_, _24145_, _23706_);
  and (_15230_, _15229_, _24027_);
  not (_15231_, _15229_);
  and (_15232_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or (_26930_, _15232_, _15230_);
  and (_15233_, _07484_, _23715_);
  and (_15234_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_06311_, _15234_, _15233_);
  and (_26871_, _22773_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_15236_, _25482_, _23983_);
  and (_15237_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_27230_, _15237_, _15236_);
  and (_15238_, _24108_, _23706_);
  and (_15239_, _15238_, _24053_);
  not (_15240_, _15238_);
  and (_15241_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_06333_, _15241_, _15239_);
  and (_15242_, _04767_, _23751_);
  and (_15243_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_06340_, _15243_, _15242_);
  and (_15244_, _08435_, _23920_);
  and (_15245_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or (_06346_, _15245_, _15244_);
  and (_15246_, _24068_, _23706_);
  and (_15247_, _15246_, _23983_);
  not (_15248_, _15246_);
  and (_15249_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_06359_, _15249_, _15247_);
  and (_15251_, _12702_, _23983_);
  and (_15252_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or (_06366_, _15252_, _15251_);
  and (_15253_, _23707_, _23693_);
  and (_15254_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_06371_, _15254_, _15253_);
  and (_15255_, _23938_, _23706_);
  and (_15256_, _15255_, _23983_);
  not (_15257_, _15255_);
  and (_15258_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or (_06374_, _15258_, _15256_);
  and (_15259_, _08240_, _23693_);
  and (_15260_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_06375_, _15260_, _15259_);
  and (_15261_, _06631_, _23715_);
  and (_15262_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or (_26923_, _15262_, _15261_);
  and (_15263_, _06631_, _24053_);
  and (_15264_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or (_06382_, _15264_, _15263_);
  and (_15266_, _07484_, _23693_);
  and (_15267_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_27219_, _15267_, _15266_);
  and (_15268_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _01548_);
  and (_15269_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_15270_, _15269_, _15268_);
  and (_26870_[7], _15270_, _22773_);
  not (_15271_, _24490_);
  nand (_15272_, _24533_, _15271_);
  nor (_15273_, _15272_, _24661_);
  nor (_15274_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  nand (_15275_, _15274_, _23761_);
  nor (_15276_, _15275_, _24629_);
  and (_15277_, _24514_, _24556_);
  and (_15278_, _15277_, _15276_);
  not (_15279_, _24580_);
  and (_15280_, _24605_, _15279_);
  and (_15281_, _15280_, _15278_);
  and (_26869_, _15281_, _15273_);
  and (_15282_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_15284_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_15285_, _15284_, _15282_);
  and (_15286_, _15285_, _04832_);
  and (_15287_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_15288_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_15289_, _15288_, _15287_);
  and (_15290_, _15289_, _10928_);
  or (_15291_, _15290_, _15286_);
  or (_15292_, _15291_, _10926_);
  and (_15293_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_15294_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_15295_, _15294_, _15293_);
  and (_15296_, _15295_, _04832_);
  and (_15297_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_15298_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_15299_, _15298_, _15297_);
  and (_15300_, _15299_, _10928_);
  or (_15301_, _15300_, _15296_);
  or (_15302_, _15301_, _04868_);
  and (_15303_, _15302_, _10945_);
  and (_15304_, _15303_, _15292_);
  or (_15305_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_15306_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_15307_, _15306_, _15305_);
  and (_15308_, _15307_, _04832_);
  or (_15309_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_15310_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_15311_, _15310_, _15309_);
  and (_15312_, _15311_, _10928_);
  or (_15313_, _15312_, _15308_);
  or (_15314_, _15313_, _10926_);
  or (_15315_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_15316_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_15317_, _15316_, _15315_);
  and (_15318_, _15317_, _04832_);
  or (_15319_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_15320_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_15321_, _15320_, _15319_);
  and (_15322_, _15321_, _10928_);
  or (_15323_, _15322_, _15318_);
  or (_15325_, _15323_, _04868_);
  and (_15326_, _15325_, _04859_);
  and (_15327_, _15326_, _15314_);
  or (_15328_, _15327_, _15304_);
  and (_15329_, _15328_, _04849_);
  and (_15330_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_15331_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_15332_, _15331_, _15330_);
  and (_15333_, _15332_, _04832_);
  and (_15334_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_15335_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_15336_, _15335_, _15334_);
  and (_15337_, _15336_, _10928_);
  or (_15338_, _15337_, _15333_);
  or (_15339_, _15338_, _10926_);
  and (_15340_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_15341_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_15342_, _15341_, _15340_);
  and (_15343_, _15342_, _04832_);
  and (_15344_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_15345_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_15346_, _15345_, _15344_);
  and (_15347_, _15346_, _10928_);
  or (_15348_, _15347_, _15343_);
  or (_15349_, _15348_, _04868_);
  and (_15350_, _15349_, _10945_);
  and (_15351_, _15350_, _15339_);
  or (_15352_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_15353_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and (_15354_, _15353_, _10928_);
  and (_15355_, _15354_, _15352_);
  or (_15356_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_15357_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and (_15358_, _15357_, _04832_);
  and (_15359_, _15358_, _15356_);
  or (_15360_, _15359_, _15355_);
  or (_15361_, _15360_, _10926_);
  or (_15362_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_15363_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_15364_, _15363_, _10928_);
  and (_15365_, _15364_, _15362_);
  or (_15366_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_15367_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_15368_, _15367_, _04832_);
  and (_15369_, _15368_, _15366_);
  or (_15370_, _15369_, _15365_);
  or (_15371_, _15370_, _04868_);
  and (_15372_, _15371_, _04859_);
  and (_15373_, _15372_, _15361_);
  or (_15374_, _15373_, _15351_);
  and (_15375_, _15374_, _10997_);
  or (_15376_, _15375_, _15329_);
  and (_15377_, _15376_, _10996_);
  and (_15378_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_15379_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_15380_, _15379_, _15378_);
  and (_15381_, _15380_, _04832_);
  and (_15382_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_15383_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_15384_, _15383_, _15382_);
  and (_15385_, _15384_, _10928_);
  or (_15386_, _15385_, _15381_);
  and (_15387_, _15386_, _04868_);
  and (_15388_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_15389_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_15390_, _15389_, _15388_);
  and (_15391_, _15390_, _04832_);
  and (_15392_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_15393_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_15394_, _15393_, _15392_);
  and (_15395_, _15394_, _10928_);
  or (_15396_, _15395_, _15391_);
  and (_15397_, _15396_, _10926_);
  or (_15398_, _15397_, _15387_);
  and (_15399_, _15398_, _10945_);
  or (_15400_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_15401_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_15402_, _15401_, _10928_);
  and (_15403_, _15402_, _15400_);
  or (_15404_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_15405_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_15406_, _15405_, _04832_);
  and (_15407_, _15406_, _15404_);
  or (_15408_, _15407_, _15403_);
  and (_15409_, _15408_, _04868_);
  or (_15410_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_15411_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_15412_, _15411_, _10928_);
  and (_15413_, _15412_, _15410_);
  or (_15414_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_15415_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_15416_, _15415_, _04832_);
  and (_15417_, _15416_, _15414_);
  or (_15418_, _15417_, _15413_);
  and (_15419_, _15418_, _10926_);
  or (_15420_, _15419_, _15409_);
  and (_15421_, _15420_, _04859_);
  or (_15422_, _15421_, _15399_);
  and (_15423_, _15422_, _10997_);
  and (_15424_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_15425_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_15426_, _15425_, _15424_);
  and (_15427_, _15426_, _04832_);
  and (_15428_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and (_15429_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_15430_, _15429_, _15428_);
  and (_15431_, _15430_, _10928_);
  or (_15432_, _15431_, _15427_);
  and (_15433_, _15432_, _04868_);
  and (_15434_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_15435_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_15436_, _15435_, _15434_);
  and (_15437_, _15436_, _04832_);
  and (_15438_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_15439_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_15440_, _15439_, _15438_);
  and (_15441_, _15440_, _10928_);
  or (_15442_, _15441_, _15437_);
  and (_15443_, _15442_, _10926_);
  or (_15444_, _15443_, _15433_);
  and (_15445_, _15444_, _10945_);
  or (_15446_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_15447_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_15448_, _15447_, _15446_);
  and (_15449_, _15448_, _04832_);
  or (_15450_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_15451_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_15452_, _15451_, _15450_);
  and (_15453_, _15452_, _10928_);
  or (_15454_, _15453_, _15449_);
  and (_15455_, _15454_, _04868_);
  or (_15456_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_15457_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_15458_, _15457_, _15456_);
  and (_15459_, _15458_, _04832_);
  or (_15460_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_15461_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_15462_, _15461_, _15460_);
  and (_15463_, _15462_, _10928_);
  or (_15464_, _15463_, _15459_);
  and (_15466_, _15464_, _10926_);
  or (_15467_, _15466_, _15455_);
  and (_15468_, _15467_, _04859_);
  or (_15469_, _15468_, _15445_);
  and (_15470_, _15469_, _04849_);
  or (_15471_, _15470_, _15423_);
  and (_15472_, _15471_, _04839_);
  or (_15473_, _15472_, _15377_);
  or (_15474_, _15473_, _04843_);
  and (_15475_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_15476_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_15477_, _15476_, _15475_);
  and (_15478_, _15477_, _04832_);
  and (_15479_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_15480_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_15481_, _15480_, _15479_);
  and (_15482_, _15481_, _10928_);
  or (_15483_, _15482_, _15478_);
  or (_15484_, _15483_, _10926_);
  and (_15485_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_15487_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_15488_, _15487_, _15485_);
  and (_15489_, _15488_, _04832_);
  and (_15490_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_15491_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_15492_, _15491_, _15490_);
  and (_15493_, _15492_, _10928_);
  or (_15494_, _15493_, _15489_);
  or (_15495_, _15494_, _04868_);
  and (_15496_, _15495_, _10945_);
  and (_15497_, _15496_, _15484_);
  or (_15498_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_15499_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_15500_, _15499_, _10928_);
  and (_15501_, _15500_, _15498_);
  or (_15502_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_15503_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_15504_, _15503_, _04832_);
  and (_15505_, _15504_, _15502_);
  or (_15506_, _15505_, _15501_);
  or (_15508_, _15506_, _10926_);
  or (_15509_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_15510_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_15511_, _15510_, _10928_);
  and (_15512_, _15511_, _15509_);
  or (_15513_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_15514_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and (_15515_, _15514_, _04832_);
  and (_15516_, _15515_, _15513_);
  or (_15517_, _15516_, _15512_);
  or (_15518_, _15517_, _04868_);
  and (_15519_, _15518_, _04859_);
  and (_15520_, _15519_, _15508_);
  or (_15521_, _15520_, _15497_);
  and (_15522_, _15521_, _10997_);
  and (_15523_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_15524_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_15525_, _15524_, _15523_);
  and (_15526_, _15525_, _04832_);
  and (_15527_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_15528_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_15529_, _15528_, _15527_);
  and (_15530_, _15529_, _10928_);
  or (_15531_, _15530_, _15526_);
  or (_15532_, _15531_, _10926_);
  and (_15533_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_15534_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_15535_, _15534_, _15533_);
  and (_15536_, _15535_, _04832_);
  and (_15537_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_15538_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_15539_, _15538_, _15537_);
  and (_15540_, _15539_, _10928_);
  or (_15541_, _15540_, _15536_);
  or (_15542_, _15541_, _04868_);
  and (_15543_, _15542_, _10945_);
  and (_15544_, _15543_, _15532_);
  or (_15545_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_15546_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_15547_, _15546_, _15545_);
  and (_15548_, _15547_, _04832_);
  or (_15549_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_15550_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_15551_, _15550_, _15549_);
  and (_15552_, _15551_, _10928_);
  or (_15553_, _15552_, _15548_);
  or (_15554_, _15553_, _10926_);
  or (_15555_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_15556_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_15557_, _15556_, _15555_);
  and (_15558_, _15557_, _04832_);
  or (_15559_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_15560_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_15561_, _15560_, _15559_);
  and (_15562_, _15561_, _10928_);
  or (_15563_, _15562_, _15558_);
  or (_15564_, _15563_, _04868_);
  and (_15565_, _15564_, _04859_);
  and (_15566_, _15565_, _15554_);
  or (_15567_, _15566_, _15544_);
  and (_15568_, _15567_, _04849_);
  or (_15569_, _15568_, _15522_);
  and (_15570_, _15569_, _10996_);
  or (_15571_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_15572_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_15573_, _15572_, _15571_);
  and (_15574_, _15573_, _04832_);
  or (_15575_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_15576_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and (_15577_, _15576_, _15575_);
  and (_15578_, _15577_, _10928_);
  or (_15579_, _15578_, _15574_);
  and (_15580_, _15579_, _10926_);
  or (_15581_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_15582_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_15583_, _15582_, _15581_);
  and (_15584_, _15583_, _04832_);
  or (_15585_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_15586_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_15587_, _15586_, _15585_);
  and (_15588_, _15587_, _10928_);
  or (_15589_, _15588_, _15584_);
  and (_15590_, _15589_, _04868_);
  or (_15591_, _15590_, _15580_);
  and (_15592_, _15591_, _04859_);
  and (_15593_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_15594_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_15595_, _15594_, _15593_);
  and (_15596_, _15595_, _04832_);
  and (_15597_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_15598_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_15599_, _15598_, _15597_);
  and (_15600_, _15599_, _10928_);
  or (_15601_, _15600_, _15596_);
  and (_15602_, _15601_, _10926_);
  and (_15603_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_15604_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_15605_, _15604_, _15603_);
  and (_15606_, _15605_, _04832_);
  and (_15607_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_15608_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_15609_, _15608_, _15607_);
  and (_15610_, _15609_, _10928_);
  or (_15611_, _15610_, _15606_);
  and (_15612_, _15611_, _04868_);
  or (_15613_, _15612_, _15602_);
  and (_15614_, _15613_, _10945_);
  or (_15615_, _15614_, _15592_);
  and (_15616_, _15615_, _04849_);
  or (_15617_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_15618_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and (_15619_, _15618_, _10928_);
  and (_15620_, _15619_, _15617_);
  or (_15621_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_15622_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_15623_, _15622_, _04832_);
  and (_15624_, _15623_, _15621_);
  or (_15625_, _15624_, _15620_);
  and (_15626_, _15625_, _10926_);
  or (_15627_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_15628_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and (_15629_, _15628_, _10928_);
  and (_15630_, _15629_, _15627_);
  or (_15631_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_15632_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_15633_, _15632_, _04832_);
  and (_15634_, _15633_, _15631_);
  or (_15635_, _15634_, _15630_);
  and (_15636_, _15635_, _04868_);
  or (_15637_, _15636_, _15626_);
  and (_15638_, _15637_, _04859_);
  and (_15639_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_15640_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_15641_, _15640_, _15639_);
  and (_15642_, _15641_, _04832_);
  and (_15643_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and (_15644_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_15645_, _15644_, _15643_);
  and (_15646_, _15645_, _10928_);
  or (_15647_, _15646_, _15642_);
  and (_15648_, _15647_, _10926_);
  and (_15649_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and (_15650_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_15651_, _15650_, _15649_);
  and (_15652_, _15651_, _04832_);
  and (_15653_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_15654_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_15655_, _15654_, _15653_);
  and (_15656_, _15655_, _10928_);
  or (_15657_, _15656_, _15652_);
  and (_15658_, _15657_, _04868_);
  or (_15659_, _15658_, _15648_);
  and (_15660_, _15659_, _10945_);
  or (_15661_, _15660_, _15638_);
  and (_15662_, _15661_, _10997_);
  or (_15663_, _15662_, _15616_);
  and (_15664_, _15663_, _04839_);
  or (_15665_, _15664_, _15570_);
  or (_15666_, _15665_, _11204_);
  and (_15667_, _15666_, _15474_);
  or (_15668_, _15667_, _26153_);
  and (_15669_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_15670_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_15671_, _15670_, _15669_);
  and (_15672_, _15671_, _04832_);
  and (_15673_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_15674_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_15675_, _15674_, _15673_);
  and (_15676_, _15675_, _10928_);
  or (_15677_, _15676_, _15672_);
  or (_15678_, _15677_, _10926_);
  and (_15679_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_15680_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_15681_, _15680_, _15679_);
  and (_15682_, _15681_, _04832_);
  and (_15683_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_15684_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_15685_, _15684_, _15683_);
  and (_15686_, _15685_, _10928_);
  or (_15687_, _15686_, _15682_);
  or (_15688_, _15687_, _04868_);
  and (_15689_, _15688_, _10945_);
  and (_15690_, _15689_, _15678_);
  or (_15691_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_15692_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_15693_, _15692_, _15691_);
  and (_15694_, _15693_, _04832_);
  or (_15695_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_15696_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_15697_, _15696_, _15695_);
  and (_15698_, _15697_, _10928_);
  or (_15699_, _15698_, _15694_);
  or (_15700_, _15699_, _10926_);
  or (_15701_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_15702_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_15703_, _15702_, _15701_);
  and (_15704_, _15703_, _04832_);
  or (_15705_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_15706_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_15707_, _15706_, _15705_);
  and (_15708_, _15707_, _10928_);
  or (_15709_, _15708_, _15704_);
  or (_15710_, _15709_, _04868_);
  and (_15711_, _15710_, _04859_);
  and (_15712_, _15711_, _15700_);
  or (_15713_, _15712_, _15690_);
  and (_15714_, _15713_, _04849_);
  and (_15715_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_15716_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_15717_, _15716_, _15715_);
  and (_15718_, _15717_, _04832_);
  and (_15719_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_15720_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_15721_, _15720_, _15719_);
  and (_15722_, _15721_, _10928_);
  or (_15723_, _15722_, _15718_);
  or (_15724_, _15723_, _10926_);
  and (_15725_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_15726_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_15727_, _15726_, _15725_);
  and (_15728_, _15727_, _04832_);
  and (_15729_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_15730_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_15731_, _15730_, _15729_);
  and (_15732_, _15731_, _10928_);
  or (_15733_, _15732_, _15728_);
  or (_15734_, _15733_, _04868_);
  and (_15735_, _15734_, _10945_);
  and (_15736_, _15735_, _15724_);
  or (_15737_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_15738_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_15739_, _15738_, _10928_);
  and (_15740_, _15739_, _15737_);
  or (_15741_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_15742_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_15743_, _15742_, _04832_);
  and (_15744_, _15743_, _15741_);
  or (_15745_, _15744_, _15740_);
  or (_15746_, _15745_, _10926_);
  or (_15747_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_15749_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_15750_, _15749_, _10928_);
  and (_15751_, _15750_, _15747_);
  or (_15752_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_15753_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_15754_, _15753_, _04832_);
  and (_15755_, _15754_, _15752_);
  or (_15756_, _15755_, _15751_);
  or (_15757_, _15756_, _04868_);
  and (_15758_, _15757_, _04859_);
  and (_15759_, _15758_, _15746_);
  or (_15760_, _15759_, _15736_);
  and (_15761_, _15760_, _10997_);
  or (_15762_, _15761_, _15714_);
  and (_15763_, _15762_, _10996_);
  and (_15764_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_15765_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_15766_, _15765_, _15764_);
  and (_15767_, _15766_, _04832_);
  and (_15768_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_15770_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_15771_, _15770_, _15768_);
  and (_15772_, _15771_, _10928_);
  or (_15773_, _15772_, _15767_);
  and (_15774_, _15773_, _04868_);
  and (_15775_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and (_15776_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_15777_, _15776_, _15775_);
  and (_15778_, _15777_, _04832_);
  and (_15779_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_15780_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_15781_, _15780_, _15779_);
  and (_15782_, _15781_, _10928_);
  or (_15783_, _15782_, _15778_);
  and (_15784_, _15783_, _10926_);
  or (_15785_, _15784_, _15774_);
  and (_15786_, _15785_, _10945_);
  or (_15787_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_15788_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and (_15789_, _15788_, _10928_);
  and (_15791_, _15789_, _15787_);
  or (_15792_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_15793_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and (_15794_, _15793_, _04832_);
  and (_15795_, _15794_, _15792_);
  or (_15796_, _15795_, _15791_);
  and (_15797_, _15796_, _04868_);
  or (_15798_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_15799_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and (_15800_, _15799_, _10928_);
  and (_15801_, _15800_, _15798_);
  or (_15802_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_15803_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_15804_, _15803_, _04832_);
  and (_15805_, _15804_, _15802_);
  or (_15806_, _15805_, _15801_);
  and (_15807_, _15806_, _10926_);
  or (_15808_, _15807_, _15797_);
  and (_15809_, _15808_, _04859_);
  or (_15810_, _15809_, _15786_);
  and (_15811_, _15810_, _10997_);
  and (_15812_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_15813_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_15814_, _15813_, _15812_);
  and (_15815_, _15814_, _04832_);
  and (_15816_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_15817_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_15818_, _15817_, _15816_);
  and (_15819_, _15818_, _10928_);
  or (_15820_, _15819_, _15815_);
  and (_15821_, _15820_, _04868_);
  and (_15822_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_15823_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_15824_, _15823_, _15822_);
  and (_15825_, _15824_, _04832_);
  and (_15826_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_15827_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_15828_, _15827_, _15826_);
  and (_15829_, _15828_, _10928_);
  or (_15830_, _15829_, _15825_);
  and (_15831_, _15830_, _10926_);
  or (_15832_, _15831_, _15821_);
  and (_15833_, _15832_, _10945_);
  or (_15834_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_15835_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_15836_, _15835_, _15834_);
  and (_15837_, _15836_, _04832_);
  or (_15838_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_15839_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_15840_, _15839_, _15838_);
  and (_15841_, _15840_, _10928_);
  or (_15842_, _15841_, _15837_);
  and (_15843_, _15842_, _04868_);
  or (_15844_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_15845_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_15846_, _15845_, _15844_);
  and (_15847_, _15846_, _04832_);
  or (_15848_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_15849_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_15850_, _15849_, _15848_);
  and (_15851_, _15850_, _10928_);
  or (_15852_, _15851_, _15847_);
  and (_15853_, _15852_, _10926_);
  or (_15854_, _15853_, _15843_);
  and (_15855_, _15854_, _04859_);
  or (_15856_, _15855_, _15833_);
  and (_15857_, _15856_, _04849_);
  or (_15858_, _15857_, _15811_);
  and (_15859_, _15858_, _04839_);
  or (_15860_, _15859_, _15763_);
  or (_15861_, _15860_, _04843_);
  and (_15862_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_15863_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_15864_, _15863_, _15862_);
  and (_15865_, _15864_, _04832_);
  and (_15866_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_15867_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_15868_, _15867_, _15866_);
  and (_15869_, _15868_, _10928_);
  or (_15870_, _15869_, _15865_);
  or (_15871_, _15870_, _10926_);
  and (_15872_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_15873_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_15874_, _15873_, _15872_);
  and (_15875_, _15874_, _04832_);
  and (_15876_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_15877_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_15878_, _15877_, _15876_);
  and (_15879_, _15878_, _10928_);
  or (_15880_, _15879_, _15875_);
  or (_15882_, _15880_, _04868_);
  and (_15883_, _15882_, _10945_);
  and (_15884_, _15883_, _15871_);
  or (_15885_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_15886_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_15887_, _15886_, _10928_);
  and (_15888_, _15887_, _15885_);
  or (_15889_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_15890_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_15891_, _15890_, _04832_);
  and (_15892_, _15891_, _15889_);
  or (_15893_, _15892_, _15888_);
  or (_15894_, _15893_, _10926_);
  or (_15895_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_15896_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_15897_, _15896_, _10928_);
  and (_15898_, _15897_, _15895_);
  or (_15899_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_15900_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_15901_, _15900_, _04832_);
  and (_15902_, _15901_, _15899_);
  or (_15903_, _15902_, _15898_);
  or (_15904_, _15903_, _04868_);
  and (_15905_, _15904_, _04859_);
  and (_15906_, _15905_, _15894_);
  or (_15907_, _15906_, _15884_);
  and (_15908_, _15907_, _10997_);
  and (_15909_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_15910_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_15911_, _15910_, _15909_);
  and (_15912_, _15911_, _04832_);
  and (_15913_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_15914_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_15915_, _15914_, _15913_);
  and (_15916_, _15915_, _10928_);
  or (_15917_, _15916_, _15912_);
  or (_15918_, _15917_, _10926_);
  and (_15919_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_15920_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_15921_, _15920_, _15919_);
  and (_15922_, _15921_, _04832_);
  and (_15923_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_15924_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_15925_, _15924_, _15923_);
  and (_15926_, _15925_, _10928_);
  or (_15927_, _15926_, _15922_);
  or (_15928_, _15927_, _04868_);
  and (_15929_, _15928_, _10945_);
  and (_15930_, _15929_, _15918_);
  or (_15931_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_15932_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_15933_, _15932_, _15931_);
  and (_15934_, _15933_, _04832_);
  or (_15935_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_15936_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_15937_, _15936_, _15935_);
  and (_15938_, _15937_, _10928_);
  or (_15939_, _15938_, _15934_);
  or (_15940_, _15939_, _10926_);
  or (_15941_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_15942_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_15943_, _15942_, _15941_);
  and (_15944_, _15943_, _04832_);
  or (_15945_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_15946_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_15947_, _15946_, _15945_);
  and (_15948_, _15947_, _10928_);
  or (_15949_, _15948_, _15944_);
  or (_15950_, _15949_, _04868_);
  and (_15951_, _15950_, _04859_);
  and (_15953_, _15951_, _15940_);
  or (_15954_, _15953_, _15930_);
  and (_15955_, _15954_, _04849_);
  or (_15956_, _15955_, _15908_);
  and (_15957_, _15956_, _10996_);
  or (_15958_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_15959_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_15960_, _15959_, _15958_);
  and (_15961_, _15960_, _04832_);
  or (_15962_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_15963_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_15964_, _15963_, _15962_);
  and (_15965_, _15964_, _10928_);
  or (_15966_, _15965_, _15961_);
  and (_15967_, _15966_, _10926_);
  or (_15968_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_15969_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_15970_, _15969_, _15968_);
  and (_15971_, _15970_, _04832_);
  or (_15972_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_15973_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_15974_, _15973_, _15972_);
  and (_15975_, _15974_, _10928_);
  or (_15976_, _15975_, _15971_);
  and (_15977_, _15976_, _04868_);
  or (_15978_, _15977_, _15967_);
  and (_15979_, _15978_, _04859_);
  and (_15980_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_15981_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_15982_, _15981_, _15980_);
  and (_15983_, _15982_, _04832_);
  and (_15984_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_15985_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_15986_, _15985_, _15984_);
  and (_15987_, _15986_, _10928_);
  or (_15988_, _15987_, _15983_);
  and (_15989_, _15988_, _10926_);
  and (_15990_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_15991_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_15992_, _15991_, _15990_);
  and (_15993_, _15992_, _04832_);
  and (_15994_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_15995_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_15996_, _15995_, _15994_);
  and (_15997_, _15996_, _10928_);
  or (_15998_, _15997_, _15993_);
  and (_15999_, _15998_, _04868_);
  or (_16000_, _15999_, _15989_);
  and (_16001_, _16000_, _10945_);
  or (_16002_, _16001_, _15979_);
  and (_16004_, _16002_, _04849_);
  or (_16005_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_16006_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_16007_, _16006_, _10928_);
  and (_16008_, _16007_, _16005_);
  or (_16009_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_16010_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_16011_, _16010_, _04832_);
  and (_16012_, _16011_, _16009_);
  or (_16013_, _16012_, _16008_);
  and (_16014_, _16013_, _10926_);
  or (_16015_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_16016_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_16017_, _16016_, _10928_);
  and (_16018_, _16017_, _16015_);
  or (_16019_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_16020_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_16021_, _16020_, _04832_);
  and (_16022_, _16021_, _16019_);
  or (_16023_, _16022_, _16018_);
  and (_16024_, _16023_, _04868_);
  or (_16025_, _16024_, _16014_);
  and (_16026_, _16025_, _04859_);
  and (_16027_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_16028_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_16029_, _16028_, _16027_);
  and (_16030_, _16029_, _04832_);
  and (_16031_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_16032_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_16033_, _16032_, _16031_);
  and (_16034_, _16033_, _10928_);
  or (_16035_, _16034_, _16030_);
  and (_16036_, _16035_, _10926_);
  and (_16037_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_16038_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_16039_, _16038_, _16037_);
  and (_16040_, _16039_, _04832_);
  and (_16041_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_16042_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_16043_, _16042_, _16041_);
  and (_16044_, _16043_, _10928_);
  or (_16045_, _16044_, _16040_);
  and (_16046_, _16045_, _04868_);
  or (_16047_, _16046_, _16036_);
  and (_16048_, _16047_, _10945_);
  or (_16049_, _16048_, _16026_);
  and (_16050_, _16049_, _10997_);
  or (_16051_, _16050_, _16004_);
  and (_16052_, _16051_, _04839_);
  or (_16053_, _16052_, _15957_);
  or (_16054_, _16053_, _11204_);
  and (_16055_, _16054_, _15861_);
  or (_16056_, _16055_, _03196_);
  and (_16057_, _16056_, _15668_);
  or (_16058_, _16057_, _04876_);
  or (_16059_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_16060_, _16059_, _22773_);
  and (_06407_, _16060_, _16058_);
  and (_16061_, _10669_, _24061_);
  not (_16062_, _16061_);
  and (_16063_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  and (_16064_, _16061_, _23919_);
  or (_06433_, _16064_, _16063_);
  and (_16065_, _10669_, _24123_);
  not (_16066_, _16065_);
  and (_16067_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_16068_, _16065_, _23919_);
  or (_06436_, _16068_, _16067_);
  and (_16069_, _24975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_16070_, _25008_, _24984_);
  nor (_16071_, _16070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_16072_, _16071_, _02626_);
  and (_16073_, _10280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_16074_, _16073_, _16072_);
  and (_16075_, _16074_, _24976_);
  nor (_16076_, _16075_, _16069_);
  nor (_16077_, _16076_, _24192_);
  and (_16078_, _24192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_16079_, _16078_, _16077_);
  and (_16080_, _16079_, _24188_);
  nor (_16081_, _24188_, _24017_);
  or (_16082_, _16081_, _16080_);
  and (_06441_, _16082_, _22773_);
  or (_16083_, _23253_, _23205_);
  nor (_16084_, _10187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_16085_, _16084_, _10218_);
  and (_16086_, _16085_, _10189_);
  and (_16087_, _10191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_16088_, _24294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_16089_, _16088_, _23210_);
  or (_16090_, _16089_, _16087_);
  or (_16091_, _16090_, _16086_);
  or (_16092_, _16091_, _23252_);
  and (_16093_, _16092_, _22773_);
  and (_06454_, _16093_, _16083_);
  and (_16094_, _24274_, _23706_);
  and (_16095_, _16094_, _23900_);
  not (_16096_, _16094_);
  and (_16097_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or (_06460_, _16097_, _16095_);
  and (_16098_, _12702_, _23900_);
  and (_16099_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or (_06465_, _16099_, _16098_);
  and (_16100_, _24740_, _23920_);
  and (_16101_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_06477_, _16101_, _16100_);
  and (_16102_, _01745_, _23715_);
  and (_16103_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or (_06480_, _16103_, _16102_);
  and (_16104_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_16105_, _15079_, _23919_);
  or (_06481_, _16105_, _16104_);
  and (_16106_, _07484_, _23751_);
  and (_16107_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_06483_, _16107_, _16106_);
  and (_16108_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_16109_, _15079_, _23899_);
  or (_06520_, _16109_, _16108_);
  and (_16110_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  and (_16111_, _10799_, _23899_);
  or (_06523_, _16111_, _16110_);
  and (_16113_, _15080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_16114_, _15079_, _23714_);
  or (_06526_, _16114_, _16113_);
  and (_16115_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and (_16116_, _15184_, _23692_);
  or (_06528_, _16116_, _16115_);
  and (_16117_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and (_16118_, _15188_, _23692_);
  or (_06535_, _16118_, _16117_);
  and (_16119_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nor (_16120_, _15210_, _23982_);
  or (_06537_, _16120_, _16119_);
  and (_16121_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_16122_, _03161_, _24027_);
  or (_06538_, _16122_, _16121_);
  and (_16123_, _15229_, _23983_);
  and (_16124_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or (_26931_, _16124_, _16123_);
  and (_16125_, _04767_, _24027_);
  and (_16126_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_06546_, _16126_, _16125_);
  and (_16127_, _15246_, _23693_);
  and (_16128_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_26912_, _16128_, _16127_);
  and (_16129_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_16130_, _03161_, _23920_);
  or (_06550_, _16130_, _16129_);
  and (_16131_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_16132_, _03161_, _23900_);
  or (_06556_, _16132_, _16131_);
  and (_16133_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_16134_, _15184_, _23899_);
  or (_06559_, _16134_, _16133_);
  and (_16135_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_16136_, _15184_, _23714_);
  or (_06565_, _16136_, _16135_);
  and (_16137_, _08240_, _23983_);
  and (_16138_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_06601_, _16138_, _16137_);
  and (_16139_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  and (_16140_, _02748_, _23751_);
  or (_06604_, _16140_, _16139_);
  and (_16141_, _08240_, _23920_);
  and (_16142_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_06620_, _16142_, _16141_);
  and (_16143_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  nor (_16144_, _15185_, _23982_);
  or (_06622_, _16144_, _16143_);
  and (_16145_, _12702_, _24027_);
  and (_16146_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or (_06624_, _16146_, _16145_);
  and (_16147_, _02749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  and (_16148_, _02748_, _24053_);
  or (_27158_, _16148_, _16147_);
  and (_16149_, _06631_, _23751_);
  and (_16150_, _06633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or (_06634_, _16150_, _16149_);
  and (_16151_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  nor (_16152_, _15185_, _24026_);
  or (_06638_, _16152_, _16151_);
  and (_16153_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_16154_, _15184_, _23919_);
  or (_06640_, _16154_, _16153_);
  and (_16155_, _26273_, _25315_);
  nand (_16156_, _16155_, _24405_);
  or (_16157_, _16156_, _00619_);
  nand (_16158_, _16156_, _03513_);
  and (_16159_, _16158_, _22915_);
  and (_16160_, _16159_, _16157_);
  nor (_16161_, _22914_, _03513_);
  and (_16162_, _16155_, _24341_);
  nand (_16163_, _16162_, _23681_);
  or (_16164_, _16162_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_16165_, _16164_, _24330_);
  and (_16166_, _16165_, _16163_);
  or (_16167_, _16166_, _16161_);
  or (_16168_, _16167_, _16160_);
  and (_06644_, _16168_, _22773_);
  and (_16169_, _25190_, _23983_);
  and (_16170_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_06647_, _16170_, _16169_);
  and (_16171_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_16172_, _03161_, _23983_);
  or (_06650_, _16172_, _16171_);
  and (_16173_, _15255_, _24027_);
  and (_16174_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or (_06652_, _16174_, _16173_);
  and (_16175_, _08240_, _23900_);
  and (_16176_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_06660_, _16176_, _16175_);
  and (_16177_, _24027_, _23707_);
  and (_16178_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_06662_, _16178_, _16177_);
  and (_16179_, _23900_, _23707_);
  and (_16180_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_26910_, _16180_, _16179_);
  and (_16181_, _15246_, _23751_);
  and (_16182_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_06665_, _16182_, _16181_);
  and (_16183_, _25190_, _24027_);
  and (_16184_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_06668_, _16184_, _16183_);
  and (_16185_, _15246_, _23900_);
  and (_16186_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_06671_, _16186_, _16185_);
  and (_16187_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_16188_, _06621_, _23920_);
  or (_06673_, _16188_, _16187_);
  and (_16189_, _10669_, _23930_);
  not (_16190_, _16189_);
  and (_16191_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  nor (_16192_, _16190_, _24026_);
  or (_06677_, _16192_, _16191_);
  and (_16193_, _01745_, _23693_);
  and (_16194_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or (_06680_, _16194_, _16193_);
  and (_16195_, _01745_, _24053_);
  and (_16196_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or (_06682_, _16196_, _16195_);
  and (_16197_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  and (_16198_, _16189_, _23919_);
  or (_06683_, _16198_, _16197_);
  and (_16199_, _08435_, _24053_);
  and (_16200_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or (_06685_, _16200_, _16199_);
  and (_16201_, _01745_, _24027_);
  and (_16202_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or (_06687_, _16202_, _16201_);
  and (_16203_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and (_16204_, _16189_, _23899_);
  or (_06693_, _16204_, _16203_);
  and (_16205_, _08435_, _23715_);
  and (_16206_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or (_06695_, _16206_, _16205_);
  and (_16207_, _24740_, _24053_);
  and (_16208_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_06697_, _16208_, _16207_);
  and (_16209_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_16210_, _06621_, _24027_);
  or (_27155_, _16210_, _16209_);
  and (_16211_, _24740_, _23900_);
  and (_16212_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_06701_, _16212_, _16211_);
  and (_16213_, _04767_, _23920_);
  and (_16214_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_06708_, _16214_, _16213_);
  and (_16215_, _04767_, _23715_);
  and (_16216_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_06729_, _16216_, _16215_);
  and (_16217_, _15185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_16218_, _15184_, _24052_);
  or (_06731_, _16218_, _16217_);
  and (_16219_, _24157_, _23706_);
  and (_16220_, _16219_, _23751_);
  not (_16221_, _16219_);
  and (_16222_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or (_06734_, _16222_, _16220_);
  and (_16223_, _16219_, _23920_);
  and (_16224_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or (_06742_, _16224_, _16223_);
  and (_16225_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  nor (_16226_, _16190_, _23982_);
  or (_06744_, _16226_, _16225_);
  and (_16227_, _15238_, _24027_);
  and (_16228_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_06746_, _16228_, _16227_);
  and (_16229_, _12702_, _23715_);
  and (_16230_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or (_06749_, _16230_, _16229_);
  and (_16231_, _23905_, _23706_);
  and (_16232_, _16231_, _23920_);
  not (_16233_, _16231_);
  and (_16234_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_26927_, _16234_, _16232_);
  and (_16235_, _16231_, _23693_);
  and (_16236_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_26926_, _16236_, _16235_);
  and (_16237_, _16094_, _24053_);
  and (_16238_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or (_06757_, _16238_, _16237_);
  and (_16239_, _15229_, _24053_);
  and (_16240_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or (_06759_, _16240_, _16239_);
  and (_16241_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_16242_, _06621_, _23983_);
  or (_06761_, _16242_, _16241_);
  and (_16243_, _15229_, _23715_);
  and (_16244_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or (_06763_, _16244_, _16243_);
  and (_16245_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_16246_, _03161_, _23751_);
  or (_06766_, _16246_, _16245_);
  nand (_16247_, _24186_, _23357_);
  nand (_16248_, _16070_, _24976_);
  or (_16249_, _16248_, _24192_);
  and (_16250_, _16249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand (_16251_, _10280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_16252_, _16070_, _24975_);
  nand (_16253_, _16252_, _24989_);
  and (_16254_, _16253_, _16251_);
  nor (_16255_, _16254_, _24192_);
  or (_16256_, _16255_, _24186_);
  or (_16257_, _16256_, _16250_);
  and (_16258_, _16257_, _22773_);
  and (_06770_, _16258_, _16247_);
  and (_16259_, _24740_, _23715_);
  and (_16260_, _24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_26916_, _16260_, _16259_);
  and (_16261_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_16262_, _03161_, _24053_);
  or (_06774_, _16262_, _16261_);
  and (_16263_, _10669_, _23938_);
  not (_16264_, _16263_);
  and (_16265_, _16264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and (_16266_, _23938_, _23423_);
  and (_16267_, _23986_, _22856_);
  and (_16268_, _16267_, _16266_);
  and (_16269_, _16268_, _23919_);
  or (_26933_, _16269_, _16265_);
  and (_16270_, _10669_, _23700_);
  not (_16271_, _16270_);
  and (_16272_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_16273_, _16270_, _23714_);
  or (_06780_, _16273_, _16272_);
  and (_16274_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_16275_, _16270_, _24052_);
  or (_06781_, _16275_, _16274_);
  and (_16276_, _10669_, _24068_);
  not (_16277_, _16276_);
  and (_16278_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_16279_, _16276_, _23750_);
  or (_06784_, _16279_, _16278_);
  and (_16280_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  nor (_16281_, _16062_, _23982_);
  or (_06787_, _16281_, _16280_);
  and (_16282_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_16283_, _16276_, _23899_);
  or (_06790_, _16283_, _16282_);
  and (_16284_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nor (_16285_, _16062_, _24026_);
  or (_06793_, _16285_, _16284_);
  and (_16286_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and (_16287_, _15205_, _23692_);
  or (_06796_, _16287_, _16286_);
  and (_16288_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_16289_, _16065_, _23899_);
  or (_26939_, _16289_, _16288_);
  and (_16290_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_16291_, _16065_, _23750_);
  or (_26938_, _16291_, _16290_);
  and (_16292_, _10669_, _24157_);
  not (_16293_, _16292_);
  and (_16294_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and (_16295_, _16292_, _23899_);
  or (_06806_, _16295_, _16294_);
  and (_16296_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  nor (_16297_, _16293_, _23982_);
  or (_06826_, _16297_, _16296_);
  and (_16298_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  nor (_16299_, _15189_, _23982_);
  or (_06829_, _16299_, _16298_);
  and (_16300_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and (_16301_, _16061_, _23899_);
  or (_06835_, _16301_, _16300_);
  and (_16302_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and (_16303_, _16189_, _23692_);
  or (_06837_, _16303_, _16302_);
  and (_16304_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  and (_16305_, _16061_, _23692_);
  or (_06839_, _16305_, _16304_);
  and (_16306_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and (_16307_, _16189_, _23714_);
  or (_06841_, _16307_, _16306_);
  and (_16308_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  and (_16309_, _16189_, _24052_);
  or (_06843_, _16309_, _16308_);
  and (_16310_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  and (_16311_, _02756_, _23983_);
  or (_27152_, _16311_, _16310_);
  and (_16312_, _16190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and (_16313_, _16189_, _23750_);
  or (_26941_, _16313_, _16312_);
  and (_16314_, _12689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and (_16315_, _12688_, _23919_);
  or (_06848_, _16315_, _16314_);
  and (_16316_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  and (_16317_, _02756_, _24027_);
  or (_06852_, _16317_, _16316_);
  and (_16318_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  and (_16319_, _02756_, _23920_);
  or (_06854_, _16319_, _16318_);
  and (_16320_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and (_16321_, _10670_, _23692_);
  or (_06857_, _16321_, _16320_);
  and (_16322_, _10801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  nor (_16323_, _10801_, _23982_);
  or (_06859_, _16323_, _16322_);
  and (_16324_, _10671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor (_16325_, _10671_, _24026_);
  or (_06866_, _16325_, _16324_);
  and (_16326_, _02509_, _23900_);
  and (_16327_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_06875_, _16327_, _16326_);
  and (_16328_, _10432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  and (_16329_, _10431_, _23715_);
  or (_06877_, _16329_, _16328_);
  and (_16330_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  and (_16331_, _10303_, _23715_);
  or (_06879_, _16331_, _16330_);
  and (_16332_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  and (_16333_, _10303_, _24053_);
  or (_26951_, _16333_, _16332_);
  and (_16334_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_16335_, _10090_, _23751_);
  or (_26952_, _16335_, _16334_);
  and (_16336_, _10304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  and (_16337_, _10303_, _23983_);
  or (_06884_, _16337_, _16336_);
  and (_16338_, _10092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_16339_, _10090_, _23983_);
  or (_06888_, _16339_, _16338_);
  and (_16340_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  and (_16341_, _16061_, _23750_);
  or (_06890_, _16341_, _16340_);
  and (_16342_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  and (_16343_, _16061_, _24052_);
  or (_06893_, _16343_, _16342_);
  and (_16344_, _08240_, _23715_);
  and (_16345_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_06895_, _16345_, _16344_);
  and (_16346_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_16347_, _06621_, _23751_);
  or (_06898_, _16347_, _16346_);
  and (_16348_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_16349_, _09579_, _23900_);
  or (_06899_, _16349_, _16348_);
  and (_16350_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_16351_, _09579_, _23751_);
  or (_06902_, _16351_, _16350_);
  and (_16352_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_16353_, _06621_, _23715_);
  or (_27154_, _16353_, _16352_);
  and (_16354_, _06623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_16355_, _06621_, _23693_);
  or (_27153_, _16355_, _16354_);
  and (_16356_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  and (_16357_, _16061_, _23714_);
  or (_06948_, _16357_, _16356_);
  and (_16358_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_16359_, _02763_, _23983_);
  or (_06965_, _16359_, _16358_);
  and (_16360_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_16361_, _02763_, _24027_);
  or (_06971_, _16361_, _16360_);
  and (_16362_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_16363_, _15188_, _23919_);
  or (_06978_, _16363_, _16362_);
  or (_16364_, _23744_, _23211_);
  and (_16365_, _23284_, _23255_);
  nor (_16366_, _16365_, _23285_);
  or (_16367_, _16366_, _23210_);
  and (_16368_, _16367_, _23253_);
  and (_16369_, _16368_, _16364_);
  and (_16370_, _23252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_16371_, _16370_, _16369_);
  and (_06986_, _16371_, _22773_);
  and (_16372_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_16373_, _15188_, _23899_);
  or (_06992_, _16373_, _16372_);
  and (_16374_, _09463_, _23900_);
  and (_16375_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_07012_, _16375_, _16374_);
  and (_16376_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_16377_, _15188_, _23714_);
  or (_07017_, _16377_, _16376_);
  and (_16378_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  and (_16379_, _02756_, _24053_);
  or (_07023_, _16379_, _16378_);
  and (_16380_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  and (_16381_, _02756_, _23693_);
  or (_07031_, _16381_, _16380_);
  and (_16382_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nor (_16383_, _15189_, _24026_);
  or (_07035_, _16383_, _16382_);
  and (_16384_, _02758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  and (_16385_, _02756_, _23751_);
  or (_07039_, _16385_, _16384_);
  and (_16386_, _10273_, _23900_);
  and (_16387_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or (_07045_, _16387_, _16386_);
  and (_16388_, _07087_, _24053_);
  and (_16389_, _07089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_07061_, _16389_, _16388_);
  nand (_16390_, _02481_, _24017_);
  and (_16391_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_16392_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_16393_, _16392_, _16391_);
  or (_16394_, _16393_, _02481_);
  and (_16395_, _16394_, _05576_);
  and (_16396_, _16395_, _16390_);
  and (_16397_, _02473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_16398_, _16397_, _16396_);
  and (_07063_, _16398_, _22773_);
  and (_16399_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and (_16400_, _16292_, _23919_);
  or (_07065_, _16400_, _16399_);
  and (_16401_, _10273_, _23715_);
  and (_16402_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  or (_07070_, _16402_, _16401_);
  and (_16403_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  nor (_16404_, _16293_, _24026_);
  or (_07074_, _16404_, _16403_);
  and (_16405_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_16406_, _02763_, _23693_);
  or (_07099_, _16406_, _16405_);
  and (_16407_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_16408_, _02763_, _23751_);
  or (_27150_, _16408_, _16407_);
  and (_16409_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_16410_, _02763_, _24053_);
  or (_27149_, _16410_, _16409_);
  and (_16411_, _15189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_16412_, _15188_, _24052_);
  or (_26940_, _16412_, _16411_);
  and (_16413_, _05705_, _22895_);
  or (_16414_, _16413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_16415_, _16414_, _09813_);
  nand (_16416_, _16413_, _23681_);
  and (_16417_, _16416_, _16415_);
  and (_16418_, _05713_, _23744_);
  or (_16419_, _16418_, _16417_);
  and (_07143_, _16419_, _22773_);
  and (_16420_, _05705_, _24405_);
  or (_16421_, _16420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_16422_, _16421_, _09813_);
  nand (_16423_, _16420_, _23681_);
  and (_16424_, _16423_, _16422_);
  and (_16425_, _05713_, _24788_);
  or (_16426_, _16425_, _16424_);
  and (_07150_, _16426_, _22773_);
  and (_16427_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_16428_, _09579_, _23983_);
  or (_07153_, _16428_, _16427_);
  and (_16429_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_16430_, _09579_, _24027_);
  or (_07154_, _16430_, _16429_);
  or (_16431_, _23211_, _23205_);
  and (_16432_, _23364_, _23257_);
  nor (_16433_, _23376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand (_16434_, _16433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_16435_, _16434_, _16432_);
  nor (_16436_, _23364_, _23280_);
  and (_16437_, _23375_, _23373_);
  or (_16438_, _16437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_16439_, _16438_, _16436_);
  and (_16440_, _16439_, _16435_);
  or (_16441_, _16440_, _23210_);
  and (_16442_, _16441_, _23253_);
  and (_16443_, _16442_, _16431_);
  and (_16444_, _23252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_16445_, _16444_, _16443_);
  and (_07159_, _16445_, _22773_);
  and (_16446_, _02403_, _23983_);
  and (_16447_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_07161_, _16447_, _16446_);
  and (_16448_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_16449_, _02763_, _23900_);
  or (_07163_, _16449_, _16448_);
  not (_16450_, _05705_);
  or (_16451_, _16450_, _24426_);
  and (_16452_, _16451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_16453_, _16452_, _05713_);
  and (_16454_, _24432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_16455_, _16454_, _24431_);
  and (_16456_, _16455_, _05705_);
  or (_16457_, _16456_, _16453_);
  or (_16458_, _09813_, _23205_);
  and (_16459_, _16458_, _22773_);
  and (_07165_, _16459_, _16457_);
  and (_16460_, _10273_, _23693_);
  and (_16461_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or (_27217_, _16461_, _16460_);
  and (_16462_, _02476_, _05719_);
  or (_16463_, _16462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_16464_, _16463_, _05705_);
  nand (_16465_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_16466_, _16465_, _05705_);
  or (_16467_, _16466_, _03230_);
  and (_16468_, _16467_, _16464_);
  or (_16469_, _16468_, _05713_);
  nand (_16470_, _05713_, _24017_);
  and (_16471_, _16470_, _22773_);
  and (_07173_, _16471_, _16469_);
  and (_16472_, _24130_, _23924_);
  and (_16473_, _16472_, _24027_);
  not (_16474_, _16472_);
  and (_16475_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or (_07176_, _16475_, _16473_);
  and (_16476_, _05705_, _23208_);
  or (_16478_, _16476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_16479_, _16478_, _09813_);
  nand (_16480_, _16476_, _23681_);
  and (_16481_, _16480_, _16479_);
  nor (_16482_, _09813_, _23357_);
  or (_16483_, _16482_, _16481_);
  and (_07178_, _16483_, _22773_);
  and (_16484_, _05705_, _23250_);
  or (_16485_, _16484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_16486_, _16485_, _09813_);
  nand (_16487_, _16484_, _23681_);
  and (_16488_, _16487_, _16486_);
  and (_16489_, _05713_, _23413_);
  or (_16490_, _16489_, _16488_);
  and (_07180_, _16490_, _22773_);
  and (_16491_, _10273_, _23751_);
  and (_16492_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  or (_07182_, _16492_, _16491_);
  and (_16493_, _05662_, _05616_);
  and (_16494_, _16493_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_16495_, _16494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_16496_, _16495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_16497_, _16495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_16498_, _16497_, _16496_);
  and (_16499_, _05659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or (_16500_, _16499_, _05656_);
  or (_16501_, _16500_, _16498_);
  nand (_16502_, _05656_, _02475_);
  and (_16503_, _16502_, _05619_);
  and (_16504_, _16503_, _16501_);
  and (_16506_, _05618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_16507_, _16506_, _16504_);
  nor (_16508_, _05679_, _23357_);
  or (_16509_, _16508_, _16507_);
  and (_07204_, _16509_, _22773_);
  and (_16510_, _16472_, _24053_);
  and (_16511_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or (_07206_, _16511_, _16510_);
  and (_16512_, _05618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_16513_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_16514_, _16494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_16515_, _16514_, _16495_);
  and (_16516_, _05659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_16517_, _16516_, _05656_);
  or (_16518_, _16517_, _16515_);
  and (_16519_, _16518_, _16513_);
  and (_16520_, _16519_, _05619_);
  or (_16521_, _16520_, _16512_);
  and (_16522_, _05617_, _23205_);
  or (_16523_, _16522_, _16521_);
  and (_07209_, _16523_, _22773_);
  or (_16524_, _05682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_16525_, _16524_, _05679_);
  and (_16526_, _05617_, _23413_);
  or (_16527_, _16526_, _16525_);
  or (_16528_, _16493_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_16529_, _05656_, _16494_);
  and (_16530_, _16529_, _16528_);
  and (_16531_, _09797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_16532_, _16531_, _16530_);
  nand (_16533_, _16532_, _05619_);
  and (_16534_, _16533_, _22773_);
  and (_07211_, _16534_, _16527_);
  or (_16535_, _05679_, _23247_);
  or (_16536_, _05682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_16537_, _09797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_16538_, _05631_, _05616_);
  or (_16539_, _16538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_16540_, _05656_, _16493_);
  or (_16541_, _16540_, _05618_);
  and (_16542_, _16541_, _16539_);
  or (_16543_, _16542_, _16537_);
  and (_16544_, _16543_, _16536_);
  or (_16545_, _16544_, _05617_);
  and (_16546_, _16545_, _22773_);
  and (_07214_, _16546_, _16535_);
  and (_16547_, _05618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  not (_16548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nand (_16549_, _05656_, _16548_);
  and (_16550_, _05658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_16551_, _16550_, _05637_);
  not (_16552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_16553_, _05630_, _05616_);
  and (_16554_, _16553_, _16552_);
  nor (_16555_, _16554_, _16538_);
  or (_16556_, _16555_, _05656_);
  or (_16557_, _16556_, _16551_);
  and (_16558_, _16557_, _16549_);
  and (_16559_, _16558_, _05619_);
  or (_16560_, _16559_, _16547_);
  and (_16561_, _05617_, _23744_);
  or (_16562_, _16561_, _16560_);
  and (_07217_, _16562_, _22773_);
  or (_16563_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_16564_, _05658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_16565_, _16564_, _05637_);
  not (_16566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_16567_, _05687_, _16566_);
  and (_16568_, _16567_, _16553_);
  or (_16569_, _16568_, _05656_);
  or (_16570_, _16569_, _16565_);
  and (_16571_, _16570_, _16563_);
  and (_16572_, _16571_, _05619_);
  and (_16573_, _05618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_16574_, _05617_, _24788_);
  or (_16575_, _16574_, _16573_);
  or (_16576_, _16575_, _16572_);
  and (_07220_, _16576_, _22773_);
  and (_16577_, _24145_, _24130_);
  and (_16578_, _16577_, _23900_);
  not (_16579_, _16577_);
  and (_16580_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_07224_, _16580_, _16578_);
  and (_16581_, _02764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_16582_, _02763_, _23715_);
  or (_07227_, _16582_, _16581_);
  and (_16583_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nor (_16584_, _16066_, _24026_);
  or (_07229_, _16584_, _16583_);
  and (_16585_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  and (_16586_, _16292_, _24052_);
  or (_07231_, _16586_, _16585_);
  and (_16587_, _04033_, _23715_);
  and (_16588_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or (_07233_, _16588_, _16587_);
  and (_16589_, _24274_, _24130_);
  and (_16590_, _16589_, _23900_);
  not (_16591_, _16589_);
  and (_16592_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_07236_, _16592_, _16590_);
  and (_16593_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nor (_16594_, _16066_, _23982_);
  or (_07243_, _16594_, _16593_);
  and (_16595_, _24130_, _23905_);
  and (_16596_, _16595_, _23920_);
  not (_16597_, _16595_);
  and (_16598_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_07246_, _16598_, _16596_);
  and (_16599_, _08240_, _24027_);
  and (_16600_, _08242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_07248_, _16600_, _16599_);
  nand (_16601_, _24017_, _23210_);
  nor (_16602_, _10724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_16603_, _16602_, _10726_);
  or (_16604_, _16603_, _23210_);
  and (_16605_, _16604_, _25049_);
  and (_16606_, _16605_, _16601_);
  and (_16607_, _23252_, _22773_);
  and (_16608_, _16607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_07250_, _16608_, _16606_);
  and (_16609_, _16595_, _24053_);
  and (_16610_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or (_07252_, _16610_, _16609_);
  and (_16611_, _24130_, _23444_);
  and (_16612_, _16611_, _23900_);
  not (_16613_, _16611_);
  and (_16614_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or (_07256_, _16614_, _16612_);
  and (_16615_, _16611_, _24053_);
  and (_16616_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or (_07259_, _16616_, _16615_);
  nor (_16617_, _05682_, _24017_);
  or (_16618_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_16619_, _05627_, _05616_);
  not (_16620_, _16619_);
  nor (_16621_, _16620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_16622_, _16620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_16623_, _16622_, _05656_);
  or (_16624_, _16623_, _16621_);
  and (_16625_, _05659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_16626_, _16625_, _16624_);
  and (_16627_, _16626_, _16618_);
  and (_16628_, _16627_, _05619_);
  and (_16629_, _05617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_16630_, _16629_, _16628_);
  or (_16631_, _16630_, _16617_);
  and (_07261_, _16631_, _22773_);
  and (_16632_, _24130_, _23930_);
  and (_16633_, _16632_, _23983_);
  not (_16634_, _16632_);
  and (_16635_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_07264_, _16635_, _16633_);
  and (_16636_, _16632_, _23920_);
  and (_16637_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_07266_, _16637_, _16636_);
  nor (_16638_, _05682_, _23357_);
  and (_16639_, _05626_, _05616_);
  or (_16640_, _16639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_16641_, _16619_, _05656_);
  and (_16642_, _16641_, _16640_);
  and (_16643_, _09797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_16644_, _16643_, _16642_);
  and (_16645_, _16644_, _05619_);
  and (_16646_, _05617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_16647_, _16646_, _16645_);
  or (_16648_, _16647_, _16638_);
  and (_07269_, _16648_, _22773_);
  and (_16649_, _05618_, _23205_);
  and (_16650_, _05625_, _05616_);
  or (_16651_, _16650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_16652_, _16639_, _05656_);
  and (_16653_, _16652_, _16651_);
  and (_16654_, _09797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_16655_, _16654_, _16653_);
  and (_16656_, _16655_, _05619_);
  and (_16657_, _05617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_16658_, _16657_, _16656_);
  or (_16659_, _16658_, _16649_);
  and (_07271_, _16659_, _22773_);
  or (_16660_, _10723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_16661_, _16607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_16662_, _10724_);
  and (_16663_, _16662_, _25050_);
  or (_16664_, _16663_, _16661_);
  and (_16665_, _16664_, _16660_);
  nand (_16666_, _25049_, _23210_);
  nor (_16667_, _16666_, _23357_);
  or (_07273_, _16667_, _16665_);
  and (_16668_, _05618_, _23413_);
  and (_16669_, _05658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_16670_, _16669_, _05637_);
  not (_16671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_16672_, _09760_, _16671_);
  nor (_16673_, _16672_, _16650_);
  or (_16674_, _16673_, _05656_);
  or (_16675_, _16674_, _16670_);
  or (_16676_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_16677_, _16676_, _16675_);
  and (_16678_, _16677_, _05619_);
  and (_16679_, _05617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_16680_, _16679_, _16678_);
  or (_16681_, _16680_, _16668_);
  and (_07275_, _16681_, _22773_);
  and (_16682_, _24130_, _24108_);
  and (_16683_, _16682_, _23900_);
  not (_16684_, _16682_);
  and (_16685_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or (_07277_, _16685_, _16683_);
  and (_16686_, _16682_, _23693_);
  and (_16687_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or (_26890_, _16687_, _16686_);
  and (_16688_, _24157_, _24130_);
  and (_16689_, _16688_, _23983_);
  not (_16690_, _16688_);
  and (_16691_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_07282_, _16691_, _16689_);
  and (_16692_, _16688_, _23715_);
  and (_16693_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_07288_, _16693_, _16692_);
  and (_16694_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and (_16695_, _03165_, _23693_);
  or (_07292_, _16695_, _16694_);
  and (_16696_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  and (_16697_, _16292_, _23714_);
  or (_07295_, _16697_, _16696_);
  and (_16698_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  and (_16699_, _03165_, _23751_);
  or (_07299_, _16699_, _16698_);
  and (_16700_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and (_16701_, _16292_, _23692_);
  or (_07306_, _16701_, _16700_);
  nand (_16702_, _02473_, _24017_);
  and (_16703_, _05646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_16704_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_16705_, _16704_, _16703_);
  or (_16706_, _16705_, _02473_);
  and (_16707_, _16706_, _22773_);
  and (_07308_, _16707_, _16702_);
  and (_16708_, _16293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and (_16709_, _16292_, _23750_);
  or (_07310_, _16709_, _16708_);
  and (_16710_, _24130_, _24123_);
  and (_16711_, _16710_, _23693_);
  not (_16712_, _16710_);
  and (_16713_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or (_26889_, _16713_, _16711_);
  and (_16714_, _25169_, _23920_);
  and (_16715_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_07332_, _16715_, _16714_);
  and (_16716_, _09480_, _23983_);
  and (_16717_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or (_07335_, _16717_, _16716_);
  and (_16718_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  and (_16719_, _03165_, _24053_);
  or (_07337_, _16719_, _16718_);
  and (_16720_, _24130_, _24061_);
  and (_16721_, _16720_, _24027_);
  not (_16722_, _16720_);
  and (_16723_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_07341_, _16723_, _16721_);
  and (_16724_, _24098_, _23693_);
  and (_16725_, _24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or (_07344_, _16725_, _16724_);
  and (_16726_, _05618_, _23744_);
  and (_16727_, _05616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_16728_, _16727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor (_16729_, _09758_, _05656_);
  and (_16730_, _16729_, _16728_);
  and (_16731_, _09797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_16732_, _16731_, _16730_);
  and (_16733_, _16732_, _05619_);
  and (_16734_, _05617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_16735_, _16734_, _16733_);
  or (_16736_, _16735_, _16726_);
  and (_07345_, _16736_, _22773_);
  or (_16737_, _05616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_16738_, _05657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_16739_, _16738_, _05637_);
  nand (_16740_, _16739_, _16727_);
  and (_16741_, _16740_, _16737_);
  or (_16742_, _16741_, _05656_);
  or (_16743_, _05674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_16744_, _16743_, _16742_);
  and (_16745_, _16744_, _05619_);
  and (_16746_, _05618_, _24788_);
  and (_16747_, _05617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_16748_, _16747_, _16746_);
  or (_16749_, _16748_, _16745_);
  and (_07348_, _16749_, _22773_);
  and (_16750_, _16720_, _23751_);
  and (_16751_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_07350_, _16751_, _16750_);
  and (_16752_, _16720_, _23715_);
  and (_16753_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_07353_, _16753_, _16752_);
  and (_16754_, _15255_, _23693_);
  and (_16755_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or (_26907_, _16755_, _16754_);
  and (_16756_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_16757_, _16065_, _24052_);
  or (_07360_, _16757_, _16756_);
  and (_16758_, _16472_, _23693_);
  and (_16759_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or (_07363_, _16759_, _16758_);
  and (_16760_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  nor (_16761_, _15206_, _23982_);
  or (_07368_, _16761_, _16760_);
  and (_16762_, _16577_, _23751_);
  and (_16763_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_07371_, _16763_, _16762_);
  and (_16764_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  and (_16765_, _03165_, _23900_);
  or (_07374_, _16765_, _16764_);
  and (_16766_, _16589_, _23751_);
  and (_16767_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_07375_, _16767_, _16766_);
  or (_16768_, _05576_, _23247_);
  and (_16769_, _05646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_16770_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_16771_, _16770_, _16769_);
  or (_16772_, _16771_, _02473_);
  and (_16773_, _16772_, _22773_);
  and (_07378_, _16773_, _16768_);
  or (_16774_, _05576_, _23744_);
  nor (_16775_, _02482_, _16548_);
  and (_16776_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_16777_, _16776_, _16775_);
  or (_16778_, _16777_, _02473_);
  and (_16779_, _16778_, _22773_);
  and (_07380_, _16779_, _16774_);
  or (_16780_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_16781_, _02482_, _16566_);
  and (_16782_, _16781_, _16780_);
  or (_16783_, _16782_, _02473_);
  nand (_16784_, _02473_, _24047_);
  and (_16785_, _16784_, _22773_);
  and (_07385_, _16785_, _16783_);
  and (_16786_, _16595_, _23693_);
  and (_16787_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or (_07387_, _16787_, _16786_);
  and (_16788_, _03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  and (_16789_, _03165_, _23920_);
  or (_27147_, _16789_, _16788_);
  and (_16790_, _16682_, _24027_);
  and (_16791_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or (_26891_, _16791_, _16790_);
  and (_16792_, _25440_, _24053_);
  and (_16793_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or (_07395_, _16793_, _16792_);
  and (_16794_, _16688_, _23751_);
  and (_16795_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_07403_, _16795_, _16794_);
  and (_16796_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_16797_, _16065_, _23714_);
  or (_07405_, _16797_, _16796_);
  and (_16798_, _16066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_16799_, _16065_, _23692_);
  or (_07407_, _16799_, _16798_);
  and (_16800_, _16710_, _24027_);
  and (_16801_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or (_07409_, _16801_, _16800_);
  not (_16802_, _02481_);
  or (_16803_, _16802_, _23205_);
  and (_16804_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_16805_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_16806_, _16805_, _16804_);
  or (_16807_, _16806_, _02481_);
  and (_16808_, _16807_, _05576_);
  and (_16809_, _16808_, _16803_);
  and (_16810_, _02473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_16811_, _16810_, _16809_);
  and (_07412_, _16811_, _22773_);
  or (_16812_, _16802_, _23413_);
  and (_16813_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_16814_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_16815_, _16814_, _16813_);
  or (_16816_, _16815_, _02481_);
  and (_16817_, _16816_, _05576_);
  and (_16818_, _16817_, _16812_);
  and (_16819_, _02473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_16820_, _16819_, _16818_);
  and (_07414_, _16820_, _22773_);
  or (_16821_, _16802_, _23247_);
  and (_16822_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_16823_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_16824_, _16823_, _16822_);
  or (_16825_, _16824_, _02481_);
  and (_16826_, _16825_, _05576_);
  and (_16827_, _16826_, _16821_);
  and (_16828_, _02473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_16829_, _16828_, _16827_);
  and (_07417_, _16829_, _22773_);
  or (_16830_, _16802_, _23744_);
  and (_16831_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_16832_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_16833_, _16832_, _16831_);
  or (_16834_, _16833_, _02481_);
  and (_16835_, _16834_, _05576_);
  and (_16836_, _16835_, _16830_);
  and (_16837_, _02473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_16838_, _16837_, _16836_);
  and (_07420_, _16838_, _22773_);
  or (_16839_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_16840_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_16841_, _16840_, _16839_);
  or (_16842_, _16841_, _02481_);
  nand (_16843_, _02481_, _24047_);
  and (_16844_, _16843_, _16842_);
  or (_16845_, _16844_, _02473_);
  or (_16846_, _05576_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_16847_, _16846_, _22773_);
  and (_07439_, _16847_, _16845_);
  and (_16848_, _16632_, _23751_);
  and (_16849_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_07441_, _16849_, _16848_);
  and (_16850_, _16577_, _23920_);
  and (_16851_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_07446_, _16851_, _16850_);
  and (_16852_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and (_16853_, _03169_, _23900_);
  or (_07448_, _16853_, _16852_);
  and (_16854_, _16589_, _23920_);
  and (_16855_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_07450_, _16855_, _16854_);
  or (_16856_, _16156_, _26798_);
  not (_16857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_16858_, _16156_, _16857_);
  and (_16859_, _16858_, _22915_);
  and (_16860_, _16859_, _16856_);
  nor (_16861_, _22914_, _16857_);
  or (_16862_, _16156_, _23708_);
  and (_16863_, _16858_, _24330_);
  and (_16864_, _16863_, _16862_);
  or (_16865_, _16864_, _16861_);
  or (_16866_, _16865_, _16860_);
  and (_07452_, _16866_, _22773_);
  and (_16867_, _16595_, _24027_);
  and (_16868_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or (_07454_, _16868_, _16867_);
  and (_16869_, _16611_, _23751_);
  and (_16870_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or (_26895_, _16870_, _16869_);
  or (_16871_, _16156_, _00183_);
  not (_16872_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_16873_, _16156_, _16872_);
  and (_16874_, _16873_, _22915_);
  and (_16875_, _16874_, _16871_);
  nor (_16876_, _22914_, _16872_);
  and (_16877_, _16155_, _24184_);
  nand (_16878_, _16877_, _23681_);
  or (_16879_, _16877_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_16880_, _16879_, _24330_);
  and (_16881_, _16880_, _16878_);
  or (_16882_, _16881_, _16876_);
  or (_16883_, _16882_, _16875_);
  and (_07458_, _16883_, _22773_);
  or (_16884_, _16156_, _00101_);
  not (_16885_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_16886_, _16156_, _16885_);
  and (_16887_, _16886_, _22915_);
  and (_16888_, _16887_, _16884_);
  nor (_16889_, _22914_, _16885_);
  and (_16890_, _16155_, _22895_);
  nand (_16891_, _16890_, _23681_);
  or (_16892_, _16890_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_16893_, _16892_, _24330_);
  and (_16894_, _16893_, _16891_);
  or (_16895_, _16894_, _16889_);
  or (_16896_, _16895_, _16888_);
  and (_07460_, _16896_, _22773_);
  or (_16897_, _16156_, _00443_);
  nand (_16898_, _16156_, _03530_);
  and (_16899_, _16898_, _22915_);
  and (_16900_, _16899_, _16897_);
  nor (_16901_, _22914_, _03530_);
  and (_16902_, _16155_, _23208_);
  nand (_16903_, _16902_, _23681_);
  or (_16904_, _16902_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_16905_, _16904_, _24330_);
  and (_16906_, _16905_, _16903_);
  or (_16907_, _16906_, _16901_);
  or (_16908_, _16907_, _16900_);
  and (_07462_, _16908_, _22773_);
  or (_16909_, _16156_, _00352_);
  nand (_16910_, _16156_, _03525_);
  and (_16911_, _16910_, _22915_);
  and (_16912_, _16911_, _16909_);
  nor (_16913_, _22914_, _03525_);
  and (_16914_, _16155_, _24190_);
  nand (_16915_, _16914_, _23681_);
  or (_16916_, _16914_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_16917_, _16916_, _24330_);
  and (_16918_, _16917_, _16915_);
  or (_16919_, _16918_, _16913_);
  or (_16920_, _16919_, _16912_);
  and (_07464_, _16920_, _22773_);
  or (_16921_, _16156_, _00277_);
  not (_16922_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_16923_, _16156_, _16922_);
  and (_16924_, _16923_, _22915_);
  and (_16925_, _16924_, _16921_);
  nor (_16926_, _22914_, _16922_);
  and (_16927_, _16155_, _23250_);
  nand (_16928_, _16927_, _23681_);
  or (_16929_, _16927_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_16930_, _16929_, _24330_);
  and (_16931_, _16930_, _16928_);
  or (_16932_, _16931_, _16926_);
  or (_16933_, _16932_, _16925_);
  and (_07466_, _16933_, _22773_);
  and (_16934_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_16935_, _15205_, _23750_);
  or (_07468_, _16935_, _16934_);
  or (_16936_, _16156_, _00564_);
  nand (_16937_, _16156_, _03517_);
  and (_16938_, _16937_, _22915_);
  and (_16939_, _16938_, _16936_);
  nor (_16940_, _22914_, _03517_);
  and (_16941_, _16155_, _24373_);
  nand (_16942_, _16941_, _23681_);
  or (_16943_, _16941_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_16944_, _16943_, _24330_);
  and (_16945_, _16944_, _16942_);
  or (_16946_, _16945_, _16940_);
  or (_16947_, _16946_, _16939_);
  and (_07470_, _16947_, _22773_);
  and (_16948_, _16710_, _23715_);
  and (_16949_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or (_07473_, _16949_, _16948_);
  and (_16950_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_16951_, _15205_, _24052_);
  or (_07475_, _16951_, _16950_);
  and (_16952_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and (_16953_, _03169_, _23715_);
  or (_07477_, _16953_, _16952_);
  and (_16954_, _09480_, _24027_);
  and (_16955_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or (_27042_, _16955_, _16954_);
  and (_16956_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  and (_16957_, _03169_, _23693_);
  or (_07480_, _16957_, _16956_);
  and (_16958_, _16611_, _23983_);
  and (_16959_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or (_07486_, _16959_, _16958_);
  and (_16960_, _16632_, _23693_);
  and (_16961_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_26893_, _16961_, _16960_);
  and (_16962_, _16589_, _24027_);
  and (_16963_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_07493_, _16963_, _16962_);
  and (_16964_, _02244_, _23693_);
  and (_16965_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or (_07499_, _16965_, _16964_);
  and (_16966_, _10273_, _24027_);
  and (_16967_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  or (_07503_, _16967_, _16966_);
  and (_16968_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_16969_, _15205_, _23714_);
  or (_07508_, _16969_, _16968_);
  and (_16970_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_16971_, _15205_, _23919_);
  or (_07510_, _16971_, _16970_);
  and (_16972_, _15206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_16973_, _15205_, _23899_);
  or (_07514_, _16973_, _16972_);
  and (_16974_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and (_16975_, _03169_, _23983_);
  or (_07533_, _16975_, _16974_);
  and (_16976_, _02326_, _23920_);
  and (_16977_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or (_07535_, _16977_, _16976_);
  and (_16978_, _04771_, _23983_);
  and (_16979_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or (_07540_, _16979_, _16978_);
  and (_16980_, _04771_, _24053_);
  and (_16981_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_27248_, _16981_, _16980_);
  and (_16982_, _03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and (_16983_, _03169_, _24027_);
  or (_07544_, _16983_, _16982_);
  and (_16984_, _24027_, _23925_);
  and (_16985_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_07546_, _16985_, _16984_);
  and (_16986_, _05731_, _24053_);
  and (_16987_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or (_27241_, _16987_, _16986_);
  and (_16988_, _24108_, _23891_);
  and (_16989_, _16988_, _24053_);
  not (_16990_, _16988_);
  and (_16991_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_07559_, _16991_, _16989_);
  and (_16992_, _24157_, _23891_);
  and (_16993_, _16992_, _23715_);
  not (_16994_, _16992_);
  and (_16995_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or (_07562_, _16995_, _16993_);
  and (_16996_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and (_16997_, _15209_, _24052_);
  or (_07565_, _16997_, _16996_);
  and (_16998_, _24123_, _23891_);
  and (_17000_, _16998_, _24027_);
  not (_17001_, _16998_);
  and (_17002_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_07570_, _17002_, _17000_);
  and (_17003_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and (_17004_, _15209_, _23750_);
  or (_07572_, _17004_, _17003_);
  and (_17005_, _16998_, _23751_);
  and (_17006_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_07575_, _17006_, _17005_);
  and (_17007_, _23892_, _23693_);
  and (_17008_, _23902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or (_07577_, _17008_, _17007_);
  and (_17009_, _24069_, _23693_);
  and (_17010_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or (_07579_, _17010_, _17009_);
  and (_17011_, _01759_, _23693_);
  and (_17012_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  or (_07586_, _17012_, _17011_);
  and (_17013_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_17014_, _02769_, _24027_);
  or (_27145_, _17014_, _17013_);
  and (_17015_, _15246_, _23715_);
  and (_17016_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_07591_, _17016_, _17015_);
  and (_17017_, _24145_, _23453_);
  and (_17018_, _17017_, _23751_);
  not (_17019_, _17017_);
  and (_17020_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_07595_, _17020_, _17018_);
  and (_17021_, _04033_, _23693_);
  and (_17022_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or (_07596_, _17022_, _17021_);
  and (_17023_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_17024_, _02769_, _23920_);
  or (_07603_, _17024_, _17023_);
  and (_17025_, _02248_, _23751_);
  and (_17026_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or (_07606_, _17026_, _17025_);
  and (_17027_, _01759_, _23900_);
  and (_17028_, _01761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  or (_07608_, _17028_, _17027_);
  and (_17029_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and (_17030_, _15209_, _23692_);
  or (_07611_, _17030_, _17029_);
  and (_17031_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and (_17032_, _15209_, _23919_);
  or (_07613_, _17032_, _17031_);
  and (_17033_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and (_17034_, _15209_, _23899_);
  or (_07641_, _17034_, _17033_);
  and (_17035_, _02423_, _23751_);
  and (_17036_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or (_07643_, _17036_, _17035_);
  and (_17037_, _25428_, _23693_);
  and (_17038_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_27197_, _17038_, _17037_);
  and (_07647_, _26125_, _22773_);
  and (_17039_, _24319_, _23920_);
  and (_17040_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_07649_, _17040_, _17039_);
  and (_07651_, _26880_, _26021_);
  and (_17041_, _24319_, _23751_);
  and (_17042_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_07654_, _17042_, _17041_);
  and (_17043_, _15210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  and (_17044_, _15209_, _23714_);
  or (_07657_, _17044_, _17043_);
  and (_17045_, _16998_, _24053_);
  and (_17046_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_07662_, _17046_, _17045_);
  and (_17047_, _02853_, _23715_);
  and (_17048_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or (_07664_, _17048_, _17047_);
  and (_17049_, _01952_, _23920_);
  and (_17050_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or (_07667_, _17050_, _17049_);
  and (_17051_, _23715_, _23454_);
  and (_17052_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or (_07673_, _17052_, _17051_);
  and (_17053_, _24062_, _23983_);
  and (_17054_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_07679_, _17054_, _17053_);
  and (_17055_, _24062_, _23900_);
  and (_17056_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_07682_, _17056_, _17055_);
  and (_17057_, _23932_, _23900_);
  and (_17058_, _23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_27210_, _17058_, _17057_);
  and (_17059_, _23987_, _23890_);
  and (_17060_, _17059_, _23983_);
  not (_17061_, _17059_);
  and (_17062_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_27258_, _17062_, _17060_);
  and (_17063_, _10669_, _24097_);
  not (_17064_, _17063_);
  and (_17065_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  and (_17066_, _17063_, _23714_);
  or (_07688_, _17066_, _17065_);
  and (_17067_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and (_17068_, _17063_, _23692_);
  or (_07692_, _17068_, _17067_);
  and (_17069_, _24097_, _23987_);
  and (_17070_, _17069_, _23715_);
  not (_17071_, _17069_);
  and (_17072_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_07695_, _17072_, _17070_);
  and (_17073_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  and (_17074_, _17063_, _23750_);
  or (_07696_, _17074_, _17073_);
  and (_17075_, _23988_, _23715_);
  and (_17076_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_07700_, _17076_, _17075_);
  and (_17077_, _02244_, _23983_);
  and (_17078_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or (_07702_, _17078_, _17077_);
  and (_17079_, _09552_, _23715_);
  and (_17080_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_07705_, _17080_, _17079_);
  and (_17081_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  and (_17082_, _17063_, _24052_);
  or (_07707_, _17082_, _17081_);
  and (_17083_, _24061_, _23891_);
  and (_17084_, _17083_, _23983_);
  not (_17085_, _17083_);
  and (_17086_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or (_07710_, _17086_, _17084_);
  and (_17087_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_17088_, _02769_, _23983_);
  or (_07716_, _17088_, _17087_);
  and (_17089_, _25482_, _23751_);
  and (_17090_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_27226_, _17090_, _17089_);
  and (_17091_, _02455_, _23715_);
  and (_17092_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or (_07719_, _17092_, _17091_);
  and (_17093_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  nor (_17094_, _17064_, _23982_);
  or (_07742_, _17094_, _17093_);
  and (_17095_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  nor (_17096_, _17064_, _24026_);
  or (_07744_, _17096_, _17095_);
  and (_17097_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  and (_17098_, _17063_, _23919_);
  or (_07748_, _17098_, _17097_);
  and (_17099_, _24274_, _23453_);
  and (_17100_, _17099_, _23900_);
  not (_17101_, _17099_);
  and (_17102_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_07751_, _17102_, _17100_);
  and (_17103_, _17064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and (_17104_, _17063_, _23899_);
  or (_07763_, _17104_, _17103_);
  and (_17105_, _09507_, _23920_);
  and (_17106_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_07765_, _17106_, _17105_);
  and (_17107_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_17108_, _02769_, _24053_);
  or (_07767_, _17108_, _17107_);
  and (_17109_, _25428_, _23983_);
  and (_17110_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_27198_, _17110_, _17109_);
  and (_17111_, _24069_, _24027_);
  and (_17112_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or (_07784_, _17112_, _17111_);
  and (_17113_, _25159_, _23900_);
  and (_17114_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or (_27193_, _17114_, _17113_);
  and (_17115_, _25190_, _23715_);
  and (_17116_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_07801_, _17116_, _17115_);
  and (_17117_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_17118_, _16276_, _23714_);
  or (_07803_, _17118_, _17117_);
  and (_17119_, _01952_, _23751_);
  and (_17120_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or (_07805_, _17120_, _17119_);
  and (_17121_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_17122_, _16276_, _23692_);
  or (_08024_, _17122_, _17121_);
  and (_17123_, _09621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  and (_17124_, _09620_, _24053_);
  or (_08026_, _17124_, _17123_);
  and (_17125_, _16988_, _23751_);
  and (_17126_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_08029_, _17126_, _17125_);
  and (_17127_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_17128_, _02769_, _23715_);
  or (_08036_, _17128_, _17127_);
  and (_17129_, _17017_, _24027_);
  and (_17130_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_08039_, _17130_, _17129_);
  and (_17131_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_17132_, _16276_, _23919_);
  or (_08041_, _17132_, _17131_);
  and (_17133_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  nor (_17134_, _16277_, _23982_);
  or (_08044_, _17134_, _17133_);
  and (_17135_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_17136_, _02769_, _23693_);
  or (_27143_, _17136_, _17135_);
  and (_17137_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  nor (_17138_, _16277_, _24026_);
  or (_08047_, _17138_, _17137_);
  and (_17139_, _10525_, _23715_);
  and (_17140_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or (_08050_, _17140_, _17139_);
  and (_17141_, _24319_, _24027_);
  and (_17142_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_08051_, _17142_, _17141_);
  and (_17143_, _02771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_17144_, _02769_, _23751_);
  or (_08055_, _17144_, _17143_);
  and (_17145_, _16988_, _23693_);
  and (_17146_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_08110_, _17146_, _17145_);
  and (_17147_, _24235_, _24124_);
  and (_17148_, _17147_, _23900_);
  not (_17149_, _17147_);
  and (_17150_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_08116_, _17150_, _17148_);
  and (_17151_, _24124_, _23890_);
  and (_17152_, _17151_, _23920_);
  not (_17153_, _17151_);
  and (_17154_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_08123_, _17154_, _17152_);
  and (_17155_, _17151_, _23751_);
  and (_17156_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or (_08125_, _17156_, _17155_);
  and (_17157_, _24124_, _24097_);
  and (_17158_, _17157_, _24027_);
  not (_17159_, _17157_);
  and (_17160_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or (_08129_, _17160_, _17158_);
  and (_17161_, _17157_, _23693_);
  and (_17162_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or (_08132_, _17162_, _17161_);
  and (_17163_, _24124_, _24068_);
  and (_17164_, _17163_, _23983_);
  not (_17165_, _17163_);
  and (_17166_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_27290_, _17166_, _17164_);
  and (_17167_, _17163_, _23693_);
  and (_17168_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_08136_, _17168_, _17167_);
  and (_17169_, _24124_, _23700_);
  and (_17170_, _17169_, _23983_);
  not (_17171_, _17169_);
  and (_17172_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_08139_, _17172_, _17170_);
  and (_17173_, _17169_, _23715_);
  and (_17174_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_08142_, _17174_, _17173_);
  and (_17175_, _09580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_17176_, _09579_, _23920_);
  or (_26956_, _17176_, _17175_);
  and (_17177_, _24124_, _23938_);
  and (_17178_, _17177_, _23920_);
  not (_17179_, _17177_);
  and (_17180_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_08148_, _17180_, _17178_);
  and (_17182_, _17177_, _23751_);
  and (_17183_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or (_08150_, _17183_, _17182_);
  and (_17184_, _23987_, _23924_);
  and (_17185_, _17184_, _24027_);
  not (_17186_, _17184_);
  and (_17187_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or (_08154_, _17187_, _17185_);
  and (_17188_, _10525_, _23693_);
  and (_17189_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or (_08156_, _17189_, _17188_);
  and (_17190_, _24274_, _23987_);
  and (_17191_, _17190_, _23920_);
  not (_17192_, _17190_);
  and (_17193_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_08160_, _17193_, _17191_);
  and (_17194_, _17190_, _23715_);
  and (_17195_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_08162_, _17195_, _17194_);
  and (_17196_, _23987_, _23905_);
  and (_17197_, _17196_, _23983_);
  not (_17198_, _17196_);
  and (_17199_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or (_08166_, _17199_, _17197_);
  and (_17200_, _17196_, _23715_);
  and (_17201_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_27279_, _17201_, _17200_);
  and (_17202_, _17196_, _23751_);
  and (_17203_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_08169_, _17203_, _17202_);
  and (_17204_, _24215_, _23900_);
  and (_17205_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_08172_, _17205_, _17204_);
  and (_17206_, _17184_, _23751_);
  and (_17207_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_27283_, _17207_, _17206_);
  and (_17208_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  nor (_17209_, _16271_, _23982_);
  or (_08386_, _17209_, _17208_);
  and (_17210_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nor (_17211_, _16271_, _24026_);
  or (_08389_, _17211_, _17210_);
  and (_17212_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_17213_, _16270_, _23919_);
  or (_08392_, _17213_, _17212_);
  and (_17214_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_17215_, _16270_, _23899_);
  or (_08394_, _17215_, _17214_);
  and (_17216_, _24145_, _23987_);
  and (_17217_, _17216_, _23693_);
  not (_17218_, _17216_);
  and (_17219_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_08398_, _17219_, _17217_);
  and (_17220_, _17216_, _23920_);
  and (_17221_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_08399_, _17221_, _17220_);
  and (_17222_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_17223_, _02775_, _23715_);
  or (_08403_, _17223_, _17222_);
  and (_17224_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_17225_, _02775_, _23693_);
  or (_08406_, _17225_, _17224_);
  and (_17226_, _17147_, _24027_);
  and (_17227_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_27293_, _17227_, _17226_);
  and (_17228_, _17147_, _24053_);
  and (_17229_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_27292_, _17229_, _17228_);
  and (_17230_, _23983_, _23721_);
  and (_17231_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_08412_, _17231_, _17230_);
  and (_17232_, _16277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_17233_, _16276_, _24052_);
  or (_08414_, _17233_, _17232_);
  and (_17234_, _17169_, _24053_);
  and (_17235_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_08420_, _17235_, _17234_);
  and (_17236_, _10341_, _23983_);
  and (_17237_, _10343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_08554_, _17237_, _17236_);
  and (_17238_, _01908_, _24053_);
  and (_17239_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or (_08577_, _17239_, _17238_);
  and (_17240_, _01908_, _23751_);
  and (_17241_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or (_08593_, _17241_, _17240_);
  and (_17242_, _24319_, _24053_);
  and (_17243_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_08604_, _17243_, _17242_);
  and (_17244_, _01932_, _23983_);
  and (_17245_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_08617_, _17245_, _17244_);
  and (_17246_, _24235_, _23453_);
  and (_17247_, _17246_, _23751_);
  not (_17248_, _17246_);
  and (_17249_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or (_27199_, _17249_, _17247_);
  and (_17250_, _04033_, _24053_);
  and (_17251_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or (_08649_, _17251_, _17250_);
  nor (_26831_[5], _24495_, rst);
  and (_17252_, _02403_, _23900_);
  and (_17253_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_08663_, _17253_, _17252_);
  and (_17254_, _02403_, _23715_);
  and (_17255_, _02405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_08667_, _17255_, _17254_);
  and (_26831_[4], _24664_, _22773_);
  and (_17256_, _02509_, _24053_);
  and (_17257_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_08685_, _17257_, _17256_);
  and (_17258_, _02509_, _23751_);
  and (_17259_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_08702_, _17259_, _17258_);
  and (_17260_, _17246_, _24053_);
  and (_17261_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or (_08707_, _17261_, _17260_);
  and (_17262_, _04771_, _23751_);
  and (_17263_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_27249_, _17263_, _17262_);
  and (_17264_, _04771_, _23693_);
  and (_17265_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_27250_, _17265_, _17264_);
  and (_17266_, _04771_, _23715_);
  and (_17267_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_08729_, _17267_, _17266_);
  and (_17268_, _04207_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_17269_, _04231_, _24725_);
  or (_17270_, _17269_, _24675_);
  and (_17271_, _04210_, _24566_);
  or (_17272_, _17271_, _06146_);
  or (_17273_, _17272_, _17270_);
  or (_17274_, _17273_, _04236_);
  or (_17275_, _17274_, _06143_);
  and (_17276_, _17275_, _01886_);
  or (_26838_[1], _17276_, _17268_);
  and (_17277_, _25924_, _24672_);
  or (_17278_, _17277_, _05791_);
  or (_17279_, _17278_, _24710_);
  and (_17280_, _25876_, _24615_);
  or (_17281_, _17280_, _05442_);
  or (_17282_, _17281_, _17279_);
  or (_17283_, _06310_, _06146_);
  or (_17284_, _17283_, _17282_);
  or (_17285_, _17284_, _05466_);
  or (_17286_, _17285_, _05437_);
  and (_17287_, _17286_, _23760_);
  and (_17288_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17289_, _17288_, _05455_);
  or (_17290_, _17289_, _17287_);
  and (_26844_, _17290_, _22773_);
  and (_17291_, _01250_, _01127_);
  and (_17292_, _01221_, _24610_);
  and (_17293_, _01144_, _01139_);
  or (_17294_, _17293_, _17292_);
  or (_17295_, _17294_, _17291_);
  or (_17296_, _01281_, _01235_);
  or (_17297_, _17296_, _01264_);
  or (_17298_, _17297_, _17295_);
  nand (_17299_, _01261_, _01194_);
  or (_17300_, _17299_, _17298_);
  and (_17301_, _01215_, _01156_);
  or (_17302_, _01250_, _01136_);
  or (_17303_, _17302_, _01118_);
  and (_17304_, _17303_, _01122_);
  or (_17305_, _17304_, _07873_);
  or (_17306_, _17305_, _17301_);
  or (_17307_, _17306_, _07872_);
  or (_17308_, _17307_, _17300_);
  and (_17309_, _17308_, _23761_);
  nor (_17310_, _07866_, _04965_);
  or (_17311_, _17310_, rst);
  or (_26834_[1], _17311_, _17309_);
  and (_17312_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17313_, _17312_, _05450_);
  and (_17314_, _17313_, _22773_);
  or (_17315_, _04231_, _24691_);
  or (_17316_, _17280_, _05771_);
  or (_17317_, _17316_, _17315_);
  or (_17318_, _17317_, _24675_);
  and (_17319_, _17318_, _01886_);
  or (_26837_[1], _17319_, _17314_);
  and (_17320_, _04207_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_17321_, _25914_, _25898_);
  or (_17322_, _17321_, _25875_);
  or (_17323_, _06057_, _25920_);
  or (_17324_, _17323_, _17322_);
  or (_17325_, _06061_, _06048_);
  or (_17326_, _17325_, _17280_);
  or (_17327_, _17326_, _06068_);
  or (_17328_, _17327_, _17324_);
  and (_17329_, _17328_, _01886_);
  or (_26841_[1], _17329_, _17320_);
  or (_17330_, _06603_, _04210_);
  and (_17331_, _17330_, _23760_);
  nor (_17332_, _25859_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_17333_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17334_, _17333_, _17332_);
  or (_17335_, _17334_, _17331_);
  and (_26843_[1], _17335_, _22773_);
  and (_17336_, _24319_, _23693_);
  and (_17337_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_08790_, _17337_, _17336_);
  and (_17338_, _02423_, _24053_);
  and (_17339_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or (_08812_, _17339_, _17338_);
  and (_17340_, _17059_, _23751_);
  and (_17341_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_08817_, _17341_, _17340_);
  and (_17342_, _02853_, _23920_);
  and (_17343_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or (_27133_, _17343_, _17342_);
  and (_17344_, _17246_, _23983_);
  and (_17345_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or (_27200_, _17345_, _17344_);
  and (_17346_, _01908_, _23983_);
  and (_17347_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or (_08854_, _17347_, _17346_);
  and (_17348_, _01908_, _24027_);
  and (_17349_, _01910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or (_27033_, _17349_, _17348_);
  and (_17350_, _10273_, _23920_);
  and (_17351_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or (_08884_, _17351_, _17350_);
  and (_17352_, _10411_, _23920_);
  and (_17353_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or (_08886_, _17353_, _17352_);
  and (_17354_, _17190_, _24053_);
  and (_17355_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_08912_, _17355_, _17354_);
  and (_17356_, _17196_, _23920_);
  and (_17357_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or (_08914_, _17357_, _17356_);
  and (_17358_, _24215_, _23983_);
  and (_17359_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_08917_, _17359_, _17358_);
  and (_17360_, _17184_, _23715_);
  and (_17361_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_08920_, _17361_, _17360_);
  and (_17362_, _17151_, _23693_);
  and (_17363_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or (_08925_, _17363_, _17362_);
  and (_17364_, _17157_, _23715_);
  and (_17365_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or (_08927_, _17365_, _17364_);
  and (_17366_, _17163_, _23715_);
  and (_17367_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_27289_, _17367_, _17366_);
  and (_17368_, _17169_, _23900_);
  and (_17369_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_08930_, _17369_, _17368_);
  and (_17370_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_17371_, _02775_, _23920_);
  or (_08934_, _17371_, _17370_);
  and (_17372_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_17373_, _02775_, _23900_);
  or (_27141_, _17373_, _17372_);
  and (_17374_, _10411_, _24027_);
  and (_17375_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or (_08938_, _17375_, _17374_);
  and (_17376_, _24053_, _23721_);
  and (_17377_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_08950_, _17377_, _17376_);
  and (_17378_, _17059_, _23693_);
  and (_17379_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_08963_, _17379_, _17378_);
  and (_17380_, _17163_, _23900_);
  and (_17381_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_08973_, _17381_, _17380_);
  and (_17382_, _16264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  and (_17383_, _16263_, _23983_);
  or (_08979_, _17383_, _17382_);
  and (_17384_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_17385_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_17386_, _17385_, _17384_);
  and (_17387_, _17386_, _04832_);
  and (_17388_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_17389_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_17390_, _17389_, _17388_);
  and (_17391_, _17390_, _10928_);
  or (_17392_, _17391_, _17387_);
  or (_17393_, _17392_, _10926_);
  and (_17394_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and (_17395_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_17396_, _17395_, _17394_);
  and (_17397_, _17396_, _04832_);
  and (_17398_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_17399_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_17400_, _17399_, _17398_);
  and (_17401_, _17400_, _10928_);
  or (_17402_, _17401_, _17397_);
  or (_17403_, _17402_, _04868_);
  and (_17404_, _17403_, _10945_);
  and (_17405_, _17404_, _17393_);
  or (_17406_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_17407_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_17408_, _17407_, _17406_);
  and (_17409_, _17408_, _04832_);
  or (_17410_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_17411_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_17412_, _17411_, _17410_);
  and (_17413_, _17412_, _10928_);
  or (_17414_, _17413_, _17409_);
  or (_17415_, _17414_, _10926_);
  or (_17416_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_17417_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_17418_, _17417_, _17416_);
  and (_17419_, _17418_, _04832_);
  or (_17420_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_17421_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and (_17422_, _17421_, _17420_);
  and (_17423_, _17422_, _10928_);
  or (_17424_, _17423_, _17419_);
  or (_17425_, _17424_, _04868_);
  and (_17426_, _17425_, _04859_);
  and (_17427_, _17426_, _17415_);
  or (_17428_, _17427_, _17405_);
  and (_17429_, _17428_, _04849_);
  and (_17430_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_17431_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_17432_, _17431_, _17430_);
  and (_17433_, _17432_, _04832_);
  and (_17434_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_17435_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_17436_, _17435_, _17434_);
  and (_17437_, _17436_, _10928_);
  or (_17438_, _17437_, _17433_);
  or (_17439_, _17438_, _10926_);
  and (_17440_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_17441_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_17442_, _17441_, _17440_);
  and (_17443_, _17442_, _04832_);
  and (_17444_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_17445_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_17446_, _17445_, _17444_);
  and (_17447_, _17446_, _10928_);
  or (_17448_, _17447_, _17443_);
  or (_17449_, _17448_, _04868_);
  and (_17450_, _17449_, _10945_);
  and (_17451_, _17450_, _17439_);
  or (_17452_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_17453_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_17454_, _17453_, _10928_);
  and (_17455_, _17454_, _17452_);
  or (_17456_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_17457_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_17458_, _17457_, _04832_);
  and (_17459_, _17458_, _17456_);
  or (_17460_, _17459_, _17455_);
  or (_17461_, _17460_, _10926_);
  or (_17462_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_17463_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and (_17464_, _17463_, _10928_);
  and (_17465_, _17464_, _17462_);
  or (_17466_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_17467_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and (_17468_, _17467_, _04832_);
  and (_17469_, _17468_, _17466_);
  or (_17470_, _17469_, _17465_);
  or (_17471_, _17470_, _04868_);
  and (_17472_, _17471_, _04859_);
  and (_17473_, _17472_, _17461_);
  or (_17474_, _17473_, _17451_);
  and (_17475_, _17474_, _10997_);
  or (_17476_, _17475_, _17429_);
  and (_17477_, _17476_, _10996_);
  and (_17478_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_17479_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_17480_, _17479_, _17478_);
  and (_17481_, _17480_, _04832_);
  and (_17482_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_17483_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_17484_, _17483_, _17482_);
  and (_17485_, _17484_, _10928_);
  or (_17486_, _17485_, _17481_);
  and (_17487_, _17486_, _04868_);
  and (_17488_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_17489_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_17490_, _17489_, _17488_);
  and (_17491_, _17490_, _04832_);
  and (_17492_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_17493_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_17494_, _17493_, _17492_);
  and (_17495_, _17494_, _10928_);
  or (_17496_, _17495_, _17491_);
  and (_17497_, _17496_, _10926_);
  or (_17498_, _17497_, _17487_);
  and (_17499_, _17498_, _10945_);
  or (_17500_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_17501_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_17502_, _17501_, _10928_);
  and (_17503_, _17502_, _17500_);
  or (_17504_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_17505_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_17506_, _17505_, _04832_);
  and (_17507_, _17506_, _17504_);
  or (_17508_, _17507_, _17503_);
  and (_17509_, _17508_, _04868_);
  or (_17510_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_17512_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_17513_, _17512_, _10928_);
  and (_17514_, _17513_, _17510_);
  or (_17515_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_17516_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_17517_, _17516_, _04832_);
  and (_17518_, _17517_, _17515_);
  or (_17519_, _17518_, _17514_);
  and (_17520_, _17519_, _10926_);
  or (_17521_, _17520_, _17509_);
  and (_17522_, _17521_, _04859_);
  or (_17523_, _17522_, _17499_);
  and (_17524_, _17523_, _10997_);
  and (_17525_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_17526_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_17527_, _17526_, _17525_);
  and (_17528_, _17527_, _04832_);
  and (_17529_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_17530_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_17531_, _17530_, _17529_);
  and (_17532_, _17531_, _10928_);
  or (_17533_, _17532_, _17528_);
  and (_17534_, _17533_, _04868_);
  and (_17535_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and (_17536_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_17537_, _17536_, _17535_);
  and (_17538_, _17537_, _04832_);
  and (_17539_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_17540_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_17541_, _17540_, _17539_);
  and (_17542_, _17541_, _10928_);
  or (_17543_, _17542_, _17538_);
  and (_17544_, _17543_, _10926_);
  or (_17545_, _17544_, _17534_);
  and (_17546_, _17545_, _10945_);
  or (_17547_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_17548_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_17549_, _17548_, _17547_);
  and (_17550_, _17549_, _04832_);
  or (_17551_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_17552_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_17553_, _17552_, _17551_);
  and (_17554_, _17553_, _10928_);
  or (_17555_, _17554_, _17550_);
  and (_17556_, _17555_, _04868_);
  or (_17557_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_17558_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_17559_, _17558_, _17557_);
  and (_17560_, _17559_, _04832_);
  or (_17561_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_17563_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_17564_, _17563_, _17561_);
  and (_17565_, _17564_, _10928_);
  or (_17566_, _17565_, _17560_);
  and (_17567_, _17566_, _10926_);
  or (_17568_, _17567_, _17556_);
  and (_17569_, _17568_, _04859_);
  or (_17570_, _17569_, _17546_);
  and (_17571_, _17570_, _04849_);
  or (_17572_, _17571_, _17524_);
  and (_17573_, _17572_, _04839_);
  or (_17574_, _17573_, _17477_);
  or (_17575_, _17574_, _04843_);
  and (_17576_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and (_17577_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_17578_, _17577_, _17576_);
  and (_17579_, _17578_, _04832_);
  and (_17580_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_17581_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_17582_, _17581_, _17580_);
  and (_17584_, _17582_, _10928_);
  or (_17585_, _17584_, _17579_);
  or (_17586_, _17585_, _10926_);
  and (_17587_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and (_17588_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_17589_, _17588_, _17587_);
  and (_17590_, _17589_, _04832_);
  and (_17591_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_17592_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_17593_, _17592_, _17591_);
  and (_17594_, _17593_, _10928_);
  or (_17595_, _17594_, _17590_);
  or (_17596_, _17595_, _04868_);
  and (_17597_, _17596_, _10945_);
  and (_17598_, _17597_, _17586_);
  or (_17599_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_17600_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_17601_, _17600_, _10928_);
  and (_17602_, _17601_, _17599_);
  or (_17603_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_17604_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and (_17605_, _17604_, _04832_);
  and (_17606_, _17605_, _17603_);
  or (_17607_, _17606_, _17602_);
  or (_17608_, _17607_, _10926_);
  or (_17609_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_17610_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_17611_, _17610_, _10928_);
  and (_17612_, _17611_, _17609_);
  or (_17613_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_17614_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and (_17615_, _17614_, _04832_);
  and (_17616_, _17615_, _17613_);
  or (_17617_, _17616_, _17612_);
  or (_17618_, _17617_, _04868_);
  and (_17619_, _17618_, _04859_);
  and (_17620_, _17619_, _17608_);
  or (_17621_, _17620_, _17598_);
  and (_17622_, _17621_, _10997_);
  and (_17623_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_17624_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_17625_, _17624_, _17623_);
  and (_17626_, _17625_, _04832_);
  and (_17627_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_17628_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_17629_, _17628_, _17627_);
  and (_17630_, _17629_, _10928_);
  or (_17631_, _17630_, _17626_);
  or (_17632_, _17631_, _10926_);
  and (_17633_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_17635_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_17636_, _17635_, _17633_);
  and (_17637_, _17636_, _04832_);
  and (_17638_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_17639_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_17640_, _17639_, _17638_);
  and (_17641_, _17640_, _10928_);
  or (_17642_, _17641_, _17637_);
  or (_17643_, _17642_, _04868_);
  and (_17644_, _17643_, _10945_);
  and (_17645_, _17644_, _17632_);
  or (_17646_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_17647_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_17648_, _17647_, _17646_);
  and (_17649_, _17648_, _04832_);
  or (_17650_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_17651_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_17652_, _17651_, _17650_);
  and (_17653_, _17652_, _10928_);
  or (_17654_, _17653_, _17649_);
  or (_17656_, _17654_, _10926_);
  or (_17657_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_17658_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_17659_, _17658_, _17657_);
  and (_17660_, _17659_, _04832_);
  or (_17661_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_17662_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_17663_, _17662_, _17661_);
  and (_17664_, _17663_, _10928_);
  or (_17665_, _17664_, _17660_);
  or (_17666_, _17665_, _04868_);
  and (_17667_, _17666_, _04859_);
  and (_17668_, _17667_, _17656_);
  or (_17669_, _17668_, _17645_);
  and (_17670_, _17669_, _04849_);
  or (_17671_, _17670_, _17622_);
  and (_17672_, _17671_, _10996_);
  or (_17673_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_17674_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_17675_, _17674_, _17673_);
  and (_17676_, _17675_, _04832_);
  or (_17677_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_17678_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and (_17679_, _17678_, _17677_);
  and (_17680_, _17679_, _10928_);
  or (_17681_, _17680_, _17676_);
  and (_17682_, _17681_, _10926_);
  or (_17683_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_17684_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_17685_, _17684_, _17683_);
  and (_17686_, _17685_, _04832_);
  or (_17687_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_17688_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_17689_, _17688_, _17687_);
  and (_17690_, _17689_, _10928_);
  or (_17691_, _17690_, _17686_);
  and (_17692_, _17691_, _04868_);
  or (_17693_, _17692_, _17682_);
  and (_17694_, _17693_, _04859_);
  and (_17695_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_17696_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_17697_, _17696_, _17695_);
  and (_17698_, _17697_, _04832_);
  and (_17699_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_17700_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_17701_, _17700_, _17699_);
  and (_17702_, _17701_, _10928_);
  or (_17703_, _17702_, _17698_);
  and (_17704_, _17703_, _10926_);
  and (_17705_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and (_17706_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_17707_, _17706_, _17705_);
  and (_17708_, _17707_, _04832_);
  and (_17709_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and (_17710_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_17711_, _17710_, _17709_);
  and (_17712_, _17711_, _10928_);
  or (_17713_, _17712_, _17708_);
  and (_17714_, _17713_, _04868_);
  or (_17715_, _17714_, _17704_);
  and (_17716_, _17715_, _10945_);
  or (_17717_, _17716_, _17694_);
  and (_17718_, _17717_, _04849_);
  or (_17719_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_17720_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_17721_, _17720_, _10928_);
  and (_17722_, _17721_, _17719_);
  or (_17723_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_17724_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_17725_, _17724_, _04832_);
  and (_17726_, _17725_, _17723_);
  or (_17727_, _17726_, _17722_);
  and (_17728_, _17727_, _10926_);
  or (_17729_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_17730_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and (_17731_, _17730_, _10928_);
  and (_17732_, _17731_, _17729_);
  or (_17733_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_17734_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_17735_, _17734_, _04832_);
  and (_17736_, _17735_, _17733_);
  or (_17737_, _17736_, _17732_);
  and (_17738_, _17737_, _04868_);
  or (_17739_, _17738_, _17728_);
  and (_17740_, _17739_, _04859_);
  and (_17741_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and (_17742_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_17743_, _17742_, _17741_);
  and (_17744_, _17743_, _04832_);
  and (_17745_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_17746_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_17747_, _17746_, _17745_);
  and (_17748_, _17747_, _10928_);
  or (_17749_, _17748_, _17744_);
  and (_17750_, _17749_, _10926_);
  and (_17751_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_17752_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_17753_, _17752_, _17751_);
  and (_17754_, _17753_, _04832_);
  and (_17755_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_17756_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_17757_, _17756_, _17755_);
  and (_17758_, _17757_, _10928_);
  or (_17759_, _17758_, _17754_);
  and (_17760_, _17759_, _04868_);
  or (_17761_, _17760_, _17750_);
  and (_17762_, _17761_, _10945_);
  or (_17763_, _17762_, _17740_);
  and (_17764_, _17763_, _10997_);
  or (_17765_, _17764_, _17718_);
  and (_17766_, _17765_, _04839_);
  or (_17767_, _17766_, _17672_);
  or (_17768_, _17767_, _11204_);
  and (_17769_, _17768_, _17575_);
  or (_17770_, _17769_, _26153_);
  and (_17771_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_17772_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_17773_, _17772_, _17771_);
  and (_17774_, _17773_, _10928_);
  and (_17775_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_17776_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_17777_, _17776_, _17775_);
  and (_17778_, _17777_, _04832_);
  or (_17779_, _17778_, _17774_);
  or (_17780_, _17779_, _10926_);
  and (_17781_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_17782_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_17783_, _17782_, _17781_);
  and (_17784_, _17783_, _10928_);
  and (_17785_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_17786_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_17787_, _17786_, _17785_);
  and (_17788_, _17787_, _04832_);
  or (_17789_, _17788_, _17784_);
  or (_17790_, _17789_, _04868_);
  and (_17791_, _17790_, _10945_);
  and (_17792_, _17791_, _17780_);
  or (_17793_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_17794_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_17795_, _17794_, _04832_);
  and (_17796_, _17795_, _17793_);
  or (_17797_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_17798_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_17799_, _17798_, _10928_);
  and (_17800_, _17799_, _17797_);
  or (_17801_, _17800_, _17796_);
  or (_17802_, _17801_, _10926_);
  or (_17803_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_17804_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_17805_, _17804_, _04832_);
  and (_17806_, _17805_, _17803_);
  or (_17807_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_17808_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_17809_, _17808_, _10928_);
  and (_17810_, _17809_, _17807_);
  or (_17811_, _17810_, _17806_);
  or (_17812_, _17811_, _04868_);
  and (_17813_, _17812_, _04859_);
  and (_17814_, _17813_, _17802_);
  or (_17815_, _17814_, _17792_);
  and (_17816_, _17815_, _10997_);
  and (_17817_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_17818_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_17819_, _17818_, _04832_);
  or (_17820_, _17819_, _17817_);
  and (_17821_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_17822_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_17823_, _17822_, _10928_);
  or (_17824_, _17823_, _17821_);
  and (_17825_, _17824_, _17820_);
  or (_17826_, _17825_, _10926_);
  and (_17827_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_17828_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_17829_, _17828_, _04832_);
  or (_17830_, _17829_, _17827_);
  and (_17831_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_17832_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_17833_, _17832_, _10928_);
  or (_17834_, _17833_, _17831_);
  and (_17835_, _17834_, _17830_);
  or (_17836_, _17835_, _04868_);
  and (_17837_, _17836_, _10945_);
  and (_17838_, _17837_, _17826_);
  or (_17839_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_17840_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_17841_, _17840_, _17839_);
  or (_17842_, _17841_, _10928_);
  or (_17843_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_17844_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_17845_, _17844_, _17843_);
  or (_17846_, _17845_, _04832_);
  and (_17847_, _17846_, _17842_);
  or (_17848_, _17847_, _10926_);
  or (_17849_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_17850_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_17851_, _17850_, _17849_);
  or (_17852_, _17851_, _10928_);
  or (_17853_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_17854_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_17855_, _17854_, _17853_);
  or (_17856_, _17855_, _04832_);
  and (_17857_, _17856_, _17852_);
  or (_17858_, _17857_, _04868_);
  and (_17859_, _17858_, _04859_);
  and (_17860_, _17859_, _17848_);
  or (_17861_, _17860_, _17838_);
  and (_17862_, _17861_, _04849_);
  or (_17863_, _17862_, _17816_);
  and (_17864_, _17863_, _10996_);
  and (_17865_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  and (_17866_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or (_17867_, _17866_, _17865_);
  and (_17868_, _17867_, _04832_);
  and (_17869_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  and (_17870_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or (_17871_, _17870_, _17869_);
  and (_17872_, _17871_, _10928_);
  or (_17873_, _17872_, _17868_);
  and (_17874_, _17873_, _04868_);
  and (_17875_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and (_17876_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or (_17877_, _17876_, _17875_);
  and (_17878_, _17877_, _04832_);
  and (_17879_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and (_17880_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or (_17881_, _17880_, _17879_);
  and (_17882_, _17881_, _10928_);
  or (_17883_, _17882_, _17878_);
  and (_17884_, _17883_, _10926_);
  or (_17885_, _17884_, _17874_);
  and (_17886_, _17885_, _10945_);
  or (_17887_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or (_17888_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and (_17889_, _17888_, _17887_);
  and (_17890_, _17889_, _04832_);
  or (_17891_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or (_17892_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and (_17893_, _17892_, _17891_);
  and (_17894_, _17893_, _10928_);
  or (_17895_, _17894_, _17890_);
  and (_17896_, _17895_, _04868_);
  or (_17897_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or (_17898_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and (_17899_, _17898_, _17897_);
  and (_17900_, _17899_, _04832_);
  or (_17901_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or (_17902_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and (_17903_, _17902_, _17901_);
  and (_17904_, _17903_, _10928_);
  or (_17905_, _17904_, _17900_);
  and (_17906_, _17905_, _10926_);
  or (_17907_, _17906_, _17896_);
  and (_17908_, _17907_, _04859_);
  or (_17909_, _17908_, _17886_);
  and (_17910_, _17909_, _10997_);
  and (_17911_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_17912_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_17913_, _17912_, _17911_);
  and (_17914_, _17913_, _04832_);
  and (_17915_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_17916_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_17917_, _17916_, _17915_);
  and (_17918_, _17917_, _10928_);
  or (_17919_, _17918_, _17914_);
  and (_17920_, _17919_, _04868_);
  and (_17921_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_17922_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_17923_, _17922_, _17921_);
  and (_17924_, _17923_, _04832_);
  and (_17925_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_17926_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_17927_, _17926_, _17925_);
  and (_17928_, _17927_, _10928_);
  or (_17929_, _17928_, _17924_);
  and (_17930_, _17929_, _10926_);
  or (_17931_, _17930_, _17920_);
  and (_17932_, _17931_, _10945_);
  or (_17933_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_17934_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_17935_, _17934_, _17933_);
  and (_17936_, _17935_, _04832_);
  or (_17937_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_17938_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_17939_, _17938_, _17937_);
  and (_17940_, _17939_, _10928_);
  or (_17941_, _17940_, _17936_);
  and (_17942_, _17941_, _04868_);
  or (_17943_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_17944_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_17945_, _17944_, _17943_);
  and (_17946_, _17945_, _04832_);
  or (_17947_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_17948_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_17949_, _17948_, _17947_);
  and (_17950_, _17949_, _10928_);
  or (_17951_, _17950_, _17946_);
  and (_17952_, _17951_, _10926_);
  or (_17953_, _17952_, _17942_);
  and (_17954_, _17953_, _04859_);
  or (_17955_, _17954_, _17932_);
  and (_17956_, _17955_, _04849_);
  or (_17957_, _17956_, _17910_);
  and (_17958_, _17957_, _04839_);
  or (_17959_, _17958_, _17864_);
  or (_17960_, _17959_, _04843_);
  and (_17961_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_17962_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_17963_, _17962_, _17961_);
  and (_17964_, _17963_, _04832_);
  and (_17965_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_17966_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_17967_, _17966_, _17965_);
  and (_17968_, _17967_, _10928_);
  or (_17969_, _17968_, _17964_);
  or (_17970_, _17969_, _10926_);
  and (_17971_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_17972_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_17973_, _17972_, _17971_);
  and (_17974_, _17973_, _04832_);
  and (_17975_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_17976_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_17977_, _17976_, _17975_);
  and (_17978_, _17977_, _10928_);
  or (_17979_, _17978_, _17974_);
  or (_17980_, _17979_, _04868_);
  and (_17981_, _17980_, _10945_);
  and (_17982_, _17981_, _17970_);
  or (_17983_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_17984_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_17985_, _17984_, _10928_);
  and (_17986_, _17985_, _17983_);
  or (_17987_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_17988_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_17989_, _17988_, _04832_);
  and (_17990_, _17989_, _17987_);
  or (_17991_, _17990_, _17986_);
  or (_17992_, _17991_, _10926_);
  or (_17993_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_17994_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_17995_, _17994_, _10928_);
  and (_17996_, _17995_, _17993_);
  or (_17997_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_17998_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_17999_, _17998_, _04832_);
  and (_18000_, _17999_, _17997_);
  or (_18001_, _18000_, _17996_);
  or (_18002_, _18001_, _04868_);
  and (_18003_, _18002_, _04859_);
  and (_18004_, _18003_, _17992_);
  or (_18005_, _18004_, _17982_);
  and (_18006_, _18005_, _10997_);
  and (_18007_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_18008_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_18009_, _18008_, _18007_);
  and (_18010_, _18009_, _04832_);
  and (_18011_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_18012_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_18013_, _18012_, _18011_);
  and (_18014_, _18013_, _10928_);
  or (_18015_, _18014_, _18010_);
  or (_18016_, _18015_, _10926_);
  and (_18017_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_18018_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_18019_, _18018_, _18017_);
  and (_18020_, _18019_, _04832_);
  and (_18021_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_18022_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_18023_, _18022_, _18021_);
  and (_18024_, _18023_, _10928_);
  or (_18025_, _18024_, _18020_);
  or (_18026_, _18025_, _04868_);
  and (_18027_, _18026_, _10945_);
  and (_18028_, _18027_, _18016_);
  or (_18029_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_18030_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_18031_, _18030_, _18029_);
  and (_18032_, _18031_, _04832_);
  or (_18033_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_18034_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_18035_, _18034_, _18033_);
  and (_18036_, _18035_, _10928_);
  or (_18037_, _18036_, _18032_);
  or (_18038_, _18037_, _10926_);
  or (_18039_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_18040_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_18041_, _18040_, _18039_);
  and (_18042_, _18041_, _04832_);
  or (_18043_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_18044_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_18045_, _18044_, _18043_);
  and (_18046_, _18045_, _10928_);
  or (_18047_, _18046_, _18042_);
  or (_18048_, _18047_, _04868_);
  and (_18049_, _18048_, _04859_);
  and (_18050_, _18049_, _18038_);
  or (_18051_, _18050_, _18028_);
  and (_18052_, _18051_, _04849_);
  or (_18053_, _18052_, _18006_);
  and (_18054_, _18053_, _10996_);
  or (_18055_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_18056_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_18057_, _18056_, _18055_);
  and (_18058_, _18057_, _04832_);
  or (_18059_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_18060_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_18061_, _18060_, _18059_);
  and (_18062_, _18061_, _10928_);
  or (_18063_, _18062_, _18058_);
  and (_18064_, _18063_, _10926_);
  or (_18065_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_18066_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_18067_, _18066_, _18065_);
  and (_18068_, _18067_, _04832_);
  or (_18069_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_18070_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_18071_, _18070_, _18069_);
  and (_18072_, _18071_, _10928_);
  or (_18073_, _18072_, _18068_);
  and (_18074_, _18073_, _04868_);
  or (_18075_, _18074_, _18064_);
  and (_18076_, _18075_, _04859_);
  and (_18077_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_18078_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_18079_, _18078_, _18077_);
  and (_18080_, _18079_, _04832_);
  and (_18081_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_18082_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_18083_, _18082_, _18081_);
  and (_18084_, _18083_, _10928_);
  or (_18085_, _18084_, _18080_);
  and (_18086_, _18085_, _10926_);
  and (_18087_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_18088_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_18089_, _18088_, _18087_);
  and (_18090_, _18089_, _04832_);
  and (_18091_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_18092_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_18093_, _18092_, _18091_);
  and (_18094_, _18093_, _10928_);
  or (_18095_, _18094_, _18090_);
  and (_18096_, _18095_, _04868_);
  or (_18097_, _18096_, _18086_);
  and (_18098_, _18097_, _10945_);
  or (_18099_, _18098_, _18076_);
  and (_18100_, _18099_, _04849_);
  or (_18101_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_18102_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and (_18103_, _18102_, _10928_);
  and (_18104_, _18103_, _18101_);
  or (_18105_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_18106_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_18107_, _18106_, _04832_);
  and (_18108_, _18107_, _18105_);
  or (_18109_, _18108_, _18104_);
  and (_18110_, _18109_, _10926_);
  or (_18111_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_18112_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_18113_, _18112_, _10928_);
  and (_18114_, _18113_, _18111_);
  or (_18115_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_18116_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and (_18117_, _18116_, _04832_);
  and (_18118_, _18117_, _18115_);
  or (_18119_, _18118_, _18114_);
  and (_18120_, _18119_, _04868_);
  or (_18121_, _18120_, _18110_);
  and (_18122_, _18121_, _04859_);
  and (_18123_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_18124_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_18125_, _18124_, _18123_);
  and (_18126_, _18125_, _04832_);
  and (_18127_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_18128_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_18129_, _18128_, _18127_);
  and (_18130_, _18129_, _10928_);
  or (_18131_, _18130_, _18126_);
  and (_18132_, _18131_, _10926_);
  and (_18133_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_18134_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_18135_, _18134_, _18133_);
  and (_18136_, _18135_, _04832_);
  and (_18137_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_18138_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_18139_, _18138_, _18137_);
  and (_18140_, _18139_, _10928_);
  or (_18141_, _18140_, _18136_);
  and (_18142_, _18141_, _04868_);
  or (_18143_, _18142_, _18132_);
  and (_18144_, _18143_, _10945_);
  or (_18145_, _18144_, _18122_);
  and (_18146_, _18145_, _10997_);
  or (_18147_, _18146_, _18100_);
  and (_18148_, _18147_, _04839_);
  or (_18149_, _18148_, _18054_);
  or (_18150_, _18149_, _11204_);
  and (_18151_, _18150_, _17960_);
  or (_18152_, _18151_, _03196_);
  and (_18153_, _18152_, _17770_);
  or (_18154_, _18153_, _04876_);
  or (_18155_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_18156_, _18155_, _22773_);
  and (_08982_, _18156_, _18154_);
  and (_18157_, _23924_, _23453_);
  and (_18158_, _18157_, _24027_);
  not (_18159_, _18157_);
  and (_18160_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or (_08989_, _18160_, _18158_);
  and (_18161_, _18157_, _23920_);
  and (_18162_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_08991_, _18162_, _18161_);
  and (_18163_, _24130_, _23700_);
  and (_18164_, _18163_, _23751_);
  not (_18165_, _18163_);
  and (_18166_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or (_27311_, _18166_, _18164_);
  and (_18167_, _24130_, _23938_);
  and (_18168_, _18167_, _24027_);
  not (_18169_, _18167_);
  and (_18170_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_09010_, _18170_, _18168_);
  and (_18171_, _18167_, _23693_);
  and (_18172_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_09013_, _18172_, _18171_);
  and (_18173_, _02853_, _23900_);
  and (_18174_, _02856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or (_09015_, _18174_, _18173_);
  and (_18175_, _24124_, _23924_);
  and (_18176_, _18175_, _24027_);
  not (_18177_, _18175_);
  and (_18178_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_09019_, _18178_, _18176_);
  and (_18179_, _18175_, _23715_);
  and (_18180_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_09022_, _18180_, _18179_);
  and (_18181_, _18175_, _24053_);
  and (_18182_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_09025_, _18182_, _18181_);
  or (_18183_, _16264_, _24027_);
  or (_18184_, _16263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and (_09029_, _18184_, _18183_);
  and (_18185_, _24145_, _24124_);
  and (_18186_, _18185_, _23983_);
  not (_18187_, _18185_);
  and (_18188_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_09032_, _18188_, _18186_);
  and (_18189_, _18185_, _23920_);
  and (_18190_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or (_09034_, _18190_, _18189_);
  and (_18191_, _18185_, _23751_);
  and (_18192_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or (_27308_, _18192_, _18191_);
  and (_18193_, _18157_, _23900_);
  and (_18194_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or (_09045_, _18194_, _18193_);
  and (_18195_, _24274_, _24124_);
  and (_18196_, _18195_, _24027_);
  not (_18197_, _18195_);
  and (_18198_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or (_27307_, _18198_, _18196_);
  and (_18199_, _17246_, _23715_);
  and (_18200_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or (_09073_, _18200_, _18199_);
  and (_18201_, _17246_, _23900_);
  and (_18202_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or (_09083_, _18202_, _18201_);
  and (_18203_, _17246_, _23920_);
  and (_18204_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or (_09085_, _18204_, _18203_);
  and (_18205_, _02248_, _24053_);
  and (_18206_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or (_09092_, _18206_, _18205_);
  and (_18207_, _18195_, _23693_);
  and (_18208_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or (_09104_, _18208_, _18207_);
  and (_18209_, _24124_, _23905_);
  and (_18210_, _18209_, _23983_);
  not (_18211_, _18209_);
  and (_18212_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_09108_, _18212_, _18210_);
  and (_18213_, _18209_, _23715_);
  and (_18214_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_09110_, _18214_, _18213_);
  and (_18215_, _24124_, _23930_);
  and (_18216_, _18215_, _23751_);
  not (_18217_, _18215_);
  and (_18218_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or (_09114_, _18218_, _18216_);
  and (_18219_, _24124_, _24061_);
  and (_18220_, _18219_, _23900_);
  not (_18221_, _18219_);
  and (_18222_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or (_09118_, _18222_, _18220_);
  and (_18223_, _18219_, _23751_);
  and (_18224_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or (_27299_, _18224_, _18223_);
  and (_18225_, _23920_, _23721_);
  and (_18226_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_09128_, _18226_, _18225_);
  and (_18227_, _24124_, _24108_);
  and (_18228_, _18227_, _23920_);
  not (_18229_, _18227_);
  and (_18230_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_27297_, _18230_, _18228_);
  and (_18231_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and (_18232_, _16270_, _23750_);
  or (_09131_, _18232_, _18231_);
  and (_18233_, _10273_, _24053_);
  and (_18234_, _10275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or (_09134_, _18234_, _18233_);
  and (_18235_, _09480_, _23751_);
  and (_18236_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or (_09137_, _18236_, _18235_);
  and (_18237_, _09480_, _24053_);
  and (_18238_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or (_09142_, _18238_, _18237_);
  and (_18239_, _18227_, _23715_);
  and (_18240_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_09147_, _18240_, _18239_);
  and (_18241_, _18227_, _24053_);
  and (_18242_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_09149_, _18242_, _18241_);
  and (_18243_, _24219_, _24027_);
  and (_18244_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or (_09151_, _18244_, _18243_);
  and (_18245_, _24124_, _23444_);
  and (_18246_, _18245_, _23693_);
  not (_18247_, _18245_);
  and (_18248_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_09155_, _18248_, _18246_);
  and (_18249_, _18245_, _24053_);
  and (_18250_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_09157_, _18250_, _18249_);
  and (_18251_, _18215_, _23983_);
  and (_18252_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or (_27306_, _18252_, _18251_);
  and (_18253_, _18215_, _23920_);
  and (_18254_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or (_09162_, _18254_, _18253_);
  and (_18255_, _24231_, _23751_);
  and (_18256_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or (_27314_, _18256_, _18255_);
  and (_18257_, _18163_, _24027_);
  and (_18258_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or (_09165_, _18258_, _18257_);
  and (_18259_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  and (_18260_, _02838_, _24027_);
  or (_09167_, _18260_, _18259_);
  and (_18261_, _16271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_18262_, _16270_, _23692_);
  or (_09169_, _18262_, _18261_);
  and (_18263_, _18163_, _23715_);
  and (_18264_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or (_09171_, _18264_, _18263_);
  and (_18265_, _18167_, _23900_);
  and (_18266_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_09173_, _18266_, _18265_);
  and (_18267_, _25165_, _24027_);
  and (_18268_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_09187_, _18268_, _18267_);
  and (_18269_, _01932_, _23900_);
  and (_18270_, _01934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_09190_, _18270_, _18269_);
  and (_18271_, _02509_, _24027_);
  and (_18272_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_09200_, _18272_, _18271_);
  and (_18273_, _24069_, _23983_);
  and (_18274_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or (_27196_, _18274_, _18273_);
  and (_18275_, _02350_, _23751_);
  and (_18276_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_09208_, _18276_, _18275_);
  and (_18278_, _18209_, _24053_);
  and (_18279_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_09231_, _18279_, _18278_);
  and (_18280_, _17017_, _23983_);
  and (_18281_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_09235_, _18281_, _18280_);
  and (_18282_, _18227_, _23983_);
  and (_18283_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_09241_, _18283_, _18282_);
  and (_18284_, _25176_, _23715_);
  and (_18285_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or (_09245_, _18285_, _18284_);
  and (_18286_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  and (_18287_, _02838_, _23920_);
  or (_09249_, _18287_, _18286_);
  and (_18288_, _18245_, _23900_);
  and (_18289_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_09251_, _18289_, _18288_);
  and (_18290_, _18175_, _23751_);
  and (_18291_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_09265_, _18291_, _18290_);
  and (_18292_, _18157_, _24053_);
  and (_18293_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or (_09268_, _18293_, _18292_);
  and (_18294_, _09485_, _24027_);
  and (_18295_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_09275_, _18295_, _18294_);
  and (_18296_, _10411_, _24053_);
  and (_18297_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or (_27038_, _18297_, _18296_);
  and (_18298_, _18185_, _23693_);
  and (_18299_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or (_09280_, _18299_, _18298_);
  and (_18300_, _18209_, _23900_);
  and (_18301_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_09283_, _18301_, _18300_);
  and (_18302_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  and (_18303_, _02838_, _23751_);
  or (_09291_, _18303_, _18302_);
  and (_18304_, _18195_, _23715_);
  and (_18305_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or (_09293_, _18305_, _18304_);
  and (_18306_, _18245_, _23920_);
  and (_18307_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_09296_, _18307_, _18306_);
  and (_18308_, _18215_, _23900_);
  and (_18309_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or (_09305_, _18309_, _18308_);
  and (_18310_, _17216_, _23900_);
  and (_18311_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_09307_, _18311_, _18310_);
  and (_18312_, _18215_, _23693_);
  and (_18313_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or (_09309_, _18313_, _18312_);
  and (_18314_, _23751_, _23707_);
  and (_18315_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_09311_, _18315_, _18314_);
  and (_18316_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  and (_18317_, _02838_, _24053_);
  or (_09313_, _18317_, _18316_);
  and (_18318_, _17216_, _23751_);
  and (_18319_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_27281_, _18319_, _18318_);
  and (_18320_, _16264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  and (_18321_, _16268_, _24052_);
  or (_09317_, _18321_, _18320_);
  and (_18322_, _16264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and (_18323_, _16268_, _23692_);
  or (_09319_, _18323_, _18322_);
  and (_18324_, _16264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and (_18325_, _16268_, _23750_);
  or (_09321_, _18325_, _18324_);
  and (_18326_, _18215_, _23715_);
  and (_18327_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or (_09326_, _18327_, _18326_);
  and (_18328_, _09485_, _23983_);
  and (_18329_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_09363_, _18329_, _18328_);
  and (_18330_, _18157_, _23715_);
  and (_18331_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or (_09369_, _18331_, _18330_);
  or (_18332_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_18333_, _18332_, _22773_);
  or (_18334_, _23744_, _22931_);
  and (_09373_, _18334_, _18333_);
  and (_18335_, _18157_, _23693_);
  and (_18336_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or (_09380_, _18336_, _18335_);
  and (_18337_, _02839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  and (_18338_, _02838_, _23693_);
  or (_09387_, _18338_, _18337_);
  and (_18339_, _10411_, _23751_);
  and (_18340_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or (_27039_, _18340_, _18339_);
  and (_18341_, _10411_, _23715_);
  and (_18342_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or (_09447_, _18342_, _18341_);
  and (_18343_, _17017_, _23715_);
  and (_18344_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_27216_, _18344_, _18343_);
  and (_18345_, _10411_, _23693_);
  and (_18346_, _10413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or (_09464_, _18346_, _18345_);
  and (_18347_, _17017_, _23693_);
  and (_18348_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_09473_, _18348_, _18347_);
  and (_18349_, _15255_, _23920_);
  and (_18350_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or (_09474_, _18350_, _18349_);
  nand (_18351_, _24047_, _22922_);
  or (_18352_, _22922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_18353_, _18352_, _22773_);
  and (_09477_, _18353_, _18351_);
  and (_18354_, _09507_, _23751_);
  and (_18355_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_09484_, _18355_, _18354_);
  and (_18356_, _01927_, _23920_);
  and (_18357_, _01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_09521_, _18357_, _18356_);
  and (_18358_, _17069_, _23751_);
  and (_18359_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_09539_, _18359_, _18358_);
  and (_18360_, _17069_, _24053_);
  and (_18361_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_27254_, _18361_, _18360_);
  and (_18362_, _09485_, _23751_);
  and (_18363_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_09571_, _18363_, _18362_);
  and (_18364_, _01709_, _24027_);
  and (_18365_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_09591_, _18365_, _18364_);
  and (_18366_, _17017_, _23920_);
  and (_18367_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_09594_, _18367_, _18366_);
  and (_18368_, _09485_, _24053_);
  and (_18369_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_09607_, _18369_, _18368_);
  and (_18370_, _01709_, _23920_);
  and (_18371_, _01712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_09623_, _18371_, _18370_);
  and (_18372_, _17017_, _23900_);
  and (_18373_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_09633_, _18373_, _18372_);
  and (_18374_, _09507_, _24053_);
  and (_18375_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_09646_, _18375_, _18374_);
  and (_18376_, _02326_, _23751_);
  and (_18377_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_09659_, _18377_, _18376_);
  and (_18378_, _09463_, _23983_);
  and (_18379_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_27056_, _18379_, _18378_);
  and (_18380_, _17083_, _23715_);
  and (_18381_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or (_09675_, _18381_, _18380_);
  and (_18382_, _17083_, _23693_);
  and (_18383_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or (_09689_, _18383_, _18382_);
  and (_18384_, _17083_, _23751_);
  and (_18385_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or (_09708_, _18385_, _18384_);
  and (_18386_, _02829_, _24027_);
  and (_18387_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or (_09777_, _18387_, _18386_);
  and (_18388_, _17216_, _23715_);
  and (_18389_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_09781_, _18389_, _18388_);
  nand (_09789_, _26302_, _22773_);
  and (_26864_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _22773_);
  and (_18390_, _24062_, _23920_);
  and (_18391_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_09812_, _18391_, _18390_);
  nor (_09819_, _25982_, rst);
  and (_18392_, _24027_, _23721_);
  and (_18393_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_09828_, _18393_, _18392_);
  and (_18394_, _18215_, _24027_);
  and (_18395_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or (_27305_, _18395_, _18394_);
  and (_18396_, _17216_, _24027_);
  and (_18397_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_27282_, _18397_, _18396_);
  and (_18398_, _02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_18399_, _02775_, _24053_);
  or (_09834_, _18399_, _18398_);
  nor (_09841_, _26035_, rst);
  or (_18400_, _01045_, _01043_);
  or (_18401_, _01046_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_18402_, _18401_, _18400_);
  nand (_18403_, _18402_, _03274_);
  or (_18404_, _18402_, _03274_);
  and (_18405_, _18404_, _18403_);
  and (_18406_, _18405_, _00040_);
  and (_18407_, _26801_, _26149_);
  and (_18408_, _00619_, _24643_);
  and (_18409_, _03293_, _26799_);
  nor (_18410_, _01091_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_18411_, _01091_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_18412_, _18411_, _18410_);
  and (_18413_, _18412_, _00045_);
  and (_18414_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_18415_, _18414_, _18413_);
  or (_18416_, _18415_, _18409_);
  or (_18417_, _18416_, _18408_);
  nor (_18418_, _18417_, _18407_);
  nand (_18419_, _18418_, _26378_);
  or (_18420_, _18419_, _18406_);
  not (_18421_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_18422_, _01110_, _18421_);
  and (_18423_, _01110_, _18421_);
  or (_18424_, _18423_, _18422_);
  or (_18425_, _18424_, _26378_);
  and (_18426_, _18425_, _22773_);
  and (_26861_[15], _18426_, _18420_);
  and (_18427_, _17216_, _23983_);
  and (_18428_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_09846_, _18428_, _18427_);
  and (_18429_, _24053_, _23454_);
  and (_18430_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or (_09848_, _18430_, _18429_);
  nor (_26856_[4], _25661_, rst);
  and (_18431_, _23920_, _23454_);
  and (_18432_, _23695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_09859_, _18432_, _18431_);
  nor (_09862_, _26091_, rst);
  and (_18433_, _18245_, _23751_);
  and (_18434_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_09864_, _18434_, _18433_);
  and (_18435_, _17184_, _24053_);
  and (_18436_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_09874_, _18436_, _18435_);
  or (_18437_, _24664_, _01894_);
  or (_18438_, _23759_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_18439_, _18438_, _22773_);
  and (_26835_[4], _18439_, _18437_);
  and (_18440_, _18245_, _23715_);
  and (_18441_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_09883_, _18441_, _18440_);
  and (_18442_, _17184_, _23693_);
  and (_18443_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_09885_, _18443_, _18442_);
  and (_18444_, _01952_, _24053_);
  and (_18445_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or (_09895_, _18445_, _18444_);
  nor (_18446_, _01504_, rst);
  nand (_18447_, _23760_, _01368_);
  and (_18448_, _18447_, _26864_);
  or (_26865_, _18448_, _18446_);
  and (_18449_, _24219_, _23900_);
  and (_18450_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or (_09902_, _18450_, _18449_);
  nor (_18451_, _01487_, _01477_);
  nor (_18452_, _18451_, _01486_);
  or (_18453_, _18452_, _18412_);
  nand (_18454_, _18452_, _18412_);
  and (_18455_, _18454_, _24816_);
  and (_18456_, _18455_, _18453_);
  nor (_18457_, _24816_, _03274_);
  or (_18458_, _18457_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_18459_, _18458_, _18456_);
  or (_18460_, _01368_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_18461_, _18460_, _22773_);
  and (_26862_[15], _18461_, _18459_);
  and (_18462_, _24215_, _23693_);
  and (_18463_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_09909_, _18463_, _18462_);
  and (_18464_, _16264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and (_18465_, _16268_, _23899_);
  or (_09911_, _18465_, _18464_);
  nand (_09915_, _26324_, _22773_);
  and (_18466_, _16720_, _23693_);
  and (_18467_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_09917_, _18467_, _18466_);
  and (_18468_, _24342_, _22857_);
  nand (_18469_, _18468_, _23250_);
  and (_18470_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_18471_, _25234_, _23249_);
  and (_18472_, _18471_, _22857_);
  and (_18473_, _18472_, _22914_);
  and (_18474_, _18473_, _22910_);
  and (_18475_, _18474_, _00619_);
  or (_18476_, _18475_, _18470_);
  or (_18477_, _18476_, _03856_);
  not (_18478_, _03856_);
  or (_18479_, _18478_, _03293_);
  and (_18480_, _18479_, _22773_);
  and (_09919_, _18480_, _18477_);
  and (_18481_, _16682_, _23983_);
  and (_18482_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_09920_, _18482_, _18481_);
  and (_18483_, _24027_, _23939_);
  and (_18484_, _23941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or (_09923_, _18484_, _18483_);
  and (_18485_, _01504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_18486_, _18485_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_26866_[7], _18486_, _22773_);
  and (_18487_, _18468_, _24184_);
  nor (_18488_, _18487_, _03856_);
  or (_18489_, _18488_, _00619_);
  not (_18490_, _18488_);
  or (_18491_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_18492_, _18491_, _22773_);
  and (_09928_, _18492_, _18489_);
  and (_18493_, _25190_, _23693_);
  and (_18494_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_09933_, _18494_, _18493_);
  and (_18495_, _24219_, _23920_);
  and (_18496_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_09935_, _18496_, _18495_);
  and (_18498_, _24215_, _23715_);
  and (_18499_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or (_09938_, _18499_, _18498_);
  and (_18500_, _24219_, _23983_);
  and (_18501_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or (_09940_, _18501_, _18500_);
  and (_18502_, _24215_, _23920_);
  and (_18503_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or (_09943_, _18503_, _18502_);
  nor (_18504_, _25524_, _24883_);
  nor (_18505_, _01532_, _01529_);
  nor (_18506_, _18505_, _24883_);
  and (_18507_, _18506_, _24468_);
  nor (_18508_, _18506_, _24468_);
  nor (_18509_, _18508_, _18507_);
  nor (_18510_, _18509_, _18504_);
  and (_18511_, _24473_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_18512_, _18511_, _18504_);
  nor (_18513_, _18512_, _01286_);
  or (_18514_, _18513_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_18515_, _18514_, _18510_);
  and (_26867_[2], _18515_, _22773_);
  and (_26857_[7], _26147_, _22773_);
  and (_18516_, _16264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  and (_18517_, _16268_, _23714_);
  or (_09951_, _18517_, _18516_);
  and (_18518_, _25190_, _23920_);
  and (_18519_, _25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_09955_, _18519_, _18518_);
  nor (_09958_, _26053_, rst);
  and (_18520_, _25159_, _23715_);
  and (_18521_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or (_09962_, _18521_, _18520_);
  and (_18522_, _24215_, _24027_);
  and (_18523_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or (_09964_, _18523_, _18522_);
  and (_18524_, _25159_, _23751_);
  and (_18525_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or (_09966_, _18525_, _18524_);
  nor (_18526_, _24643_, rst);
  and (_26859_, _18526_, _26378_);
  and (_18527_, _18227_, _23751_);
  and (_18528_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_09970_, _18528_, _18527_);
  nand (_09974_, _26358_, _22773_);
  and (_26863_, _15274_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_18529_, _24069_, _23751_);
  and (_18530_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or (_09979_, _18530_, _18529_);
  and (_26860_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _22773_);
  and (_26855_, _26153_, _22773_);
  or (_18531_, _18488_, _26798_);
  or (_18532_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_18533_, _18532_, _22773_);
  and (_09993_, _18533_, _18531_);
  and (_18534_, _25159_, _23983_);
  and (_18535_, _25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or (_10011_, _18535_, _18534_);
  and (_18536_, _02779_, _23900_);
  and (_18537_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_10014_, _18537_, _18536_);
  and (_18538_, _24069_, _23920_);
  and (_18539_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or (_10016_, _18539_, _18538_);
  and (_18540_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_18541_, _18474_, _00101_);
  or (_18542_, _18541_, _18540_);
  or (_18543_, _18542_, _03856_);
  nand (_18544_, _03856_, _00747_);
  and (_18545_, _18544_, _22773_);
  and (_10021_, _18545_, _18543_);
  or (_18546_, _18488_, _00277_);
  or (_18547_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_18548_, _18547_, _22773_);
  and (_10023_, _18548_, _18546_);
  and (_18549_, _18227_, _23693_);
  and (_18550_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_10027_, _18550_, _18549_);
  and (_18551_, _17196_, _24053_);
  and (_18552_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_10029_, _18552_, _18551_);
  and (_18553_, _18227_, _23900_);
  and (_18554_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_10034_, _18554_, _18553_);
  and (_18555_, _02779_, _23715_);
  and (_18556_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_10037_, _18556_, _18555_);
  and (_18557_, _17196_, _23693_);
  and (_18558_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or (_10039_, _18558_, _18557_);
  and (_18559_, _18227_, _24027_);
  and (_18560_, _18229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_10041_, _18560_, _18559_);
  and (_18561_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_18562_, _18474_, _00352_);
  or (_18563_, _18562_, _18561_);
  or (_18564_, _18563_, _03856_);
  or (_18565_, _18478_, _00958_);
  and (_18566_, _18565_, _22773_);
  and (_10048_, _18566_, _18564_);
  and (_18567_, _17196_, _23900_);
  and (_18568_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or (_10050_, _18568_, _18567_);
  and (_18569_, _24319_, _23715_);
  and (_18570_, _24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_10056_, _18570_, _18569_);
  and (_18571_, _15225_, _24027_);
  and (_18572_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_26932_, _18572_, _18571_);
  and (_18573_, _18219_, _24053_);
  and (_18574_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or (_27298_, _18574_, _18573_);
  and (_18575_, _17196_, _24027_);
  and (_18576_, _17198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or (_10063_, _18576_, _18575_);
  and (_18577_, _25428_, _24053_);
  and (_18578_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_10066_, _18578_, _18577_);
  and (_18579_, _18219_, _23693_);
  and (_18580_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or (_10068_, _18580_, _18579_);
  and (_18581_, _25428_, _24027_);
  and (_18582_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_10072_, _18582_, _18581_);
  and (_18583_, _25428_, _23900_);
  and (_18584_, _25430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_10073_, _18584_, _18583_);
  and (_18585_, _17190_, _23751_);
  and (_18586_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_10076_, _18586_, _18585_);
  and (_18587_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_18588_, _18474_, _00277_);
  or (_18589_, _18588_, _18587_);
  or (_18590_, _18589_, _03856_);
  nand (_18591_, _03856_, _00878_);
  and (_18592_, _18591_, _22773_);
  and (_10082_, _18592_, _18590_);
  or (_26833_[2], _04969_, _01888_);
  and (_18593_, _17246_, _23693_);
  and (_18594_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or (_10087_, _18594_, _18593_);
  and (_18595_, _18219_, _23715_);
  and (_18596_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or (_27300_, _18596_, _18595_);
  or (_18597_, _18488_, _00564_);
  or (_18598_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_18599_, _18598_, _22773_);
  and (_10089_, _18599_, _18597_);
  and (_18600_, _15225_, _23920_);
  and (_18601_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_10091_, _18601_, _18600_);
  and (_18602_, _18219_, _23920_);
  and (_18603_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or (_10093_, _18603_, _18602_);
  and (_18604_, _17190_, _23693_);
  and (_18605_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_10095_, _18605_, _18604_);
  and (_18606_, _17246_, _24027_);
  and (_18607_, _17248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or (_10097_, _18607_, _18606_);
  and (_18608_, _18219_, _24027_);
  and (_18609_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or (_10098_, _18609_, _18608_);
  and (_18610_, _02423_, _23983_);
  and (_18611_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or (_10100_, _18611_, _18610_);
  nor (_26832_[2], _25866_, rst);
  and (_18612_, _17190_, _23900_);
  and (_18613_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_27280_, _18613_, _18612_);
  and (_18614_, _18219_, _23983_);
  and (_18615_, _18221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or (_10104_, _18615_, _18614_);
  and (_18616_, _17190_, _24027_);
  and (_18617_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_10105_, _18617_, _18616_);
  and (_18618_, _04207_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_18619_, _25877_);
  nand (_18620_, _00003_, _18619_);
  or (_18621_, _18620_, _06594_);
  or (_18622_, _04228_, _25898_);
  or (_18623_, _18622_, _26811_);
  or (_18624_, _18623_, _04227_);
  or (_18625_, _18624_, _18621_);
  and (_18626_, _18625_, _01886_);
  or (_26836_, _18626_, _18618_);
  and (_18627_, _09507_, _23693_);
  and (_18628_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_10114_, _18628_, _18627_);
  and (_18629_, _25440_, _23693_);
  and (_18630_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or (_10116_, _18630_, _18629_);
  or (_18631_, _18488_, _00443_);
  or (_18632_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_18633_, _18632_, _22773_);
  and (_10119_, _18633_, _18631_);
  and (_18634_, _17190_, _23983_);
  and (_18635_, _17192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_10121_, _18635_, _18634_);
  and (_18636_, _17216_, _24053_);
  and (_18637_, _17218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_10124_, _18637_, _18636_);
  and (_18638_, _24062_, _24053_);
  and (_18639_, _24064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_10126_, _18639_, _18638_);
  and (_18640_, _18215_, _24053_);
  and (_18641_, _18217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or (_27304_, _18641_, _18640_);
  nand (_18642_, _24518_, _23759_);
  or (_18643_, _23759_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_18644_, _18643_, _22773_);
  and (_26835_[7], _18644_, _18642_);
  and (_18645_, _25440_, _23920_);
  and (_18646_, _25442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or (_27207_, _18646_, _18645_);
  and (_18647_, _18245_, _24027_);
  and (_18648_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_10133_, _18648_, _18647_);
  and (_18649_, _01952_, _24027_);
  and (_18650_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or (_10135_, _18650_, _18649_);
  or (_18651_, _05452_, _04227_);
  and (_18652_, _18651_, _24646_);
  or (_18653_, _05453_, _04975_);
  or (_18654_, _18653_, _18652_);
  or (_18655_, _18654_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_18656_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _22781_);
  and (_18657_, _18656_, _22773_);
  and (_26840_[2], _18657_, _18655_);
  and (_18658_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18659_, _25929_, _23760_);
  or (_18660_, _18659_, _18658_);
  or (_18661_, _18660_, _05450_);
  and (_26839_[2], _18661_, _22773_);
  and (_18662_, _04207_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_18663_, _04949_, _03607_);
  or (_18664_, _18663_, _06146_);
  or (_18665_, _05771_, _04213_);
  or (_18666_, _25891_, _25880_);
  or (_18667_, _18666_, _18665_);
  or (_18668_, _18667_, _06105_);
  or (_18669_, _18668_, _18664_);
  or (_18670_, _06143_, _04225_);
  or (_18671_, _18670_, _18669_);
  and (_18672_, _18671_, _01886_);
  or (_26842_[3], _18672_, _18662_);
  and (_18673_, _17184_, _23900_);
  and (_18674_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_10142_, _18674_, _18673_);
  and (_18675_, _01952_, _23900_);
  and (_18676_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or (_10143_, _18676_, _18675_);
  or (_18677_, _18488_, _00352_);
  or (_18678_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_18679_, _18678_, _22773_);
  and (_10146_, _18679_, _18677_);
  and (_18680_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_18681_, _18474_, _00183_);
  or (_18682_, _18681_, _18680_);
  or (_18683_, _18682_, _03856_);
  nand (_18684_, _03856_, _00815_);
  and (_18685_, _18684_, _22773_);
  and (_10147_, _18685_, _18683_);
  and (_18686_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_18687_, _18474_, _00564_);
  or (_18688_, _18687_, _18686_);
  or (_18689_, _18688_, _03856_);
  or (_18690_, _18478_, _01086_);
  and (_18691_, _18690_, _22773_);
  and (_10149_, _18691_, _18689_);
  and (_18692_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_18693_, _18474_, _00443_);
  or (_18694_, _18693_, _18692_);
  or (_18695_, _18694_, _03856_);
  or (_18696_, _18478_, _01021_);
  and (_18697_, _18696_, _22773_);
  and (_10151_, _18697_, _18695_);
  and (_18698_, _17099_, _23715_);
  and (_18699_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_10157_, _18699_, _18698_);
  and (_18700_, _18245_, _23983_);
  and (_18701_, _18247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_10159_, _18701_, _18700_);
  and (_18702_, _17184_, _23920_);
  and (_18703_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or (_10161_, _18703_, _18702_);
  and (_18704_, _18209_, _23751_);
  and (_18705_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_10163_, _18705_, _18704_);
  and (_18706_, _18469_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_18707_, _18474_, _26798_);
  or (_18708_, _18707_, _18706_);
  or (_18709_, _18708_, _03856_);
  or (_18710_, _18478_, _00691_);
  and (_18711_, _18710_, _22773_);
  and (_10165_, _18711_, _18709_);
  or (_18712_, _18488_, _00183_);
  or (_18713_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_18714_, _18713_, _22773_);
  and (_10167_, _18714_, _18712_);
  and (_18715_, _17184_, _23983_);
  and (_18716_, _17186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or (_10169_, _18716_, _18715_);
  and (_18717_, _17099_, _24027_);
  and (_18718_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_27214_, _18718_, _18717_);
  nor (_18719_, _24341_, _03380_);
  or (_18720_, _18719_, _03242_);
  and (_18721_, _18720_, _26282_);
  or (_18722_, _26283_, _26282_);
  nor (_18723_, _18722_, _23681_);
  and (_18724_, _26285_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_18725_, _18724_, _25513_);
  or (_18726_, _18725_, _18723_);
  or (_18727_, _18726_, _18721_);
  nand (_18728_, _25517_, _23976_);
  and (_18729_, _18728_, _22773_);
  and (_10174_, _18729_, _18727_);
  and (_18730_, _08435_, _23983_);
  and (_18731_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or (_26914_, _18731_, _18730_);
  and (_18732_, _18209_, _23693_);
  and (_18733_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_10179_, _18733_, _18732_);
  or (_18734_, _18488_, _00101_);
  or (_18735_, _18490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_18736_, _18735_, _22773_);
  and (_10182_, _18736_, _18734_);
  and (_18737_, _18209_, _23920_);
  and (_18738_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_10185_, _18738_, _18737_);
  and (_18739_, _02779_, _23983_);
  and (_18740_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_10194_, _18740_, _18739_);
  and (_18741_, _17177_, _24053_);
  and (_18742_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or (_10197_, _18742_, _18741_);
  and (_18743_, _15225_, _23983_);
  and (_18744_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_10201_, _18744_, _18743_);
  and (_18745_, _26282_, _24190_);
  nand (_18746_, _18745_, _23681_);
  or (_18747_, _18745_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_18748_, _18747_, _25514_);
  and (_18749_, _18748_, _18746_);
  or (_18750_, _18749_, _25660_);
  and (_10202_, _18750_, _22773_);
  and (_18751_, _18157_, _23751_);
  and (_18752_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or (_10216_, _18752_, _18751_);
  and (_18753_, _17177_, _23693_);
  and (_18754_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or (_10217_, _18754_, _18753_);
  and (_18755_, _18209_, _24027_);
  and (_18756_, _18211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_10228_, _18756_, _18755_);
  and (_18757_, _18157_, _23983_);
  and (_18758_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_10231_, _18758_, _18757_);
  and (_18759_, _18195_, _24053_);
  and (_18760_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or (_10232_, _18760_, _18759_);
  and (_18761_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_18762_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_18763_, _18762_, _18761_);
  and (_18764_, _18763_, _10928_);
  and (_18765_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_18766_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_18767_, _18766_, _18765_);
  and (_18768_, _18767_, _04832_);
  or (_18769_, _18768_, _18764_);
  or (_18770_, _18769_, _10926_);
  and (_18771_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_18772_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_18773_, _18772_, _18771_);
  and (_18774_, _18773_, _10928_);
  and (_18775_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and (_18776_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_18777_, _18776_, _18775_);
  and (_18778_, _18777_, _04832_);
  or (_18779_, _18778_, _18774_);
  or (_18780_, _18779_, _04868_);
  and (_18781_, _18780_, _10945_);
  and (_18782_, _18781_, _18770_);
  or (_18783_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_18784_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_18785_, _18784_, _04832_);
  and (_18786_, _18785_, _18783_);
  or (_18787_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_18788_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_18789_, _18788_, _10928_);
  and (_18790_, _18789_, _18787_);
  or (_18791_, _18790_, _18786_);
  or (_18792_, _18791_, _10926_);
  or (_18793_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_18794_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_18795_, _18794_, _04832_);
  and (_18796_, _18795_, _18793_);
  or (_18797_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_18798_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and (_18799_, _18798_, _10928_);
  and (_18800_, _18799_, _18797_);
  or (_18801_, _18800_, _18796_);
  or (_18802_, _18801_, _04868_);
  and (_18803_, _18802_, _04859_);
  and (_18804_, _18803_, _18792_);
  or (_18805_, _18804_, _18782_);
  or (_18806_, _18805_, _04849_);
  and (_18807_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_18808_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_18809_, _18808_, _04832_);
  or (_18810_, _18809_, _18807_);
  and (_18811_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_18812_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_18813_, _18812_, _10928_);
  or (_18814_, _18813_, _18811_);
  and (_18815_, _18814_, _18810_);
  or (_18816_, _18815_, _10926_);
  and (_18817_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and (_18818_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_18819_, _18818_, _04832_);
  or (_18820_, _18819_, _18817_);
  and (_18821_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_18822_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_18823_, _18822_, _10928_);
  or (_18824_, _18823_, _18821_);
  and (_18825_, _18824_, _18820_);
  or (_18826_, _18825_, _04868_);
  and (_18827_, _18826_, _10945_);
  and (_18828_, _18827_, _18816_);
  or (_18829_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_18830_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and (_18831_, _18830_, _18829_);
  or (_18832_, _18831_, _10928_);
  or (_18833_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_18834_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_18835_, _18834_, _18833_);
  or (_18836_, _18835_, _04832_);
  and (_18837_, _18836_, _18832_);
  or (_18838_, _18837_, _10926_);
  or (_18839_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_18840_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_18841_, _18840_, _18839_);
  or (_18842_, _18841_, _10928_);
  or (_18843_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_18844_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_18845_, _18844_, _18843_);
  or (_18846_, _18845_, _04832_);
  and (_18847_, _18846_, _18842_);
  or (_18848_, _18847_, _04868_);
  and (_18849_, _18848_, _04859_);
  and (_18850_, _18849_, _18838_);
  or (_18851_, _18850_, _18828_);
  or (_18852_, _18851_, _10997_);
  and (_18853_, _18852_, _10996_);
  and (_18854_, _18853_, _18806_);
  and (_18855_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_18856_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_18857_, _18856_, _18855_);
  and (_18858_, _18857_, _04832_);
  and (_18859_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_18860_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_18861_, _18860_, _18859_);
  and (_18862_, _18861_, _10928_);
  or (_18863_, _18862_, _18858_);
  and (_18864_, _18863_, _04868_);
  and (_18865_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_18866_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_18867_, _18866_, _18865_);
  and (_18868_, _18867_, _04832_);
  and (_18869_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_18870_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_18871_, _18870_, _18869_);
  and (_18872_, _18871_, _10928_);
  or (_18873_, _18872_, _18868_);
  and (_18874_, _18873_, _10926_);
  or (_18875_, _18874_, _18864_);
  and (_18876_, _18875_, _10945_);
  or (_18877_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_18878_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_18879_, _18878_, _18877_);
  and (_18880_, _18879_, _04832_);
  or (_18881_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_18882_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_18883_, _18882_, _18881_);
  and (_18884_, _18883_, _10928_);
  or (_18885_, _18884_, _18880_);
  and (_18886_, _18885_, _04868_);
  or (_18887_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_18888_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_18889_, _18888_, _18887_);
  and (_18890_, _18889_, _04832_);
  or (_18891_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_18892_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_18893_, _18892_, _18891_);
  and (_18894_, _18893_, _10928_);
  or (_18895_, _18894_, _18890_);
  and (_18896_, _18895_, _10926_);
  or (_18897_, _18896_, _18886_);
  and (_18898_, _18897_, _04859_);
  or (_18899_, _18898_, _18876_);
  and (_18900_, _18899_, _10997_);
  and (_18901_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_18902_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_18903_, _18902_, _18901_);
  and (_18904_, _18903_, _04832_);
  and (_18905_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_18906_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_18907_, _18906_, _18905_);
  and (_18908_, _18907_, _10928_);
  or (_18909_, _18908_, _18904_);
  and (_18910_, _18909_, _04868_);
  and (_18911_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_18912_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_18913_, _18912_, _18911_);
  and (_18914_, _18913_, _04832_);
  and (_18915_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and (_18916_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_18917_, _18916_, _18915_);
  and (_18918_, _18917_, _10928_);
  or (_18919_, _18918_, _18914_);
  and (_18920_, _18919_, _10926_);
  or (_18921_, _18920_, _18910_);
  and (_18922_, _18921_, _10945_);
  or (_18923_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_18924_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and (_18925_, _18924_, _18923_);
  and (_18926_, _18925_, _04832_);
  or (_18927_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_18928_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_18929_, _18928_, _18927_);
  and (_18930_, _18929_, _10928_);
  or (_18931_, _18930_, _18926_);
  and (_18932_, _18931_, _04868_);
  or (_18933_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_18934_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_18935_, _18934_, _18933_);
  and (_18936_, _18935_, _04832_);
  or (_18937_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_18938_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_18939_, _18938_, _18937_);
  and (_18940_, _18939_, _10928_);
  or (_18941_, _18940_, _18936_);
  and (_18942_, _18941_, _10926_);
  or (_18943_, _18942_, _18932_);
  and (_18944_, _18943_, _04859_);
  or (_18945_, _18944_, _18922_);
  and (_18946_, _18945_, _04849_);
  or (_18947_, _18946_, _18900_);
  and (_18948_, _18947_, _04839_);
  or (_18949_, _18948_, _18854_);
  or (_18950_, _18949_, _04843_);
  and (_18951_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_18952_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_18953_, _18952_, _18951_);
  and (_18954_, _18953_, _04832_);
  and (_18955_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and (_18956_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_18957_, _18956_, _18955_);
  and (_18958_, _18957_, _10928_);
  or (_18959_, _18958_, _18954_);
  or (_18960_, _18959_, _10926_);
  and (_18961_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_18962_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_18963_, _18962_, _18961_);
  and (_18964_, _18963_, _04832_);
  and (_18965_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_18966_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_18967_, _18966_, _18965_);
  and (_18968_, _18967_, _10928_);
  or (_18969_, _18968_, _18964_);
  or (_18970_, _18969_, _04868_);
  and (_18971_, _18970_, _10945_);
  and (_18972_, _18971_, _18960_);
  or (_18973_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_18974_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and (_18975_, _18974_, _10928_);
  and (_18976_, _18975_, _18973_);
  or (_18977_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_18978_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_18979_, _18978_, _04832_);
  and (_18980_, _18979_, _18977_);
  or (_18981_, _18980_, _18976_);
  or (_18982_, _18981_, _10926_);
  or (_18983_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_18984_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and (_18985_, _18984_, _10928_);
  and (_18986_, _18985_, _18983_);
  or (_18987_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_18988_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_18989_, _18988_, _04832_);
  and (_18990_, _18989_, _18987_);
  or (_18991_, _18990_, _18986_);
  or (_18992_, _18991_, _04868_);
  and (_18993_, _18992_, _04859_);
  and (_18994_, _18993_, _18982_);
  or (_18995_, _18994_, _18972_);
  and (_18996_, _18995_, _10997_);
  and (_18997_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_18998_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_18999_, _18998_, _18997_);
  and (_19000_, _18999_, _04832_);
  and (_19001_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_19002_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_19003_, _19002_, _19001_);
  and (_19004_, _19003_, _10928_);
  or (_19005_, _19004_, _19000_);
  or (_19006_, _19005_, _10926_);
  and (_19007_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_19008_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_19009_, _19008_, _19007_);
  and (_19010_, _19009_, _04832_);
  and (_19011_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_19012_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_19013_, _19012_, _19011_);
  and (_19014_, _19013_, _10928_);
  or (_19015_, _19014_, _19010_);
  or (_19016_, _19015_, _04868_);
  and (_19017_, _19016_, _10945_);
  and (_19018_, _19017_, _19006_);
  or (_19019_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_19020_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_19021_, _19020_, _19019_);
  and (_19022_, _19021_, _04832_);
  or (_19023_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_19024_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_19025_, _19024_, _19023_);
  and (_19026_, _19025_, _10928_);
  or (_19027_, _19026_, _19022_);
  or (_19028_, _19027_, _10926_);
  or (_19029_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_19030_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_19031_, _19030_, _19029_);
  and (_19032_, _19031_, _04832_);
  or (_19033_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_19034_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_19035_, _19034_, _19033_);
  and (_19036_, _19035_, _10928_);
  or (_19037_, _19036_, _19032_);
  or (_19038_, _19037_, _04868_);
  and (_19039_, _19038_, _04859_);
  and (_19040_, _19039_, _19028_);
  or (_19041_, _19040_, _19018_);
  and (_19042_, _19041_, _04849_);
  or (_19043_, _19042_, _18996_);
  and (_19044_, _19043_, _10996_);
  or (_19045_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_19046_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_19047_, _19046_, _19045_);
  and (_19048_, _19047_, _04832_);
  or (_19049_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_19050_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and (_19051_, _19050_, _19049_);
  and (_19052_, _19051_, _10928_);
  or (_19053_, _19052_, _19048_);
  and (_19054_, _19053_, _10926_);
  or (_19055_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_19056_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_19057_, _19056_, _19055_);
  and (_19058_, _19057_, _04832_);
  or (_19059_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_19060_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_19061_, _19060_, _19059_);
  and (_19062_, _19061_, _10928_);
  or (_19063_, _19062_, _19058_);
  and (_19064_, _19063_, _04868_);
  or (_19065_, _19064_, _19054_);
  and (_19066_, _19065_, _04859_);
  and (_19067_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and (_19068_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_19069_, _19068_, _19067_);
  and (_19070_, _19069_, _04832_);
  and (_19071_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_19072_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_19073_, _19072_, _19071_);
  and (_19074_, _19073_, _10928_);
  or (_19075_, _19074_, _19070_);
  and (_19076_, _19075_, _10926_);
  and (_19077_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_19078_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_19079_, _19078_, _19077_);
  and (_19080_, _19079_, _04832_);
  and (_19081_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_19082_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_19083_, _19082_, _19081_);
  and (_19084_, _19083_, _10928_);
  or (_19085_, _19084_, _19080_);
  and (_19086_, _19085_, _04868_);
  or (_19087_, _19086_, _19076_);
  and (_19088_, _19087_, _10945_);
  or (_19089_, _19088_, _19066_);
  and (_19090_, _19089_, _04849_);
  or (_19091_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_19092_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and (_19093_, _19092_, _10928_);
  and (_19094_, _19093_, _19091_);
  or (_19095_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_19096_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and (_19097_, _19096_, _04832_);
  and (_19098_, _19097_, _19095_);
  or (_19099_, _19098_, _19094_);
  and (_19100_, _19099_, _10926_);
  or (_19101_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_19102_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_19103_, _19102_, _10928_);
  and (_19104_, _19103_, _19101_);
  or (_19105_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_19106_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and (_19107_, _19106_, _04832_);
  and (_19108_, _19107_, _19105_);
  or (_19109_, _19108_, _19104_);
  and (_19110_, _19109_, _04868_);
  or (_19111_, _19110_, _19100_);
  and (_19112_, _19111_, _04859_);
  and (_19113_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and (_19114_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_19115_, _19114_, _19113_);
  and (_19116_, _19115_, _04832_);
  and (_19117_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_19118_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_19119_, _19118_, _19117_);
  and (_19120_, _19119_, _10928_);
  or (_19121_, _19120_, _19116_);
  and (_19122_, _19121_, _10926_);
  and (_19123_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and (_19124_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_19125_, _19124_, _19123_);
  and (_19126_, _19125_, _04832_);
  and (_19127_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_19128_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_19129_, _19128_, _19127_);
  and (_19130_, _19129_, _10928_);
  or (_19131_, _19130_, _19126_);
  and (_19132_, _19131_, _04868_);
  or (_19133_, _19132_, _19122_);
  and (_19134_, _19133_, _10945_);
  or (_19135_, _19134_, _19112_);
  and (_19136_, _19135_, _10997_);
  or (_19137_, _19136_, _19090_);
  and (_19138_, _19137_, _04839_);
  or (_19139_, _19138_, _19044_);
  or (_19140_, _19139_, _11204_);
  and (_19141_, _19140_, _18950_);
  or (_19142_, _19141_, _26153_);
  and (_19143_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_19144_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_19145_, _19144_, _19143_);
  and (_19146_, _19145_, _10928_);
  and (_19147_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_19148_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_19149_, _19148_, _19147_);
  and (_19150_, _19149_, _04832_);
  or (_19151_, _19150_, _19146_);
  or (_19152_, _19151_, _10926_);
  and (_19153_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_19154_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_19155_, _19154_, _19153_);
  and (_19156_, _19155_, _10928_);
  and (_19157_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_19158_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_19159_, _19158_, _19157_);
  and (_19160_, _19159_, _04832_);
  or (_19161_, _19160_, _19156_);
  or (_19162_, _19161_, _04868_);
  and (_19163_, _19162_, _10945_);
  and (_19164_, _19163_, _19152_);
  or (_19165_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_19166_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_19167_, _19166_, _04832_);
  and (_19168_, _19167_, _19165_);
  or (_19169_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_19170_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_19171_, _19170_, _10928_);
  and (_19172_, _19171_, _19169_);
  or (_19173_, _19172_, _19168_);
  or (_19174_, _19173_, _10926_);
  or (_19175_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_19176_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_19177_, _19176_, _04832_);
  and (_19178_, _19177_, _19175_);
  or (_19179_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_19180_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_19181_, _19180_, _10928_);
  and (_19182_, _19181_, _19179_);
  or (_19183_, _19182_, _19178_);
  or (_19184_, _19183_, _04868_);
  and (_19185_, _19184_, _04859_);
  and (_19186_, _19185_, _19174_);
  or (_19187_, _19186_, _19164_);
  and (_19188_, _19187_, _10997_);
  and (_19189_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_19190_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_19191_, _19190_, _04832_);
  or (_19192_, _19191_, _19189_);
  and (_19193_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_19194_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_19195_, _19194_, _10928_);
  or (_19196_, _19195_, _19193_);
  and (_19197_, _19196_, _19192_);
  or (_19198_, _19197_, _10926_);
  and (_19199_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_19200_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_19201_, _19200_, _04832_);
  or (_19202_, _19201_, _19199_);
  and (_19203_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_19204_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_19205_, _19204_, _10928_);
  or (_19206_, _19205_, _19203_);
  and (_19207_, _19206_, _19202_);
  or (_19208_, _19207_, _04868_);
  and (_19209_, _19208_, _10945_);
  and (_19210_, _19209_, _19198_);
  or (_19211_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_19212_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_19213_, _19212_, _19211_);
  or (_19214_, _19213_, _10928_);
  or (_19215_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_19216_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_19217_, _19216_, _19215_);
  or (_19218_, _19217_, _04832_);
  and (_19219_, _19218_, _19214_);
  or (_19220_, _19219_, _10926_);
  or (_19221_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_19222_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_19223_, _19222_, _19221_);
  or (_19224_, _19223_, _10928_);
  or (_19225_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_19226_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_19227_, _19226_, _19225_);
  or (_19228_, _19227_, _04832_);
  and (_19229_, _19228_, _19224_);
  or (_19230_, _19229_, _04868_);
  and (_19231_, _19230_, _04859_);
  and (_19232_, _19231_, _19220_);
  or (_19233_, _19232_, _19210_);
  and (_19234_, _19233_, _04849_);
  or (_19235_, _19234_, _19188_);
  and (_19236_, _19235_, _10996_);
  and (_19237_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  and (_19238_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  or (_19239_, _19238_, _19237_);
  and (_19240_, _19239_, _04832_);
  and (_19241_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  and (_19242_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or (_19243_, _19242_, _19241_);
  and (_19244_, _19243_, _10928_);
  or (_19245_, _19244_, _19240_);
  and (_19246_, _19245_, _04868_);
  and (_19247_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  and (_19248_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or (_19249_, _19248_, _19247_);
  and (_19250_, _19249_, _04832_);
  and (_19251_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  and (_19252_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  or (_19253_, _19252_, _19251_);
  and (_19254_, _19253_, _10928_);
  or (_19255_, _19254_, _19250_);
  and (_19256_, _19255_, _10926_);
  or (_19257_, _19256_, _19246_);
  and (_19258_, _19257_, _10945_);
  or (_19259_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  or (_19260_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  and (_19261_, _19260_, _19259_);
  and (_19262_, _19261_, _04832_);
  or (_19263_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  or (_19264_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and (_19265_, _19264_, _19263_);
  and (_19266_, _19265_, _10928_);
  or (_19267_, _19266_, _19262_);
  and (_19268_, _19267_, _04868_);
  or (_19269_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or (_19270_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  and (_19271_, _19270_, _19269_);
  and (_19272_, _19271_, _04832_);
  or (_19273_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or (_19274_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and (_19275_, _19274_, _19273_);
  and (_19276_, _19275_, _10928_);
  or (_19277_, _19276_, _19272_);
  and (_19278_, _19277_, _10926_);
  or (_19279_, _19278_, _19268_);
  and (_19280_, _19279_, _04859_);
  or (_19281_, _19280_, _19258_);
  and (_19282_, _19281_, _10997_);
  and (_19283_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_19284_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_19285_, _19284_, _19283_);
  and (_19286_, _19285_, _04832_);
  and (_19287_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_19288_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_19289_, _19288_, _19287_);
  and (_19290_, _19289_, _10928_);
  or (_19291_, _19290_, _19286_);
  and (_19292_, _19291_, _04868_);
  and (_19293_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_19294_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_19295_, _19294_, _19293_);
  and (_19296_, _19295_, _04832_);
  and (_19297_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_19298_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_19299_, _19298_, _19297_);
  and (_19300_, _19299_, _10928_);
  or (_19301_, _19300_, _19296_);
  and (_19302_, _19301_, _10926_);
  or (_19303_, _19302_, _19292_);
  and (_19304_, _19303_, _10945_);
  or (_19305_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_19306_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_19307_, _19306_, _19305_);
  and (_19308_, _19307_, _04832_);
  or (_19309_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_19310_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_19311_, _19310_, _19309_);
  and (_19312_, _19311_, _10928_);
  or (_19313_, _19312_, _19308_);
  and (_19314_, _19313_, _04868_);
  or (_19315_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_19316_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_19317_, _19316_, _19315_);
  and (_19318_, _19317_, _04832_);
  or (_19319_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_19320_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_19321_, _19320_, _19319_);
  and (_19322_, _19321_, _10928_);
  or (_19323_, _19322_, _19318_);
  and (_19324_, _19323_, _10926_);
  or (_19325_, _19324_, _19314_);
  and (_19326_, _19325_, _04859_);
  or (_19327_, _19326_, _19304_);
  and (_19328_, _19327_, _04849_);
  or (_19329_, _19328_, _19282_);
  and (_19330_, _19329_, _04839_);
  or (_19331_, _19330_, _19236_);
  or (_19332_, _19331_, _04843_);
  and (_19333_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_19334_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_19335_, _19334_, _19333_);
  and (_19336_, _19335_, _04832_);
  and (_19337_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_19338_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_19339_, _19338_, _19337_);
  and (_19340_, _19339_, _10928_);
  or (_19341_, _19340_, _19336_);
  or (_19342_, _19341_, _10926_);
  and (_19343_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_19344_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_19345_, _19344_, _19343_);
  and (_19346_, _19345_, _04832_);
  and (_19347_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_19348_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_19349_, _19348_, _19347_);
  and (_19350_, _19349_, _10928_);
  or (_19351_, _19350_, _19346_);
  or (_19352_, _19351_, _04868_);
  and (_19353_, _19352_, _10945_);
  and (_19354_, _19353_, _19342_);
  or (_19355_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_19356_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_19357_, _19356_, _10928_);
  and (_19358_, _19357_, _19355_);
  or (_19359_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_19360_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_19361_, _19360_, _04832_);
  and (_19362_, _19361_, _19359_);
  or (_19363_, _19362_, _19358_);
  or (_19364_, _19363_, _10926_);
  or (_19365_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_19366_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_19367_, _19366_, _10928_);
  and (_19368_, _19367_, _19365_);
  or (_19369_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_19370_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_19371_, _19370_, _04832_);
  and (_19372_, _19371_, _19369_);
  or (_19373_, _19372_, _19368_);
  or (_19374_, _19373_, _04868_);
  and (_19375_, _19374_, _04859_);
  and (_19376_, _19375_, _19364_);
  or (_19377_, _19376_, _19354_);
  and (_19378_, _19377_, _10997_);
  and (_19379_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_19380_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_19381_, _19380_, _19379_);
  and (_19382_, _19381_, _04832_);
  and (_19383_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_19384_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_19385_, _19384_, _19383_);
  and (_19386_, _19385_, _10928_);
  or (_19387_, _19386_, _19382_);
  or (_19388_, _19387_, _10926_);
  and (_19389_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_19390_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_19391_, _19390_, _19389_);
  and (_19392_, _19391_, _04832_);
  and (_19393_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_19394_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_19395_, _19394_, _19393_);
  and (_19396_, _19395_, _10928_);
  or (_19397_, _19396_, _19392_);
  or (_19398_, _19397_, _04868_);
  and (_19399_, _19398_, _10945_);
  and (_19400_, _19399_, _19388_);
  or (_19401_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_19402_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_19403_, _19402_, _19401_);
  and (_19404_, _19403_, _04832_);
  or (_19405_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_19406_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_19407_, _19406_, _19405_);
  and (_19408_, _19407_, _10928_);
  or (_19409_, _19408_, _19404_);
  or (_19410_, _19409_, _10926_);
  or (_19411_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_19412_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_19413_, _19412_, _19411_);
  and (_19414_, _19413_, _04832_);
  or (_19415_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_19416_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_19417_, _19416_, _19415_);
  and (_19418_, _19417_, _10928_);
  or (_19419_, _19418_, _19414_);
  or (_19420_, _19419_, _04868_);
  and (_19421_, _19420_, _04859_);
  and (_19422_, _19421_, _19410_);
  or (_19423_, _19422_, _19400_);
  and (_19424_, _19423_, _04849_);
  or (_19425_, _19424_, _19378_);
  and (_19426_, _19425_, _10996_);
  or (_19427_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_19428_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_19429_, _19428_, _19427_);
  and (_19430_, _19429_, _04832_);
  or (_19431_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_19432_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_19433_, _19432_, _19431_);
  and (_19434_, _19433_, _10928_);
  or (_19435_, _19434_, _19430_);
  and (_19436_, _19435_, _10926_);
  or (_19437_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_19438_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_19439_, _19438_, _19437_);
  and (_19440_, _19439_, _04832_);
  or (_19441_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_19442_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_19443_, _19442_, _19441_);
  and (_19444_, _19443_, _10928_);
  or (_19445_, _19444_, _19440_);
  and (_19446_, _19445_, _04868_);
  or (_19447_, _19446_, _19436_);
  and (_19448_, _19447_, _04859_);
  and (_19449_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_19450_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_19451_, _19450_, _19449_);
  and (_19452_, _19451_, _04832_);
  and (_19453_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_19454_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_19455_, _19454_, _19453_);
  and (_19456_, _19455_, _10928_);
  or (_19457_, _19456_, _19452_);
  and (_19458_, _19457_, _10926_);
  and (_19459_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_19460_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_19461_, _19460_, _19459_);
  and (_19462_, _19461_, _04832_);
  and (_19463_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_19464_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_19465_, _19464_, _19463_);
  and (_19466_, _19465_, _10928_);
  or (_19467_, _19466_, _19462_);
  and (_19468_, _19467_, _04868_);
  or (_19469_, _19468_, _19458_);
  and (_19470_, _19469_, _10945_);
  or (_19471_, _19470_, _19448_);
  and (_19472_, _19471_, _04849_);
  or (_19473_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_19474_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_19475_, _19474_, _10928_);
  and (_19476_, _19475_, _19473_);
  or (_19477_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_19478_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_19479_, _19478_, _04832_);
  and (_19480_, _19479_, _19477_);
  or (_19481_, _19480_, _19476_);
  and (_19482_, _19481_, _10926_);
  or (_19483_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_19484_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_19485_, _19484_, _10928_);
  and (_19486_, _19485_, _19483_);
  or (_19487_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_19488_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_19489_, _19488_, _04832_);
  and (_19490_, _19489_, _19487_);
  or (_19491_, _19490_, _19486_);
  and (_19492_, _19491_, _04868_);
  or (_19493_, _19492_, _19482_);
  and (_19494_, _19493_, _04859_);
  and (_19495_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_19496_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_19497_, _19496_, _19495_);
  and (_19498_, _19497_, _04832_);
  and (_19499_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_19500_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_19501_, _19500_, _19499_);
  and (_19502_, _19501_, _10928_);
  or (_19503_, _19502_, _19498_);
  and (_19504_, _19503_, _10926_);
  and (_19505_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_19506_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_19507_, _19506_, _19505_);
  and (_19508_, _19507_, _04832_);
  and (_19509_, _10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_19510_, _04824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_19511_, _19510_, _19509_);
  and (_19512_, _19511_, _10928_);
  or (_19513_, _19512_, _19508_);
  and (_19514_, _19513_, _04868_);
  or (_19515_, _19514_, _19504_);
  and (_19516_, _19515_, _10945_);
  or (_19517_, _19516_, _19494_);
  and (_19518_, _19517_, _10997_);
  or (_19519_, _19518_, _19472_);
  and (_19520_, _19519_, _04839_);
  or (_19521_, _19520_, _19426_);
  or (_19522_, _19521_, _11204_);
  and (_19523_, _19522_, _19332_);
  or (_19524_, _19523_, _03196_);
  and (_19525_, _19524_, _19142_);
  or (_19526_, _19525_, _04876_);
  or (_19527_, _11878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_19528_, _19527_, _22773_);
  and (_10234_, _19528_, _19526_);
  and (_19529_, _02779_, _24027_);
  and (_19530_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_10236_, _19530_, _19529_);
  and (_19531_, _17177_, _23715_);
  and (_19532_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or (_27288_, _19532_, _19531_);
  and (_19533_, _07484_, _23900_);
  and (_19534_, _07487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_10254_, _19534_, _19533_);
  and (_19535_, _18195_, _23751_);
  and (_19536_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or (_10256_, _19536_, _19535_);
  and (_19537_, _17177_, _23900_);
  and (_19538_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or (_10258_, _19538_, _19537_);
  and (_19539_, _18195_, _23900_);
  and (_19540_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or (_10262_, _19540_, _19539_);
  and (_19541_, _17177_, _24027_);
  and (_19542_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or (_10264_, _19542_, _19541_);
  and (_19543_, _26282_, _22895_);
  nand (_19544_, _19543_, _23681_);
  not (_19545_, _25517_);
  or (_19546_, _19543_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_19547_, _19546_, _19545_);
  and (_19548_, _19547_, _19544_);
  and (_19549_, _25517_, _23744_);
  or (_19550_, _19549_, _19548_);
  and (_10266_, _19550_, _22773_);
  and (_19551_, _05834_, _23900_);
  and (_19552_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_10269_, _19552_, _19551_);
  and (_19553_, _17099_, _23920_);
  and (_19554_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_10281_, _19554_, _19553_);
  and (_19555_, _01701_, _23693_);
  and (_19556_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or (_10284_, _19556_, _19555_);
  and (_19557_, _05834_, _24053_);
  and (_19558_, _05836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_10287_, _19558_, _19557_);
  and (_19559_, _26282_, _23250_);
  nand (_19560_, _19559_, _23681_);
  or (_19561_, _19559_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_19562_, _19561_, _19545_);
  and (_19563_, _19562_, _19560_);
  or (_19564_, _19563_, _25518_);
  and (_10289_, _19564_, _22773_);
  and (_19565_, _15225_, _24053_);
  and (_19566_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_10296_, _19566_, _19565_);
  not (_19567_, _26282_);
  or (_19568_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_19569_, _00072_, _26777_);
  or (_19570_, _19569_, _00155_);
  or (_19571_, _19570_, _00250_);
  or (_19572_, _19571_, _00412_);
  or (_19573_, _19572_, _00533_);
  and (_19574_, _19573_, _26607_);
  or (_19575_, _23594_, _23591_);
  not (_19576_, _23488_);
  nand (_19577_, _23591_, _19576_);
  and (_19578_, _19577_, _23458_);
  and (_19579_, _19578_, _19575_);
  nand (_19580_, _23631_, _23599_);
  and (_19581_, _23632_, _23597_);
  and (_19582_, _19581_, _19580_);
  or (_19583_, _23545_, _23388_);
  or (_19584_, _19583_, _23554_);
  and (_19585_, _26379_, _23185_);
  and (_19586_, _23323_, _23538_);
  and (_19587_, _19586_, _19585_);
  nand (_19588_, _19587_, _26386_);
  or (_19589_, _19588_, _19584_);
  nand (_19590_, _19589_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_19591_, _19590_, _19582_);
  or (_19592_, _19591_, _19579_);
  nor (_19593_, _19592_, _00333_);
  nand (_19594_, _19593_, _00590_);
  or (_19595_, _19594_, _19574_);
  and (_19596_, _19595_, _19568_);
  and (_19597_, _19596_, _19567_);
  and (_19598_, _02022_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_19599_, _19598_, _02023_);
  and (_19600_, _19599_, _26282_);
  or (_19601_, _19600_, _19597_);
  or (_19602_, _19601_, _25517_);
  or (_19603_, _19545_, _23247_);
  and (_19604_, _19603_, _22773_);
  and (_10297_, _19604_, _19602_);
  and (_19605_, _02455_, _23693_);
  and (_19606_, _02457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or (_10299_, _19606_, _19605_);
  and (_19607_, _18195_, _23920_);
  and (_19608_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_10301_, _19608_, _19607_);
  and (_19609_, _17177_, _23983_);
  and (_19610_, _17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_10302_, _19610_, _19609_);
  and (_19611_, _17169_, _23751_);
  and (_19612_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_10321_, _19612_, _19611_);
  and (_19613_, _18195_, _23983_);
  and (_19614_, _18197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or (_10325_, _19614_, _19613_);
  and (_19615_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_19616_, _02848_, _23693_);
  or (_10332_, _19616_, _19615_);
  and (_19617_, _02789_, _23920_);
  and (_19618_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_10336_, _19618_, _19617_);
  and (_19619_, _25482_, _24053_);
  and (_19620_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_27225_, _19620_, _19619_);
  and (_19621_, _18185_, _24053_);
  and (_19622_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or (_10339_, _19622_, _19621_);
  and (_19623_, _17169_, _23693_);
  and (_19624_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_10340_, _19624_, _19623_);
  and (_19625_, _18185_, _23715_);
  and (_19626_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or (_10344_, _19626_, _19625_);
  and (_19627_, _17169_, _23920_);
  and (_19628_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_10346_, _19628_, _19627_);
  and (_19629_, _02789_, _24027_);
  and (_19630_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_10348_, _19630_, _19629_);
  and (_10350_, _03295_, _22773_);
  and (_19631_, _18185_, _23900_);
  and (_19632_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or (_10355_, _19632_, _19631_);
  and (_19633_, _15225_, _23715_);
  and (_19634_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_10357_, _19634_, _19633_);
  and (_19635_, _17169_, _24027_);
  and (_19636_, _17171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_10359_, _19636_, _19635_);
  and (_19637_, _17083_, _23920_);
  and (_19638_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or (_10362_, _19638_, _19637_);
  or (_19639_, _23253_, _23247_);
  and (_19640_, _23269_, _23268_);
  nor (_19641_, _19640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_19642_, _19641_, _10184_);
  and (_19643_, _19642_, _10189_);
  and (_19644_, _10191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand (_19645_, _24294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_19646_, _19645_, _23210_);
  or (_19647_, _19646_, _19644_);
  or (_19648_, _19647_, _19643_);
  or (_19649_, _19648_, _23252_);
  and (_19650_, _19649_, _22773_);
  and (_10366_, _19650_, _19639_);
  and (_19651_, _17163_, _24053_);
  and (_19652_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_10368_, _19652_, _19651_);
  and (_19653_, _09570_, _23983_);
  and (_19654_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_10369_, _19654_, _19653_);
  and (_19655_, _15225_, _23693_);
  and (_19656_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_10371_, _19656_, _19655_);
  and (_19657_, _18185_, _24027_);
  and (_19658_, _18187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or (_10373_, _19658_, _19657_);
  and (_19659_, _15225_, _23751_);
  and (_19660_, _15227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_10374_, _19660_, _19659_);
  or (_19661_, _24373_, _00257_);
  nand (_19662_, _19661_, _26282_);
  or (_19663_, _19662_, _03230_);
  and (_19664_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_19665_, _19664_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_19666_, _23587_, _23458_);
  and (_19667_, _23618_, _23597_);
  nand (_19668_, _23173_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_19669_, _19668_, _19664_);
  or (_19670_, _19669_, _19667_);
  or (_19671_, _19670_, _19666_);
  and (_19672_, _19671_, _19665_);
  or (_19673_, _19672_, _26282_);
  and (_19674_, _19673_, _19663_);
  or (_19675_, _19674_, _25517_);
  nand (_19676_, _25517_, _24017_);
  and (_19677_, _19676_, _22773_);
  and (_10377_, _19677_, _19675_);
  and (_19678_, _16992_, _23751_);
  and (_19679_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or (_10380_, _19679_, _19678_);
  and (_19680_, _17163_, _23751_);
  and (_19681_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_10386_, _19681_, _19680_);
  and (_19682_, _16992_, _24027_);
  and (_19683_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or (_10388_, _19683_, _19682_);
  and (_19684_, _17163_, _23920_);
  and (_19685_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_10389_, _19685_, _19684_);
  and (_19686_, _17083_, _24053_);
  and (_19687_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or (_10391_, _19687_, _19686_);
  and (_19688_, _18175_, _23693_);
  and (_19689_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_10393_, _19689_, _19688_);
  and (_19690_, _26282_, _23208_);
  and (_19691_, _19690_, _23681_);
  nor (_19692_, _19690_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_19693_, _19692_, _19691_);
  nand (_19694_, _19693_, _19545_);
  nand (_19695_, _25517_, _23357_);
  and (_19696_, _19695_, _22773_);
  and (_10394_, _19696_, _19694_);
  and (_19697_, _02779_, _23751_);
  and (_19698_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_27131_, _19698_, _19697_);
  and (_19699_, _01745_, _23983_);
  and (_19700_, _01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or (_10397_, _19700_, _19699_);
  and (_19701_, _16720_, _24053_);
  and (_19702_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_10401_, _19702_, _19701_);
  and (_10406_, _03223_, _22773_);
  and (_19703_, _17083_, _23900_);
  and (_19704_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or (_10408_, _19704_, _19703_);
  and (_19705_, _18175_, _23900_);
  and (_19706_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_10423_, _19706_, _19705_);
  and (_10438_, _03326_, _22773_);
  and (_19707_, _09485_, _23900_);
  and (_19708_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_27037_, _19708_, _19707_);
  and (_19709_, _17083_, _24027_);
  and (_19710_, _17085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or (_27235_, _19710_, _19709_);
  and (_19711_, _02509_, _23715_);
  and (_19712_, _02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_10460_, _19712_, _19711_);
  and (_10465_, _03341_, _22773_);
  and (_19713_, _17163_, _24027_);
  and (_19714_, _17165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_10468_, _19714_, _19713_);
  and (_10484_, _03212_, _22773_);
  nor (_10486_, _03354_, rst);
  and (_19715_, _02779_, _24053_);
  and (_19716_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_10492_, _19716_, _19715_);
  and (_19717_, _16720_, _23900_);
  and (_19718_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_10493_, _19718_, _19717_);
  and (_19719_, _17157_, _24053_);
  and (_19720_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or (_10508_, _19720_, _19719_);
  and (_19721_, _10525_, _23900_);
  and (_19722_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or (_10518_, _19722_, _19721_);
  and (_19723_, _09570_, _24027_);
  and (_19724_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_10529_, _19724_, _19723_);
  and (_19725_, _09485_, _23715_);
  and (_19726_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_10530_, _19726_, _19725_);
  and (_19727_, _18175_, _23920_);
  and (_19728_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_10535_, _19728_, _19727_);
  and (_19729_, _10525_, _23751_);
  and (_19730_, _10527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or (_10540_, _19730_, _19729_);
  and (_19731_, _18175_, _23983_);
  and (_19732_, _18177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_10555_, _19732_, _19731_);
  and (_19733_, _09485_, _23693_);
  and (_19734_, _09487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_10557_, _19734_, _19733_);
  and (_19735_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_19736_, _02848_, _23751_);
  or (_10559_, _19736_, _19735_);
  and (_19737_, _09552_, _23693_);
  and (_19738_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_10560_, _19738_, _19737_);
  and (_19739_, _16720_, _23920_);
  and (_19740_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_10571_, _19740_, _19739_);
  and (_19741_, _17157_, _23751_);
  and (_19742_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or (_10572_, _19742_, _19741_);
  and (_19743_, _16720_, _23983_);
  and (_19744_, _16722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_26892_, _19744_, _19743_);
  and (_10578_, _03313_, _22773_);
  and (_19745_, _17157_, _23900_);
  and (_19746_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or (_10582_, _19746_, _19745_);
  and (_19747_, _05883_, _23693_);
  and (_19748_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_10587_, _19748_, _19747_);
  and (_10589_, _03239_, _22773_);
  and (_19749_, _09552_, _23983_);
  and (_19750_, _09554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_10596_, _19750_, _19749_);
  and (_19751_, _18167_, _24053_);
  and (_19752_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_27309_, _19752_, _19751_);
  and (_19753_, _17157_, _23920_);
  and (_19754_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or (_10607_, _19754_, _19753_);
  and (_19755_, _05883_, _23920_);
  and (_19756_, _05886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_10608_, _19756_, _19755_);
  and (_19757_, _16988_, _23920_);
  and (_19758_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_10613_, _19758_, _19757_);
  and (_19759_, _08435_, _24027_);
  and (_19760_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or (_10614_, _19760_, _19759_);
  and (_19761_, _15229_, _23693_);
  and (_19762_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or (_10618_, _19762_, _19761_);
  and (_19763_, _17017_, _24053_);
  and (_19764_, _17019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_10621_, _19764_, _19763_);
  and (_19765_, _05731_, _23983_);
  and (_19766_, _05733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or (_10623_, _19766_, _19765_);
  and (_19767_, _18167_, _23751_);
  and (_19768_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_27310_, _19768_, _19767_);
  and (_19769_, _17157_, _23983_);
  and (_19770_, _17159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_10626_, _19770_, _19769_);
  and (_19771_, _16632_, _24053_);
  and (_19772_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_10627_, _19772_, _19771_);
  and (_19773_, _15229_, _23751_);
  and (_19774_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or (_10630_, _19774_, _19773_);
  and (_19775_, _18167_, _23715_);
  and (_19776_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_10633_, _19776_, _19775_);
  and (_19777_, _02244_, _24027_);
  and (_19778_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or (_27245_, _19778_, _19777_);
  nand (_19779_, _24017_, _23252_);
  and (_19780_, _24287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_19781_, _23268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_19782_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_19783_, _19782_, _24289_);
  and (_19784_, _24284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_19785_, _19784_, _23275_);
  or (_19786_, _19785_, _19783_);
  and (_19787_, _19786_, _19781_);
  and (_19788_, _19787_, _24286_);
  or (_19789_, _19788_, _19780_);
  or (_19790_, _19789_, _23252_);
  and (_19791_, _19790_, _22773_);
  and (_10635_, _19791_, _19779_);
  and (_19792_, _17151_, _24053_);
  and (_19793_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or (_10638_, _19793_, _19792_);
  and (_19794_, _24242_, _24027_);
  and (_19795_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or (_10640_, _19795_, _19794_);
  and (_19796_, _17151_, _23715_);
  and (_19797_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or (_10645_, _19797_, _19796_);
  and (_19798_, _18167_, _23920_);
  and (_19799_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_10653_, _19799_, _19798_);
  and (_19800_, _24242_, _23983_);
  and (_19801_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_26887_, _19801_, _19800_);
  and (_19802_, _16710_, _24053_);
  and (_19803_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or (_26888_, _19803_, _19802_);
  and (_19804_, _16988_, _23900_);
  and (_19805_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_10659_, _19805_, _19804_);
  and (_19806_, _18167_, _23983_);
  and (_19807_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_10660_, _19807_, _19806_);
  and (_19808_, _23988_, _23693_);
  and (_19809_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_10664_, _19809_, _19808_);
  and (_19810_, _17151_, _23900_);
  and (_19811_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or (_10665_, _19811_, _19810_);
  and (_19812_, _16988_, _23715_);
  and (_19813_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_10668_, _19813_, _19812_);
  and (_19814_, _17151_, _24027_);
  and (_19815_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or (_27291_, _19815_, _19814_);
  and (_19816_, _18163_, _24053_);
  and (_19817_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or (_10676_, _19817_, _19816_);
  and (_19818_, _23988_, _23920_);
  and (_19819_, _23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_10679_, _19819_, _19818_);
  and (_19820_, _18163_, _23693_);
  and (_19821_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or (_10680_, _19821_, _19820_);
  and (_19822_, _16710_, _23751_);
  and (_19823_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or (_10686_, _19823_, _19822_);
  and (_19824_, _09463_, _23693_);
  and (_19825_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_10688_, _19825_, _19824_);
  and (_19826_, _17099_, _23983_);
  and (_19827_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_27215_, _19827_, _19826_);
  and (_19828_, _17151_, _23983_);
  and (_19829_, _17153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or (_10691_, _19829_, _19828_);
  and (_19830_, _04771_, _23900_);
  and (_19831_, _04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_27251_, _19831_, _19830_);
  and (_19832_, _18163_, _23900_);
  and (_19833_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or (_10694_, _19833_, _19832_);
  and (_19834_, _16710_, _23900_);
  and (_19835_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or (_10696_, _19835_, _19834_);
  and (_19836_, _17147_, _23751_);
  and (_19837_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_10700_, _19837_, _19836_);
  and (_19838_, _02326_, _23693_);
  and (_19839_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or (_10701_, _19839_, _19838_);
  and (_19840_, _09463_, _23751_);
  and (_19841_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_10704_, _19841_, _19840_);
  and (_19842_, _16710_, _23920_);
  and (_19843_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or (_10707_, _19843_, _19842_);
  and (_19844_, _17069_, _23693_);
  and (_19845_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_27255_, _19845_, _19844_);
  and (_19846_, _09463_, _24053_);
  and (_19847_, _09466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_10712_, _19847_, _19846_);
  and (_19848_, _18163_, _23920_);
  and (_19849_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or (_27312_, _19849_, _19848_);
  and (_19850_, _17147_, _23693_);
  and (_19851_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_10715_, _19851_, _19850_);
  and (_19852_, _02326_, _24053_);
  and (_19853_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or (_27252_, _19853_, _19852_);
  and (_19854_, _18163_, _23983_);
  and (_19855_, _18165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_27313_, _19855_, _19854_);
  and (_19856_, _17059_, _24053_);
  and (_19857_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_10725_, _19857_, _19856_);
  and (_19858_, _17147_, _23715_);
  and (_19859_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_10732_, _19859_, _19858_);
  and (_19860_, _17069_, _24027_);
  and (_19861_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_10735_, _19861_, _19860_);
  and (_19862_, _24231_, _24053_);
  and (_19863_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or (_10737_, _19863_, _19862_);
  and (_19864_, _17147_, _23920_);
  and (_19865_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_10739_, _19865_, _19864_);
  and (_19866_, _17059_, _24027_);
  and (_19867_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_10741_, _19867_, _19866_);
  and (_19868_, _17059_, _23715_);
  and (_19869_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_10744_, _19869_, _19868_);
  and (_19870_, _16988_, _23983_);
  and (_19871_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_27234_, _19871_, _19870_);
  and (_19872_, _16710_, _23983_);
  and (_19873_, _16712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or (_10748_, _19873_, _19872_);
  and (_19874_, _16688_, _24053_);
  and (_19875_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_10750_, _19875_, _19874_);
  and (_19876_, _16988_, _24027_);
  and (_19877_, _16990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_10753_, _19877_, _19876_);
  and (_19878_, _02794_, _23983_);
  and (_19879_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or (_10762_, _19879_, _19878_);
  and (_19880_, _16688_, _23693_);
  and (_19881_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_10763_, _19881_, _19880_);
  and (_19882_, _16688_, _23900_);
  and (_19883_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_10767_, _19883_, _19882_);
  and (_19884_, _02829_, _23920_);
  and (_19885_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or (_10769_, _19885_, _19884_);
  and (_19886_, _02350_, _23715_);
  and (_19887_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_10773_, _19887_, _19886_);
  and (_19888_, _15229_, _23920_);
  and (_19889_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or (_26929_, _19889_, _19888_);
  and (_19890_, _02789_, _24053_);
  and (_19891_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_10778_, _19891_, _19890_);
  and (_19892_, _15229_, _23900_);
  and (_19893_, _15231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or (_26928_, _19893_, _19892_);
  and (_19894_, _02849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_19895_, _02848_, _23900_);
  or (_10783_, _19895_, _19894_);
  and (_19896_, _16688_, _23920_);
  and (_19897_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_10786_, _19897_, _19896_);
  and (_19898_, _16688_, _24027_);
  and (_19900_, _16690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_10789_, _19900_, _19898_);
  and (_19901_, _16682_, _24053_);
  and (_19902_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or (_10791_, _19902_, _19901_);
  and (_19903_, _25226_, _24341_);
  nand (_19904_, _19903_, _23681_);
  or (_19905_, _19903_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_19906_, _19905_, _24330_);
  and (_19907_, _19906_, _19904_);
  nand (_19908_, _25236_, _23976_);
  or (_19909_, _25236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_19910_, _19909_, _22915_);
  and (_19911_, _19910_, _19908_);
  and (_19912_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_19913_, _19912_, rst);
  or (_19914_, _19913_, _19911_);
  or (_10794_, _19914_, _19907_);
  and (_19915_, _16682_, _23751_);
  and (_19916_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or (_10798_, _19916_, _19915_);
  and (_19917_, _16682_, _23715_);
  and (_19918_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or (_10800_, _19918_, _19917_);
  and (_19919_, _16682_, _23920_);
  and (_19920_, _16684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or (_10804_, _19920_, _19919_);
  and (_19921_, _25316_, _24341_);
  nand (_19922_, _19921_, _23681_);
  or (_19923_, _19921_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_19924_, _19923_, _24330_);
  and (_19925_, _19924_, _19922_);
  nand (_19926_, _25321_, _23976_);
  or (_19927_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_19928_, _19927_, _22915_);
  and (_19929_, _19928_, _19926_);
  and (_19930_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_19931_, _19930_, rst);
  or (_19932_, _19931_, _19929_);
  or (_10806_, _19932_, _19925_);
  and (_19934_, _02248_, _23715_);
  and (_19935_, _02250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or (_10810_, _19935_, _19934_);
  and (_19936_, _16632_, _23715_);
  and (_19937_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_26894_, _19937_, _19936_);
  and (_19938_, _09570_, _23693_);
  and (_19939_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_27052_, _19939_, _19938_);
  and (_19940_, _25315_, _24328_);
  and (_19941_, _19940_, _24341_);
  nand (_19942_, _19941_, _23681_);
  or (_19943_, _19941_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_19944_, _19943_, _24330_);
  and (_19945_, _19944_, _19942_);
  and (_19946_, _25235_, _24340_);
  nand (_19947_, _19946_, _23976_);
  or (_19948_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_19949_, _19948_, _22915_);
  and (_19950_, _19949_, _19947_);
  and (_19951_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_19952_, _19951_, rst);
  or (_19953_, _19952_, _19950_);
  or (_10816_, _19953_, _19945_);
  and (_19954_, _25225_, _24328_);
  and (_19955_, _19954_, _24341_);
  nand (_19956_, _19955_, _23681_);
  or (_19957_, _19955_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_19958_, _19957_, _24330_);
  and (_19959_, _19958_, _19956_);
  and (_19960_, _25235_, _24404_);
  nand (_19961_, _19960_, _23976_);
  or (_19962_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_19963_, _19962_, _22915_);
  and (_19964_, _19963_, _19961_);
  and (_19965_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_19966_, _19965_, rst);
  or (_19967_, _19966_, _19964_);
  or (_10818_, _19967_, _19959_);
  and (_19968_, _16992_, _23920_);
  and (_19969_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or (_27233_, _19969_, _19968_);
  and (_19970_, _16992_, _23900_);
  and (_19971_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or (_27232_, _19971_, _19970_);
  and (_19972_, _09570_, _23751_);
  and (_19973_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_27051_, _19973_, _19972_);
  and (_19974_, _02337_, _23715_);
  and (_19975_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_27036_, _19975_, _19974_);
  and (_19976_, _15246_, _23920_);
  and (_19977_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_10832_, _19977_, _19976_);
  and (_19978_, _25169_, _24053_);
  and (_19979_, _25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_10835_, _19979_, _19978_);
  nand (_19980_, _23357_, _23252_);
  not (_19981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_19982_, _24286_, _19981_);
  nor (_19983_, _10218_, _19981_);
  and (_19984_, _10218_, _19981_);
  or (_19985_, _19984_, _19983_);
  and (_19986_, _19985_, _24286_);
  nand (_19987_, _24294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_19988_, _19987_, _23210_);
  or (_19989_, _19988_, _19986_);
  or (_19990_, _19989_, _19982_);
  or (_19991_, _19990_, _23252_);
  and (_19992_, _19991_, _22773_);
  and (_10839_, _19992_, _19980_);
  and (_19993_, _24069_, _23715_);
  and (_19994_, _24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or (_10845_, _19994_, _19993_);
  and (_19995_, _02337_, _23693_);
  and (_19996_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_10855_, _19996_, _19995_);
  and (_19997_, _16992_, _23983_);
  and (_19998_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or (_10858_, _19998_, _19997_);
  and (_19999_, _09570_, _23920_);
  and (_20000_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_10861_, _20000_, _19999_);
  and (_20001_, _16094_, _24027_);
  and (_20002_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or (_10863_, _20002_, _20001_);
  and (_20003_, _15246_, _24027_);
  and (_20004_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_10867_, _20004_, _20003_);
  and (_20005_, _16094_, _23920_);
  and (_20006_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or (_10870_, _20006_, _20005_);
  and (_20007_, _04767_, _23900_);
  and (_20008_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_10873_, _20008_, _20007_);
  and (_20009_, _09570_, _23900_);
  and (_20010_, _09574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_10875_, _20010_, _20009_);
  and (_20011_, _09507_, _23900_);
  and (_20012_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_27202_, _20012_, _20011_);
  and (_20013_, _02789_, _23715_);
  and (_20014_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_27130_, _20014_, _20013_);
  and (_20015_, _24137_, _23751_);
  and (_20016_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_10878_, _20016_, _20015_);
  and (_20017_, _16632_, _23900_);
  and (_20018_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_10885_, _20018_, _20017_);
  and (_20020_, _24109_, _23751_);
  and (_20021_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_10890_, _20021_, _20020_);
  and (_20022_, _16632_, _24027_);
  and (_20023_, _16634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_10893_, _20023_, _20022_);
  and (_20024_, _24126_, _23920_);
  and (_20025_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_10895_, _20025_, _20024_);
  and (_20026_, _24131_, _24053_);
  and (_20027_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_10898_, _20027_, _20026_);
  and (_20028_, _16611_, _23693_);
  and (_20029_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or (_26896_, _20029_, _20028_);
  and (_20030_, _24126_, _23900_);
  and (_20031_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_10903_, _20031_, _20030_);
  and (_20032_, _24131_, _23751_);
  and (_20033_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_27315_, _20033_, _20032_);
  and (_20034_, _24126_, _24027_);
  and (_20035_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_27295_, _20035_, _20034_);
  and (_20036_, _02789_, _23693_);
  and (_20037_, _02791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_10912_, _20037_, _20036_);
  and (_20038_, _24109_, _23900_);
  and (_20039_, _24111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_10917_, _20039_, _20038_);
  nor (_26858_[6], _26107_, rst);
  and (_20040_, _24137_, _23900_);
  and (_20041_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_10925_, _20041_, _20040_);
  and (_20042_, _24137_, _24027_);
  and (_20043_, _24139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_10927_, _20043_, _20042_);
  and (_20044_, _24215_, _24053_);
  and (_20045_, _24217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or (_10929_, _20045_, _20044_);
  and (_20046_, _16611_, _23715_);
  and (_20047_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or (_26897_, _20047_, _20046_);
  and (_20048_, _24219_, _23693_);
  and (_20049_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or (_10935_, _20049_, _20048_);
  and (_20050_, _16611_, _23920_);
  and (_20051_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or (_26898_, _20051_, _20050_);
  and (_20052_, _24131_, _23900_);
  and (_20053_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_10938_, _20053_, _20052_);
  and (_20054_, _24131_, _24027_);
  and (_20055_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_27316_, _20055_, _20054_);
  and (_20056_, _16611_, _24027_);
  and (_20057_, _16613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or (_10941_, _20057_, _20056_);
  and (_20058_, _24117_, _23693_);
  and (_20059_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_10944_, _20059_, _20058_);
  and (_20060_, _24219_, _24053_);
  and (_20061_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or (_10947_, _20061_, _20060_);
  and (_20062_, _24250_, _23751_);
  and (_20063_, _24252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_10949_, _20063_, _20062_);
  and (_20064_, _24131_, _23715_);
  and (_20065_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_10951_, _20065_, _20064_);
  and (_20066_, _24117_, _24027_);
  and (_20067_, _24119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_10954_, _20067_, _20066_);
  and (_20068_, _24131_, _23920_);
  and (_20069_, _24133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_10956_, _20069_, _20068_);
  and (_20070_, _16595_, _23751_);
  and (_20071_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or (_10960_, _20071_, _20070_);
  and (_20072_, _16992_, _24053_);
  and (_20073_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or (_27231_, _20073_, _20072_);
  and (_20074_, _24219_, _23751_);
  and (_20075_, _24221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or (_27296_, _20075_, _20074_);
  and (_20076_, _16595_, _23715_);
  and (_20077_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or (_10968_, _20077_, _20076_);
  and (_20078_, _16094_, _23983_);
  and (_20079_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or (_10971_, _20079_, _20078_);
  and (_20080_, _24242_, _23715_);
  and (_20081_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or (_10979_, _20081_, _20080_);
  and (_20082_, _24242_, _23920_);
  and (_20083_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or (_10981_, _20083_, _20082_);
  and (_20084_, _16595_, _23900_);
  and (_20085_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or (_10983_, _20085_, _20084_);
  and (_20086_, _16595_, _23983_);
  and (_20087_, _16597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_10988_, _20087_, _20086_);
  and (_20088_, _24397_, _23920_);
  and (_20089_, _24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_10991_, _20089_, _20088_);
  and (_20090_, _24752_, _23900_);
  and (_20091_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_10993_, _20091_, _20090_);
  and (_20092_, _24126_, _23751_);
  and (_20093_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_27294_, _20093_, _20092_);
  and (_20094_, _02794_, _23715_);
  and (_20095_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or (_10998_, _20095_, _20094_);
  and (_20096_, _24126_, _23715_);
  and (_20097_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_11000_, _20097_, _20096_);
  and (_20098_, _16589_, _24053_);
  and (_20099_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_11002_, _20099_, _20098_);
  and (_20100_, _16998_, _23983_);
  and (_20101_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_11004_, _20101_, _20100_);
  and (_20102_, _24231_, _23715_);
  and (_20103_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or (_11007_, _20103_, _20102_);
  and (_20104_, _16589_, _23693_);
  and (_20105_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_11009_, _20105_, _20104_);
  and (_20106_, _24231_, _23920_);
  and (_20107_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or (_11011_, _20107_, _20106_);
  and (_20108_, _24231_, _24027_);
  and (_20109_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or (_11014_, _20109_, _20108_);
  and (_20110_, _02794_, _23693_);
  and (_20111_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or (_27129_, _20111_, _20110_);
  and (_20112_, _24158_, _23751_);
  and (_20113_, _24160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_27267_, _20113_, _20112_);
  and (_20114_, _24126_, _23693_);
  and (_20115_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_11018_, _20115_, _20114_);
  and (_20116_, _24752_, _23983_);
  and (_20117_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or (_11020_, _20117_, _20116_);
  and (_20118_, _02794_, _23751_);
  and (_20119_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or (_11022_, _20119_, _20118_);
  and (_20120_, _16589_, _23715_);
  and (_20121_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_11024_, _20121_, _20120_);
  and (_20122_, _24231_, _23693_);
  and (_20123_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or (_11028_, _20123_, _20122_);
  and (_20124_, _17147_, _23983_);
  and (_20125_, _17149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_11030_, _20125_, _20124_);
  and (_20126_, _16589_, _23983_);
  and (_20127_, _16591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_11032_, _20127_, _20126_);
  and (_20128_, _24231_, _23900_);
  and (_20129_, _24233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or (_11036_, _20129_, _20128_);
  and (_20130_, _24752_, _23715_);
  and (_20131_, _24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or (_27265_, _20131_, _20130_);
  and (_20132_, _24126_, _24053_);
  and (_20133_, _24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_11039_, _20133_, _20132_);
  and (_20134_, _16231_, _23983_);
  and (_20135_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_11043_, _20135_, _20134_);
  and (_20136_, _16577_, _24053_);
  and (_20137_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_11045_, _20137_, _20136_);
  and (_20138_, _24242_, _24053_);
  and (_20139_, _24244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or (_11058_, _20139_, _20138_);
  and (_20140_, _24305_, _23900_);
  and (_20141_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or (_11061_, _20141_, _20140_);
  and (_20142_, _16231_, _24027_);
  and (_20143_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_11065_, _20143_, _20142_);
  and (_20144_, _04033_, _23900_);
  and (_20145_, _04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or (_11076_, _20145_, _20144_);
  and (_20146_, _24389_, _23693_);
  and (_20147_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_11078_, _20147_, _20146_);
  and (_20148_, _24389_, _24053_);
  and (_20149_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_27185_, _20149_, _20148_);
  and (_20150_, _25454_, _23983_);
  and (_20151_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or (_27184_, _20151_, _20150_);
  and (_20152_, _16577_, _23693_);
  and (_20153_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_11086_, _20153_, _20152_);
  and (_20154_, _25454_, _23715_);
  and (_20155_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or (_11088_, _20155_, _20154_);
  and (_20156_, _25454_, _23751_);
  and (_20157_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or (_11090_, _20157_, _20156_);
  and (_20158_, _25436_, _23920_);
  and (_20159_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or (_11095_, _20159_, _20158_);
  and (_20160_, _16577_, _23715_);
  and (_20161_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_11097_, _20161_, _20160_);
  and (_20162_, _16094_, _23715_);
  and (_20163_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or (_11099_, _20163_, _20162_);
  and (_20164_, _25436_, _24053_);
  and (_20165_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or (_11103_, _20165_, _20164_);
  and (_20166_, _25402_, _24027_);
  and (_20167_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_11107_, _20167_, _20166_);
  and (_20168_, _02423_, _24027_);
  and (_20169_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or (_11109_, _20169_, _20168_);
  and (_20170_, _16577_, _24027_);
  and (_20171_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_11111_, _20171_, _20170_);
  and (_20172_, _25402_, _23751_);
  and (_20173_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_11113_, _20173_, _20172_);
  and (_20174_, _25389_, _24027_);
  and (_20175_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_27168_, _20175_, _20174_);
  and (_20176_, _16577_, _23983_);
  and (_20177_, _16579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_26901_, _20177_, _20176_);
  and (_20178_, _25389_, _23751_);
  and (_20179_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_27167_, _20179_, _20178_);
  and (_20180_, _25356_, _23983_);
  and (_20181_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or (_11121_, _20181_, _20180_);
  and (_20182_, _24305_, _23715_);
  and (_20183_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or (_11124_, _20183_, _20182_);
  and (_20184_, _16094_, _23693_);
  and (_20185_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or (_11126_, _20185_, _20184_);
  and (_20186_, _02794_, _23920_);
  and (_20187_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or (_11130_, _20187_, _20186_);
  and (_20188_, _25356_, _23693_);
  and (_20189_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or (_11132_, _20189_, _20188_);
  and (_20190_, _25346_, _24027_);
  and (_20191_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or (_11134_, _20191_, _20190_);
  and (_20192_, _16094_, _23751_);
  and (_20193_, _16096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or (_11136_, _20193_, _20192_);
  and (_20194_, _25346_, _23900_);
  and (_20195_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or (_11138_, _20195_, _20194_);
  and (_20196_, _25346_, _24053_);
  and (_20197_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or (_11141_, _20197_, _20196_);
  and (_20198_, _25194_, _23983_);
  and (_20199_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_27157_, _20199_, _20198_);
  and (_20201_, _25194_, _23920_);
  and (_20202_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_11145_, _20202_, _20201_);
  and (_20203_, _24305_, _23693_);
  and (_20204_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or (_27048_, _20204_, _20203_);
  and (_20205_, _25220_, _23920_);
  and (_20206_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_11149_, _20206_, _20205_);
  and (_20207_, _25220_, _24053_);
  and (_20208_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_11154_, _20208_, _20207_);
  and (_20209_, _25210_, _24027_);
  and (_20210_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_11156_, _20210_, _20209_);
  and (_20211_, _02794_, _23900_);
  and (_20212_, _02796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or (_11159_, _20212_, _20211_);
  and (_20213_, _25198_, _24027_);
  and (_20214_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or (_11163_, _20214_, _20213_);
  and (_20215_, _25198_, _23900_);
  and (_20216_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or (_11166_, _20216_, _20215_);
  and (_20217_, _16472_, _23751_);
  and (_20218_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or (_26902_, _20218_, _20217_);
  and (_20219_, _25194_, _23751_);
  and (_20220_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_11170_, _20220_, _20219_);
  and (_20221_, _16992_, _23693_);
  and (_20222_, _16994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or (_11173_, _20222_, _20221_);
  and (_20223_, _25180_, _23920_);
  and (_20224_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or (_11176_, _20224_, _20223_);
  and (_20225_, _16472_, _23715_);
  and (_20226_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or (_11178_, _20226_, _20225_);
  and (_20228_, _25454_, _23920_);
  and (_20229_, _25456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or (_27182_, _20229_, _20228_);
  nor (_20230_, _24192_, rst);
  not (_20231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_20232_, _24984_, _20231_);
  or (_20233_, _20232_, _24993_);
  and (_20234_, _20233_, _24975_);
  or (_20235_, _24206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_20236_, _20235_, _25012_);
  or (_20237_, _20236_, _20232_);
  and (_20238_, _20237_, _24976_);
  nor (_20239_, _20238_, _20234_);
  nor (_20240_, _20239_, _24186_);
  and (_11183_, _20240_, _20230_);
  and (_20241_, _16472_, _23900_);
  and (_20242_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or (_11187_, _20242_, _20241_);
  and (_20243_, _25436_, _23693_);
  and (_20244_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or (_11190_, _20244_, _20243_);
  and (_20245_, _25402_, _23715_);
  and (_20246_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_11192_, _20246_, _20245_);
  and (_20247_, _25389_, _23715_);
  and (_20248_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_11194_, _20248_, _20247_);
  and (_20249_, _16231_, _24053_);
  and (_20250_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_11197_, _20250_, _20249_);
  nand (_20251_, _26622_, _26607_);
  or (_20252_, _26607_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_20253_, _20252_, _22773_);
  and (_11199_, _20253_, _20251_);
  and (_20254_, _25356_, _23900_);
  and (_20255_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or (_27166_, _20255_, _20254_);
  and (_20256_, _16472_, _23920_);
  and (_20257_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or (_26903_, _20257_, _20256_);
  and (_20258_, _16472_, _23983_);
  and (_20259_, _16474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or (_26904_, _20259_, _20258_);
  and (_20260_, _15255_, _24053_);
  and (_20261_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or (_26905_, _20261_, _20260_);
  and (_20262_, _25180_, _23751_);
  and (_20263_, _25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or (_27136_, _20263_, _20262_);
  and (_20264_, _25220_, _23693_);
  and (_20265_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_27120_, _20265_, _20264_);
  and (_20266_, _25210_, _23715_);
  and (_20267_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_27106_, _20267_, _20266_);
  and (_20268_, _17099_, _24053_);
  and (_20269_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_27213_, _20269_, _20268_);
  and (_20270_, _15255_, _23751_);
  and (_20271_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or (_26906_, _20271_, _20270_);
  and (_20272_, _15255_, _23715_);
  and (_20273_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or (_26908_, _20273_, _20272_);
  and (_20274_, _16231_, _23751_);
  and (_20275_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_26925_, _20275_, _20274_);
  and (_20276_, _24389_, _23900_);
  and (_20277_, _24391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_27188_, _20277_, _20276_);
  and (_20278_, _15255_, _23900_);
  and (_20279_, _15257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or (_26909_, _20279_, _20278_);
  and (_20280_, _25436_, _24027_);
  and (_20281_, _25438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or (_27175_, _20281_, _20280_);
  and (_20282_, _25402_, _23983_);
  and (_20283_, _25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_27171_, _20283_, _20282_);
  and (_20284_, _25389_, _23983_);
  and (_20285_, _25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_27169_, _20285_, _20284_);
  and (_20286_, _25356_, _24053_);
  and (_20287_, _25358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or (_27164_, _20287_, _20286_);
  and (_20288_, _25346_, _23751_);
  and (_20289_, _25348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or (_27162_, _20289_, _20288_);
  and (_20290_, _25220_, _24027_);
  and (_20291_, _25222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_27121_, _20291_, _20290_);
  and (_20292_, _25210_, _23983_);
  and (_20293_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_27109_, _20293_, _20292_);
  and (_20294_, _25210_, _24053_);
  and (_20295_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_27105_, _20295_, _20294_);
  and (_20296_, _25194_, _23693_);
  and (_20297_, _25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_27156_, _20297_, _20296_);
  and (_20298_, _06253_, _23900_);
  and (_20299_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or (_27128_, _20299_, _20298_);
  and (_20300_, _17059_, _23920_);
  and (_20301_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_27257_, _20301_, _20300_);
  and (_20302_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_27319_, _20302_, _02986_);
  and (_20303_, _01876_, _23751_);
  and (_20304_, _01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_27301_, _20304_, _20303_);
  and (_20305_, _02203_, _23900_);
  and (_20306_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_27285_, _20306_, _20305_);
  and (_20307_, _17059_, _23900_);
  and (_20308_, _17061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_27256_, _20308_, _20307_);
  and (_20309_, _02392_, _23983_);
  and (_20310_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_27239_, _20310_, _20309_);
  and (_20311_, _02392_, _24053_);
  and (_20312_, _02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_27236_, _20312_, _20311_);
  and (_20313_, _02427_, _23715_);
  and (_20314_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_27221_, _20314_, _20313_);
  and (_20315_, _02503_, _24027_);
  and (_20316_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_27203_, _20316_, _20315_);
  and (_20317_, _06253_, _23715_);
  and (_20318_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or (_27127_, _20318_, _20317_);
  and (_20319_, _06253_, _23693_);
  and (_20320_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or (_27126_, _20320_, _20319_);
  and (_20321_, _25165_, _23900_);
  and (_20322_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_26936_, _20322_, _20321_);
  and (_26878_, _01717_, _22773_);
  and (_20323_, _26871_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_26877_, _20323_, _26878_);
  and (_20324_, _02344_, _24027_);
  and (_20325_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_27263_, _20325_, _20324_);
  and (_20326_, _02650_, _23715_);
  and (_20327_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_27177_, _20327_, _20326_);
  and (_20328_, _02681_, _23751_);
  and (_20329_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_27061_, _20329_, _20328_);
  nand (_20330_, _23756_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_26876_, _20330_, _22773_);
  and (_20331_, _01952_, _23983_);
  and (_20332_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_11324_, _20332_, _20331_);
  and (_20333_, _01860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_27320_, _20333_, _02571_);
  and (_20334_, _24238_, _23751_);
  and (_20335_, _24240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or (_11331_, _20335_, _20334_);
  and (_20336_, _02503_, _23983_);
  and (_20337_, _02505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_27204_, _20337_, _20336_);
  and (_20338_, _16231_, _23900_);
  and (_20339_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_11336_, _20339_, _20338_);
  or (_20340_, _24840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_20341_, _24853_, _24859_);
  nand (_20342_, _20341_, _20340_);
  nand (_20343_, _20342_, _24879_);
  nor (_20344_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _24859_);
  or (_20345_, _24870_, _24864_);
  nor (_20346_, _20345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_20347_, _20346_, _20344_);
  and (_20348_, _20347_, _20343_);
  or (_20349_, _20348_, _24855_);
  or (_20350_, _24922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_20351_, _20350_, _22773_);
  and (_11355_, _20351_, _20349_);
  and (_20352_, _24919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_20353_, _24859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_20354_, _24859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_20355_, _20354_, _20353_);
  nor (_20356_, _20355_, _24879_);
  or (_20357_, _20356_, _24855_);
  or (_20358_, _20357_, _20352_);
  or (_20359_, _20355_, _24922_);
  and (_20360_, _20359_, _22773_);
  and (_11357_, _20360_, _20358_);
  and (_11359_, _00584_, _22773_);
  and (_20361_, _16231_, _23715_);
  and (_20362_, _16233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_11363_, _20362_, _20361_);
  or (_20363_, _24840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nand (_20364_, _24853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_20365_, _20364_, _20363_);
  nand (_20366_, _20365_, _24879_);
  nor (_20367_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_20368_, _20367_);
  or (_20369_, _20345_, _24859_);
  and (_20370_, _20369_, _20368_);
  and (_20371_, _20370_, _20366_);
  or (_20372_, _20371_, _24855_);
  or (_20373_, _24922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_20374_, _20373_, _22773_);
  and (_11365_, _20374_, _20372_);
  and (_20375_, _06253_, _24027_);
  and (_20376_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or (_11373_, _20376_, _20375_);
  and (_20377_, _02344_, _23983_);
  and (_20378_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_27264_, _20378_, _20377_);
  and (_20379_, _23721_, _23715_);
  and (_20380_, _23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_27027_, _20380_, _20379_);
  and (_20381_, _02681_, _23693_);
  and (_20382_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_11389_, _20382_, _20381_);
  and (_20383_, _06253_, _23983_);
  and (_20384_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or (_11404_, _20384_, _20383_);
  and (_20385_, _25482_, _24027_);
  and (_20386_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_11406_, _20386_, _20385_);
  nor (_20387_, _25055_, _24928_);
  nor (_20388_, _20387_, _24822_);
  and (_20389_, _20388_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor (_20390_, _01812_, _01783_);
  nor (_20391_, _20390_, _24822_);
  nor (_20392_, _20344_, _24822_);
  and (_20393_, _20392_, _20368_);
  nor (_20394_, _20393_, _20391_);
  nand (_20395_, _20394_, _20389_);
  nand (_20396_, _20395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_20397_, _20396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_20398_, _22857_, _22927_);
  nor (_20399_, _24420_, _20398_);
  or (_20400_, _20399_, _20397_);
  nand (_20401_, _20399_, _23708_);
  and (_20402_, _20401_, _20400_);
  nand (_20403_, _20402_, _24764_);
  or (_20404_, _24764_, _23744_);
  and (_20405_, _20404_, _22773_);
  and (_11415_, _20405_, _20403_);
  and (_20406_, _12702_, _24053_);
  and (_20407_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or (_11417_, _20407_, _20406_);
  not (_20408_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_20409_, _20388_, _20408_);
  nand (_20410_, _20393_, _20390_);
  or (_20411_, _20410_, _20409_);
  and (_20412_, _20411_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_20413_, _20412_, _04173_);
  and (_20414_, _24421_, _22857_);
  and (_20415_, _20414_, _24341_);
  or (_20416_, _20415_, _20413_);
  nand (_20417_, _20415_, _23681_);
  and (_20418_, _20417_, _20416_);
  or (_20419_, _20418_, _24763_);
  nand (_20420_, _24763_, _23976_);
  and (_20421_, _20420_, _22773_);
  and (_11423_, _20421_, _20419_);
  and (_20422_, _20414_, _23250_);
  and (_20423_, _20422_, _23708_);
  nand (_20424_, _02562_, _22928_);
  nand (_20425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  not (_20426_, _20393_);
  and (_20427_, _20426_, _20391_);
  and (_20428_, _20427_, _20389_);
  or (_20429_, _20428_, _20425_);
  or (_20430_, _20429_, _20422_);
  nand (_20431_, _20430_, _20424_);
  or (_20432_, _20431_, _20423_);
  or (_20433_, _24764_, _23413_);
  and (_20434_, _20433_, _22773_);
  and (_11430_, _20434_, _20432_);
  nor (_20435_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _20231_);
  not (_20436_, _20427_);
  or (_20437_, _20436_, _20409_);
  and (_20438_, _20437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_20439_, _20438_, _20435_);
  and (_20440_, _20414_, _23208_);
  or (_20441_, _20440_, _20439_);
  nand (_20442_, _20440_, _23681_);
  and (_20443_, _20442_, _20441_);
  or (_20444_, _20443_, _24763_);
  nand (_20445_, _24763_, _23357_);
  and (_20446_, _20445_, _22773_);
  and (_11440_, _20446_, _20444_);
  and (_20447_, _24341_, _24333_);
  nand (_20448_, _20447_, _23681_);
  or (_20449_, _20447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_20450_, _20449_, _24347_);
  and (_20451_, _20450_, _20448_);
  nor (_20452_, _24347_, _23976_);
  or (_20453_, _20452_, _20451_);
  and (_11444_, _20453_, _22773_);
  and (_20454_, _23763_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_20455_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_20456_, _23763_, _20455_);
  or (_20457_, _20456_, _20454_);
  and (_26853_[15], _20457_, _22773_);
  and (_20458_, _24411_, _24341_);
  or (_20459_, _20458_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_20460_, _20459_, _24417_);
  nand (_20461_, _20458_, _23681_);
  and (_20462_, _20461_, _20460_);
  nor (_20463_, _24417_, _23976_);
  or (_20464_, _20463_, _20462_);
  and (_11450_, _20464_, _22773_);
  and (_11453_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _22773_);
  and (_20465_, _24759_, _24373_);
  or (_20466_, _20465_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_20467_, _20466_, _24764_);
  nand (_20468_, _20465_, _23681_);
  and (_20469_, _20468_, _20467_);
  nor (_20470_, _24764_, _24017_);
  or (_20471_, _20470_, _20469_);
  and (_11456_, _20471_, _22773_);
  and (_20472_, _23268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_20473_, _20472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_20474_, _20473_, _19640_);
  and (_20475_, _20474_, _10189_);
  and (_20476_, _10191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_20477_, _24294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_20478_, _20477_, _23210_);
  or (_20479_, _20478_, _20476_);
  or (_20480_, _20479_, _20475_);
  and (_20481_, _20480_, _23253_);
  and (_20482_, _23744_, _23252_);
  or (_20483_, _20482_, _20481_);
  and (_11459_, _20483_, _22773_);
  nand (_20484_, _24919_, _24822_);
  nand (_20485_, _20353_, _24855_);
  and (_20486_, _20485_, _22773_);
  and (_11462_, _20486_, _20484_);
  and (_20487_, _15238_, _23983_);
  and (_20488_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_11469_, _20488_, _20487_);
  and (_20489_, _02423_, _23920_);
  and (_20490_, _02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or (_11472_, _20490_, _20489_);
  and (_20491_, _02326_, _23715_);
  and (_20492_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or (_11480_, _20492_, _20491_);
  and (_20493_, _02337_, _24027_);
  and (_20494_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_11492_, _20494_, _20493_);
  and (_20495_, _02337_, _23920_);
  and (_20496_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_11497_, _20496_, _20495_);
  and (_20497_, _17099_, _23693_);
  and (_20498_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_11500_, _20498_, _20497_);
  and (_20499_, _02337_, _23900_);
  and (_20500_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_11522_, _20500_, _20499_);
  and (_20501_, _17099_, _23751_);
  and (_20502_, _17101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_11538_, _20502_, _20501_);
  and (_20503_, _09507_, _23715_);
  and (_20504_, _09509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_11541_, _20504_, _20503_);
  and (_20505_, _19940_, _24184_);
  nand (_20506_, _20505_, _23681_);
  or (_20507_, _20505_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_20508_, _20507_, _24330_);
  and (_20509_, _20508_, _20506_);
  not (_20510_, _19946_);
  or (_20511_, _20510_, _23247_);
  or (_20512_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_20513_, _20512_, _22915_);
  and (_20514_, _20513_, _20511_);
  and (_20515_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_20516_, _20515_, rst);
  or (_20517_, _20516_, _20514_);
  or (_11552_, _20517_, _20509_);
  and (_20518_, _19940_, _23208_);
  nand (_20519_, _20518_, _23681_);
  or (_20520_, _20518_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_20521_, _20520_, _24330_);
  and (_20522_, _20521_, _20519_);
  nand (_20523_, _19946_, _23357_);
  or (_20524_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_20525_, _20524_, _22915_);
  and (_20526_, _20525_, _20523_);
  nor (_20527_, _22914_, _03640_);
  or (_20528_, _20527_, rst);
  or (_20529_, _20528_, _20526_);
  or (_11554_, _20529_, _20522_);
  and (_20530_, _08435_, _23693_);
  and (_20531_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or (_11566_, _20531_, _20530_);
  and (_20532_, _25176_, _23900_);
  and (_20533_, _25178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or (_11570_, _20533_, _20532_);
  and (_20534_, _12702_, _23751_);
  and (_20535_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or (_11572_, _20535_, _20534_);
  and (_20536_, _19940_, _23250_);
  nand (_20537_, _20536_, _23681_);
  or (_20538_, _20536_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_20539_, _20538_, _24330_);
  and (_20540_, _20539_, _20537_);
  or (_20541_, _20510_, _23413_);
  or (_20542_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_20543_, _20542_, _22915_);
  and (_20544_, _20543_, _20541_);
  nor (_20545_, _22914_, _03627_);
  or (_20546_, _20545_, rst);
  or (_20547_, _20546_, _20544_);
  or (_11591_, _20547_, _20540_);
  and (_20548_, _19940_, _24373_);
  nand (_20549_, _20548_, _23681_);
  or (_20550_, _20548_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_20551_, _20550_, _24330_);
  and (_20552_, _20551_, _20549_);
  nand (_20553_, _19946_, _24017_);
  or (_20554_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_20555_, _20554_, _22915_);
  and (_20556_, _20555_, _20553_);
  and (_20557_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_20558_, _20557_, rst);
  or (_20559_, _20558_, _20556_);
  or (_11605_, _20559_, _20552_);
  and (_20560_, _19940_, _22895_);
  nand (_20561_, _20560_, _23681_);
  or (_20562_, _20560_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_20563_, _20562_, _24330_);
  and (_20564_, _20563_, _20561_);
  or (_20565_, _20510_, _23744_);
  or (_20566_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_20567_, _20566_, _22915_);
  and (_20568_, _20567_, _20565_);
  nor (_20569_, _22914_, _03645_);
  or (_20570_, _20569_, rst);
  or (_20571_, _20570_, _20568_);
  or (_11607_, _20571_, _20564_);
  and (_20572_, _19940_, _24405_);
  nand (_20573_, _20572_, _23681_);
  or (_20574_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_20575_, _20574_, _24330_);
  and (_20576_, _20575_, _20573_);
  nand (_20577_, _19946_, _24047_);
  and (_20578_, _20574_, _22915_);
  and (_20579_, _20578_, _20577_);
  nor (_20580_, _22914_, _03620_);
  or (_20581_, _20580_, rst);
  or (_20582_, _20581_, _20579_);
  or (_11609_, _20582_, _20576_);
  and (_20583_, _12702_, _23693_);
  and (_20584_, _12704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or (_11611_, _20584_, _20583_);
  and (_20585_, _02798_, _23983_);
  and (_20586_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_11617_, _20586_, _20585_);
  or (_20587_, _02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_11619_, _20587_, _02882_);
  and (_20588_, _02681_, _24053_);
  and (_20589_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_11621_, _20589_, _20588_);
  and (_20590_, _02681_, _23983_);
  and (_20591_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_11633_, _20591_, _20590_);
  and (_20592_, _02681_, _23920_);
  and (_20593_, _02683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_11637_, _20593_, _20592_);
  and (_11639_, _00737_, _22773_);
  and (_11641_, _00794_, _22773_);
  and (_11643_, _00999_, _22773_);
  and (_11645_, _01081_, _22773_);
  and (_11647_, _26777_, _22773_);
  and (_11649_, _00072_, _22773_);
  and (_20594_, _02650_, _23693_);
  and (_20595_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_11651_, _20595_, _20594_);
  and (_11653_, _00332_, _22773_);
  and (_11655_, _00412_, _22773_);
  and (_20596_, _02650_, _24027_);
  and (_20597_, _02652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_11657_, _20597_, _20596_);
  and (_11659_, _00681_, _22773_);
  and (_11661_, _00857_, _22773_);
  and (_11663_, _03285_, _22773_);
  and (_11665_, _00155_, _22773_);
  and (_20598_, _17069_, _23920_);
  and (_20599_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_11667_, _20599_, _20598_);
  and (_11670_, _00932_, _22773_);
  and (_11674_, _00250_, _22773_);
  and (_20600_, _02427_, _24053_);
  and (_20601_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_11678_, _20601_, _20600_);
  and (_20602_, _17069_, _23900_);
  and (_20603_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_11680_, _20603_, _20602_);
  and (_20604_, _15238_, _23715_);
  and (_20605_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_11685_, _20605_, _20604_);
  and (_20606_, _02344_, _23920_);
  and (_20607_, _02346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_11689_, _20607_, _20606_);
  and (_20608_, _02203_, _23983_);
  and (_20609_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_11692_, _20609_, _20608_);
  nor (_20610_, _26607_, _26617_);
  and (_20611_, _26607_, _26617_);
  or (_20612_, _20611_, _20610_);
  and (_11716_, _20612_, _22773_);
  and (_20613_, _08435_, _23751_);
  and (_20614_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or (_11721_, _20614_, _20613_);
  and (_20615_, _01541_, _23900_);
  and (_20616_, _01543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_26900_, _20616_, _20615_);
  and (_20617_, _15238_, _23693_);
  and (_20618_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_11724_, _20618_, _20617_);
  and (_20619_, _25503_, _23983_);
  and (_20620_, _25505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_11727_, _20620_, _20619_);
  and (_20621_, _25165_, _23751_);
  and (_20622_, _25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_11829_, _20622_, _20621_);
  nor (_26858_[4], _26004_, rst);
  and (_20623_, _15238_, _23751_);
  and (_20624_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_11833_, _20624_, _20623_);
  and (_20625_, _06253_, _24053_);
  and (_20626_, _06255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or (_11836_, _20626_, _20625_);
  and (_20627_, _24305_, _23983_);
  and (_20628_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or (_11842_, _20628_, _20627_);
  and (_20629_, _24305_, _24027_);
  and (_20630_, _24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or (_27050_, _20630_, _20629_);
  and (_20631_, _16998_, _23715_);
  and (_20632_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_11845_, _20632_, _20631_);
  and (_20633_, _23983_, _23707_);
  and (_20634_, _23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_26911_, _20634_, _20633_);
  and (_20635_, _16998_, _23693_);
  and (_20636_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_11849_, _20636_, _20635_);
  and (_20637_, _17069_, _23983_);
  and (_20638_, _17071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_11851_, _20638_, _20637_);
  and (_20639_, _15238_, _23920_);
  and (_20640_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_11853_, _20640_, _20639_);
  and (_20641_, _15238_, _23900_);
  and (_20642_, _15240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_11855_, _20642_, _20641_);
  and (_26832_[1], _25942_, _22773_);
  and (_20643_, _02829_, _23751_);
  and (_20644_, _02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or (_11861_, _20644_, _20643_);
  and (_20645_, _02798_, _23693_);
  and (_20646_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_11864_, _20646_, _20645_);
  and (_20647_, _01701_, _23751_);
  and (_20648_, _01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or (_11866_, _20648_, _20647_);
  and (_20649_, _16998_, _23920_);
  and (_20650_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_11868_, _20650_, _20649_);
  and (_20651_, _01952_, _23715_);
  and (_20652_, _01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or (_27212_, _20652_, _20651_);
  and (_20653_, _19940_, _24190_);
  nand (_20654_, _20653_, _23681_);
  or (_20655_, _20653_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_20656_, _20655_, _24330_);
  and (_20657_, _20656_, _20654_);
  or (_20658_, _20510_, _23205_);
  or (_20659_, _19946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_20660_, _20659_, _22915_);
  and (_20661_, _20660_, _20658_);
  nor (_20662_, _22914_, _03615_);
  or (_20663_, _20662_, rst);
  or (_20664_, _20663_, _20661_);
  or (_11872_, _20664_, _20657_);
  and (_20665_, _24268_, _23920_);
  and (_20666_, _24270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_27045_, _20666_, _20665_);
  and (_20667_, _16998_, _23900_);
  and (_20668_, _17001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_11875_, _20668_, _20667_);
  and (_20669_, _19954_, _24373_);
  nand (_20670_, _20669_, _23681_);
  or (_20671_, _20669_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_20672_, _20671_, _24330_);
  and (_20673_, _20672_, _20670_);
  nand (_20674_, _19960_, _24017_);
  or (_20675_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_20676_, _20675_, _22915_);
  and (_20677_, _20676_, _20674_);
  and (_20678_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_20679_, _20678_, rst);
  or (_20680_, _20679_, _20677_);
  or (_12076_, _20680_, _20673_);
  and (_20681_, _19954_, _23208_);
  nand (_20682_, _20681_, _23681_);
  or (_20683_, _20681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_20684_, _20683_, _24330_);
  and (_20685_, _20684_, _20682_);
  nand (_20686_, _19960_, _23357_);
  or (_20687_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_20688_, _20687_, _22915_);
  and (_20689_, _20688_, _20686_);
  nor (_20690_, _22914_, _03692_);
  or (_20691_, _20690_, rst);
  or (_20692_, _20691_, _20689_);
  or (_12078_, _20692_, _20685_);
  and (_20693_, _16219_, _23900_);
  and (_20694_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or (_12082_, _20694_, _20693_);
  and (_20695_, _19954_, _23250_);
  nand (_20696_, _20695_, _23681_);
  or (_20697_, _20695_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_20698_, _20697_, _24330_);
  and (_20699_, _20698_, _20696_);
  not (_20700_, _19960_);
  or (_20701_, _20700_, _23413_);
  or (_20702_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_20703_, _20702_, _22915_);
  and (_20704_, _20703_, _20701_);
  nor (_20705_, _22914_, _03679_);
  or (_20706_, _20705_, rst);
  or (_20707_, _20706_, _20704_);
  or (_12086_, _20707_, _20699_);
  and (_20708_, _19954_, _24184_);
  nand (_20709_, _20708_, _23681_);
  or (_20710_, _20708_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_20711_, _20710_, _24330_);
  and (_20712_, _20711_, _20709_);
  or (_20713_, _20700_, _23247_);
  or (_20714_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_20715_, _20714_, _22915_);
  and (_20716_, _20715_, _20713_);
  and (_20717_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_20718_, _20717_, rst);
  or (_20719_, _20718_, _20716_);
  or (_12088_, _20719_, _20712_);
  and (_20720_, _19954_, _22895_);
  nand (_20721_, _20720_, _23681_);
  or (_20722_, _20720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_20723_, _20722_, _24330_);
  and (_20724_, _20723_, _20721_);
  or (_20725_, _20700_, _23744_);
  or (_20726_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_20727_, _20726_, _22915_);
  and (_20728_, _20727_, _20725_);
  nor (_20729_, _22914_, _03698_);
  or (_20730_, _20729_, rst);
  or (_20731_, _20730_, _20728_);
  or (_12090_, _20731_, _20724_);
  and (_20732_, _19954_, _24405_);
  nand (_20733_, _20732_, _23681_);
  or (_20734_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_20735_, _20734_, _24330_);
  and (_20736_, _20735_, _20733_);
  nand (_20737_, _19960_, _24047_);
  and (_20738_, _20734_, _22915_);
  and (_20739_, _20738_, _20737_);
  nor (_20740_, _22914_, _03671_);
  or (_20741_, _20740_, rst);
  or (_20742_, _20741_, _20739_);
  or (_12092_, _20742_, _20736_);
  and (_20743_, _19954_, _24190_);
  nand (_20744_, _20743_, _23681_);
  or (_20745_, _20743_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_20746_, _20745_, _24330_);
  and (_20747_, _20746_, _20744_);
  or (_20748_, _20700_, _23205_);
  or (_20749_, _19960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_20750_, _20749_, _22915_);
  and (_20751_, _20750_, _20748_);
  nor (_20752_, _22914_, _03666_);
  or (_20753_, _20752_, rst);
  or (_20754_, _20753_, _20751_);
  or (_12094_, _20754_, _20747_);
  and (_20755_, _25316_, _24373_);
  nand (_20756_, _20755_, _23681_);
  or (_20757_, _20755_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_20758_, _20757_, _24330_);
  and (_20759_, _20758_, _20756_);
  nand (_20760_, _25321_, _24017_);
  or (_20761_, _25321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_20762_, _20761_, _22915_);
  and (_20763_, _20762_, _20760_);
  and (_20764_, _25257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_20765_, _20764_, rst);
  or (_20766_, _20765_, _20763_);
  or (_12105_, _20766_, _20759_);
  and (_20767_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20768_, _20767_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20769_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_20770_, _20769_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_20771_, _20770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_20772_, _20771_, _20768_);
  and (_20773_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_20774_, _20773_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_20775_, _20774_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_20776_, _20775_, _20772_);
  and (_20777_, _20776_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_20778_, _20777_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_20779_, _20778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20780_, _20778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20781_, _20780_, _20779_);
  nor (_20782_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20783_, _20782_);
  and (_20784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _23830_);
  and (_20785_, _20767_, _23844_);
  nor (_20786_, _20767_, _23844_);
  nor (_20787_, _20786_, _20785_);
  nor (_20788_, _20787_, _23830_);
  nor (_20789_, _20788_, _20784_);
  not (_20790_, _20789_);
  nor (_20791_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20792_, _23840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20793_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _23835_);
  nor (_20794_, _20793_, _20792_);
  and (_20795_, _20794_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20796_, _20795_, _20791_);
  nor (_20797_, _20796_, _05474_);
  and (_20798_, _20796_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_20799_, _20798_, _20797_);
  nor (_20800_, _20799_, _20790_);
  nor (_20801_, _20796_, _05024_);
  and (_20802_, _20796_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_20803_, _20802_, _20801_);
  nor (_20804_, _20803_, _20789_);
  nor (_20805_, _20804_, _20800_);
  nor (_20806_, _20805_, _20783_);
  and (_20807_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _23830_);
  not (_20808_, _20807_);
  nor (_20809_, _20796_, _05011_);
  and (_20810_, _20796_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_20811_, _20810_, _20809_);
  nor (_20812_, _20811_, _20790_);
  not (_20813_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_20814_, _20796_, _20813_);
  and (_20815_, _20796_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_20816_, _20815_, _20814_);
  nor (_20817_, _20816_, _20789_);
  nor (_20818_, _20817_, _20812_);
  nor (_20819_, _20818_, _20808_);
  nor (_20820_, _20819_, _20806_);
  and (_20821_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20822_, _20821_);
  nor (_20823_, _20796_, _05035_);
  and (_20824_, _20796_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_20825_, _20824_, _20823_);
  nor (_20826_, _20825_, _20790_);
  not (_20827_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_20828_, _20796_, _20827_);
  and (_20829_, _20796_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_20830_, _20829_, _20828_);
  nor (_20831_, _20830_, _20789_);
  nor (_20832_, _20831_, _20826_);
  nor (_20833_, _20832_, _20822_);
  and (_20834_, _23835_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20835_, _20834_);
  nor (_20836_, _20796_, _05054_);
  and (_20837_, _20796_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_20838_, _20837_, _20836_);
  nor (_20839_, _20838_, _20790_);
  not (_20840_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_20841_, _20796_, _20840_);
  and (_20842_, _20796_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_20843_, _20842_, _20841_);
  nor (_20844_, _20843_, _20789_);
  nor (_20845_, _20844_, _20839_);
  nor (_20846_, _20845_, _20835_);
  nor (_20847_, _20846_, _20833_);
  and (_20848_, _20847_, _20820_);
  not (_20849_, _20796_);
  and (_20850_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_20851_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_20852_, _20851_, _20850_);
  and (_20853_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_20854_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_20855_, _20854_, _20853_);
  and (_20856_, _20855_, _20852_);
  and (_20857_, _20856_, _20849_);
  and (_20858_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_20859_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_20860_, _20859_, _20858_);
  and (_20861_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_20862_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_20863_, _20862_, _20861_);
  and (_20864_, _20863_, _20860_);
  and (_20865_, _20864_, _20796_);
  or (_20866_, _20865_, _20790_);
  nor (_20867_, _20866_, _20857_);
  and (_20868_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_20869_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_20870_, _20869_, _20868_);
  and (_20871_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_20872_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_20873_, _20872_, _20871_);
  and (_20874_, _20873_, _20870_);
  nor (_20875_, _20874_, _20796_);
  and (_20876_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_20877_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_20878_, _20877_, _20876_);
  and (_20879_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_20880_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_20881_, _20880_, _20879_);
  and (_20882_, _20881_, _20878_);
  nor (_20883_, _20882_, _20849_);
  or (_20884_, _20883_, _20875_);
  and (_20885_, _20884_, _20790_);
  nor (_20886_, _20885_, _20867_);
  nor (_20887_, _20886_, _20848_);
  and (_20888_, _20887_, _20781_);
  nor (_20889_, _20777_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_20890_, _20889_, _20778_);
  and (_20891_, _20890_, _20887_);
  nor (_20892_, _20776_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20893_, _20892_, _20777_);
  and (_20894_, _20893_, _20887_);
  nor (_20895_, _20890_, _20887_);
  nor (_20896_, _20895_, _20891_);
  and (_20897_, _20774_, _20772_);
  and (_20898_, _20897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_20899_, _20897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_20900_, _20899_, _20898_);
  and (_20901_, _20900_, _20887_);
  nor (_20902_, _20900_, _20887_);
  and (_20903_, _20773_, _20772_);
  nor (_20904_, _20903_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_20905_, _20904_, _20897_);
  and (_20906_, _20905_, _20887_);
  nor (_20907_, _20905_, _20887_);
  nor (_20908_, _20907_, _20906_);
  not (_20909_, _20908_);
  and (_20910_, _20772_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20911_, _20910_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_20912_, _20911_, _20903_);
  and (_20913_, _20912_, _20887_);
  nor (_20914_, _20772_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20915_, _20914_, _20910_);
  and (_20916_, _20915_, _20887_);
  nor (_20917_, _20912_, _20887_);
  nor (_20918_, _20917_, _20913_);
  and (_20919_, _20770_, _20768_);
  nor (_20920_, _20919_, _23860_);
  and (_20921_, _20919_, _23860_);
  nor (_20922_, _20921_, _20920_);
  not (_20923_, _20922_);
  and (_20924_, _20923_, _20887_);
  nor (_20925_, _20923_, _20887_);
  and (_20926_, _20769_, _20768_);
  nor (_20927_, _20926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_20928_, _20927_, _20919_);
  and (_20929_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_20930_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_20931_, _20930_, _20929_);
  and (_20932_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_20933_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_20934_, _20933_, _20932_);
  and (_20935_, _20934_, _20931_);
  and (_20936_, _20935_, _20849_);
  and (_20937_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_20938_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_20939_, _20938_, _20937_);
  and (_20940_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_20941_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_20942_, _20941_, _20940_);
  and (_20943_, _20942_, _20939_);
  and (_20944_, _20943_, _20796_);
  or (_20945_, _20944_, _20790_);
  nor (_20946_, _20945_, _20936_);
  and (_20947_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_20948_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_20949_, _20948_, _20947_);
  and (_20950_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_20951_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_20952_, _20951_, _20950_);
  and (_20953_, _20952_, _20949_);
  and (_20954_, _20953_, _20849_);
  and (_20955_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_20956_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_20957_, _20956_, _20955_);
  and (_20958_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_20959_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_20960_, _20959_, _20958_);
  and (_20961_, _20960_, _20957_);
  and (_20962_, _20961_, _20796_);
  nor (_20963_, _20962_, _20954_);
  and (_20964_, _20963_, _20790_);
  nor (_20965_, _20964_, _20946_);
  nor (_20966_, _20965_, _20848_);
  and (_20967_, _20966_, _20928_);
  nor (_20968_, _20966_, _20928_);
  nor (_20969_, _20968_, _20967_);
  not (_20970_, _20969_);
  and (_20971_, _20768_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20972_, _20971_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_20973_, _20972_, _20926_);
  and (_20974_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_20975_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_20976_, _20975_, _20974_);
  and (_20977_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_20978_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_20979_, _20978_, _20977_);
  and (_20980_, _20979_, _20976_);
  and (_20981_, _20980_, _20849_);
  and (_20982_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_20983_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_20984_, _20983_, _20982_);
  and (_20985_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_20986_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_20987_, _20986_, _20985_);
  and (_20988_, _20987_, _20984_);
  and (_20989_, _20988_, _20796_);
  or (_20990_, _20989_, _20790_);
  nor (_20991_, _20990_, _20981_);
  and (_20992_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_20993_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_20994_, _20993_, _20992_);
  and (_20995_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_20996_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_20997_, _20996_, _20995_);
  and (_20998_, _20997_, _20994_);
  nor (_20999_, _20998_, _20796_);
  and (_21000_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_21001_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_21002_, _21001_, _21000_);
  and (_21003_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_21004_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_21005_, _21004_, _21003_);
  and (_21006_, _21005_, _21002_);
  nor (_21007_, _21006_, _20849_);
  or (_21008_, _21007_, _20999_);
  and (_21009_, _21008_, _20790_);
  nor (_21010_, _21009_, _20991_);
  nor (_21011_, _21010_, _20848_);
  and (_21012_, _21011_, _20973_);
  nor (_21013_, _21011_, _20973_);
  nor (_21014_, _21013_, _21012_);
  not (_21015_, _21014_);
  and (_21016_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_21017_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_21018_, _21017_, _21016_);
  and (_21019_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_21020_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_21021_, _21020_, _21019_);
  and (_21022_, _21021_, _21018_);
  and (_21023_, _21022_, _20849_);
  and (_21024_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_21025_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_21026_, _21025_, _21024_);
  and (_21027_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_21028_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_21029_, _21028_, _21027_);
  and (_21030_, _21029_, _21026_);
  and (_21031_, _21030_, _20796_);
  or (_21032_, _21031_, _20790_);
  nor (_21033_, _21032_, _21023_);
  and (_21034_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_21035_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_21036_, _21035_, _21034_);
  and (_21037_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_21038_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_21039_, _21038_, _21037_);
  and (_21040_, _21039_, _21036_);
  nor (_21041_, _21040_, _20796_);
  and (_21042_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_21043_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_21044_, _21043_, _21042_);
  and (_21045_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_21046_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_21047_, _21046_, _21045_);
  and (_21048_, _21047_, _21044_);
  nor (_21049_, _21048_, _20849_);
  or (_21050_, _21049_, _21041_);
  and (_21051_, _21050_, _20790_);
  nor (_21052_, _21051_, _21033_);
  nor (_21053_, _21052_, _20848_);
  nor (_21054_, _20768_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_21055_, _21054_, _20971_);
  and (_21056_, _21055_, _21053_);
  not (_21057_, _20787_);
  and (_21058_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_21059_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_21060_, _21059_, _21058_);
  and (_21061_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_21062_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_21063_, _21062_, _21061_);
  and (_21064_, _21063_, _21060_);
  and (_21065_, _21064_, _20849_);
  and (_21066_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_21067_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_21068_, _21067_, _21066_);
  and (_21069_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_21070_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_21071_, _21070_, _21069_);
  and (_21072_, _21071_, _21068_);
  and (_21073_, _21072_, _20796_);
  or (_21074_, _21073_, _20789_);
  nor (_21075_, _21074_, _21065_);
  and (_21076_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_21077_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_21078_, _21077_, _21076_);
  and (_21079_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_21080_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_21081_, _21080_, _21079_);
  and (_21082_, _21081_, _21078_);
  nor (_21083_, _21082_, _20796_);
  and (_21084_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_21085_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_21086_, _21085_, _21084_);
  and (_21087_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_21088_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_21089_, _21088_, _21087_);
  and (_21090_, _21089_, _21086_);
  nor (_21091_, _21090_, _20849_);
  or (_21092_, _21091_, _21083_);
  and (_21093_, _21092_, _20789_);
  nor (_21094_, _21093_, _21075_);
  nor (_21095_, _21094_, _20848_);
  and (_21096_, _21095_, _21057_);
  nor (_21097_, _21095_, _21057_);
  nor (_21098_, _21097_, _21096_);
  not (_21099_, _21098_);
  not (_21100_, _20794_);
  and (_21101_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_21102_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_21103_, _21102_, _21101_);
  and (_21104_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_21105_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_21106_, _21105_, _21104_);
  and (_21107_, _21106_, _21103_);
  and (_21108_, _21107_, _20849_);
  and (_21109_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_21110_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_21111_, _21110_, _21109_);
  and (_21112_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_21113_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_21114_, _21113_, _21112_);
  and (_21115_, _21114_, _21111_);
  and (_21116_, _21115_, _20796_);
  or (_21117_, _21116_, _20790_);
  nor (_21118_, _21117_, _21108_);
  and (_21119_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_21120_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_21121_, _21120_, _21119_);
  and (_21122_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_21123_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_21124_, _21123_, _21122_);
  and (_21125_, _21124_, _21121_);
  nor (_21126_, _21125_, _20796_);
  and (_21127_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_21128_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_21129_, _21128_, _21127_);
  and (_21130_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_21131_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_21132_, _21131_, _21130_);
  and (_21133_, _21132_, _21129_);
  nor (_21134_, _21133_, _20849_);
  or (_21135_, _21134_, _21126_);
  and (_21136_, _21135_, _20790_);
  nor (_21137_, _21136_, _21118_);
  nor (_21138_, _21137_, _20848_);
  and (_21139_, _21138_, _21100_);
  and (_21140_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_21141_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_21142_, _21141_, _21140_);
  and (_21143_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_21144_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_21145_, _21144_, _21143_);
  and (_21146_, _21145_, _21142_);
  and (_21147_, _21146_, _20849_);
  and (_21148_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_21149_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_21150_, _21149_, _21148_);
  and (_21151_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_21152_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_21153_, _21152_, _21151_);
  and (_21154_, _21153_, _21150_);
  and (_21155_, _21154_, _20796_);
  or (_21156_, _21155_, _20790_);
  nor (_21157_, _21156_, _21147_);
  and (_21158_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_21159_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_21160_, _21159_, _21158_);
  and (_21161_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_21162_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_21163_, _21162_, _21161_);
  and (_21164_, _21163_, _21160_);
  and (_21165_, _21164_, _20849_);
  and (_21166_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_21167_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_21168_, _21167_, _21166_);
  and (_21169_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_21170_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_21171_, _21170_, _21169_);
  and (_21172_, _21171_, _21168_);
  and (_21173_, _21172_, _20796_);
  nor (_21174_, _21173_, _21165_);
  and (_21175_, _21174_, _20790_);
  nor (_21176_, _21175_, _21157_);
  nor (_21177_, _21176_, _20848_);
  and (_21178_, _21177_, _23835_);
  and (_21179_, _20834_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_21180_, _20821_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_21181_, _21180_, _21179_);
  and (_21182_, _20807_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_21183_, _20782_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_21184_, _21183_, _21182_);
  and (_21185_, _21184_, _21181_);
  and (_21186_, _21185_, _20849_);
  and (_21187_, _20834_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_21188_, _20821_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_21189_, _21188_, _21187_);
  and (_21190_, _20807_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_21191_, _20782_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_21192_, _21191_, _21190_);
  and (_21193_, _21192_, _21189_);
  and (_21194_, _21193_, _20796_);
  or (_21195_, _21194_, _20790_);
  nor (_21196_, _21195_, _21186_);
  and (_21197_, _20834_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_21198_, _20782_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_21199_, _21198_, _21197_);
  and (_21200_, _20807_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_21201_, _20821_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_21202_, _21201_, _21200_);
  and (_21203_, _21202_, _21199_);
  nor (_21204_, _21203_, _20796_);
  and (_21205_, _20834_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_21206_, _20821_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_21207_, _21206_, _21205_);
  and (_21208_, _20807_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_21209_, _20782_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_21210_, _21209_, _21208_);
  and (_21211_, _21210_, _21207_);
  nor (_21212_, _21211_, _20849_);
  or (_21213_, _21212_, _21204_);
  and (_21214_, _21213_, _20790_);
  nor (_21215_, _21214_, _21196_);
  nor (_21216_, _21215_, _20848_);
  and (_21217_, _21216_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21218_, _21177_, _23835_);
  nor (_21219_, _21218_, _21178_);
  and (_21220_, _21219_, _21217_);
  nor (_21221_, _21220_, _21178_);
  nor (_21222_, _21138_, _21100_);
  nor (_21223_, _21222_, _21139_);
  not (_21224_, _21223_);
  nor (_21225_, _21224_, _21221_);
  nor (_21226_, _21225_, _21139_);
  nor (_21227_, _21226_, _21099_);
  nor (_21228_, _21227_, _21096_);
  nor (_21229_, _21055_, _21053_);
  nor (_21230_, _21229_, _21056_);
  not (_21231_, _21230_);
  nor (_21232_, _21231_, _21228_);
  nor (_21233_, _21232_, _21056_);
  nor (_21234_, _21233_, _21015_);
  nor (_21235_, _21234_, _21012_);
  nor (_21236_, _21235_, _20970_);
  nor (_21237_, _21236_, _20967_);
  nor (_21238_, _21237_, _20925_);
  or (_21239_, _21238_, _20924_);
  nor (_21240_, _20915_, _20887_);
  nor (_21241_, _21240_, _20916_);
  and (_21242_, _21241_, _21239_);
  and (_21243_, _21242_, _20918_);
  or (_21244_, _21243_, _20916_);
  nor (_21245_, _21244_, _20913_);
  nor (_21246_, _21245_, _20909_);
  nor (_21247_, _21246_, _20906_);
  nor (_21248_, _21247_, _20902_);
  nor (_21249_, _21248_, _20901_);
  nor (_21250_, _20893_, _20887_);
  nor (_21251_, _21250_, _20894_);
  not (_21252_, _21251_);
  nor (_21253_, _21252_, _21249_);
  and (_21254_, _21253_, _20896_);
  or (_21255_, _21254_, _20894_);
  nor (_21256_, _21255_, _20891_);
  nor (_21257_, _20887_, _20781_);
  nor (_21258_, _21257_, _20888_);
  not (_21259_, _21258_);
  nor (_21260_, _21259_, _21256_);
  nor (_21261_, _21260_, _20888_);
  nor (_21262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_21263_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_21264_, _21263_, _21262_);
  not (_21265_, _21264_);
  and (_21266_, _21265_, _20779_);
  nor (_21267_, _21265_, _20779_);
  nor (_21268_, _21267_, _21266_);
  not (_21269_, _21268_);
  and (_21270_, _21269_, _20887_);
  nor (_21271_, _21269_, _20887_);
  nor (_21272_, _21271_, _21270_);
  not (_21273_, _21272_);
  nand (_21274_, _21273_, _21261_);
  or (_21275_, _21273_, _21261_);
  and (_21276_, _21275_, _21274_);
  and (_21277_, _21259_, _21256_);
  nor (_21278_, _21277_, _21260_);
  and (_21279_, _21278_, _23824_);
  nor (_21280_, _21278_, _23824_);
  nor (_21281_, _21253_, _20894_);
  nor (_21282_, _20890_, _23820_);
  and (_21283_, _20890_, _23820_);
  or (_21284_, _21283_, _21282_);
  nand (_21285_, _21284_, _20887_);
  or (_21286_, _21284_, _20887_);
  and (_21287_, _21286_, _21285_);
  not (_21288_, _21287_);
  nand (_21289_, _21288_, _21281_);
  or (_21290_, _21288_, _21281_);
  and (_21291_, _21290_, _21289_);
  and (_21292_, _21252_, _21249_);
  nor (_21293_, _21292_, _21253_);
  nand (_21294_, _21293_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_21295_, _21293_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_21296_, _21295_, _21294_);
  nor (_21297_, _20900_, _23811_);
  and (_21298_, _20900_, _23811_);
  or (_21299_, _21298_, _21297_);
  nand (_21300_, _21299_, _20887_);
  or (_21301_, _21299_, _20887_);
  and (_21302_, _21301_, _21300_);
  not (_21303_, _21302_);
  nand (_21304_, _21303_, _21247_);
  or (_21305_, _21303_, _21247_);
  and (_21306_, _21305_, _21304_);
  and (_21307_, _21245_, _20909_);
  nor (_21308_, _21307_, _21246_);
  nand (_21309_, _21308_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_21310_, _21308_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_21311_, _21310_, _21309_);
  nor (_21312_, _21241_, _21239_);
  nor (_21313_, _21312_, _21242_);
  nor (_21314_, _21313_, _23798_);
  nor (_21315_, _20924_, _20925_);
  nor (_21316_, _21315_, _21237_);
  and (_21317_, _21315_, _21237_);
  or (_21318_, _21317_, _21316_);
  and (_21319_, _21318_, _23794_);
  nor (_21320_, _21318_, _23794_);
  and (_21321_, _21235_, _20970_);
  nor (_21322_, _21321_, _21236_);
  nor (_21323_, _21322_, _23790_);
  and (_21324_, _21322_, _23790_);
  and (_21325_, _21233_, _21015_);
  nor (_21326_, _21325_, _21234_);
  and (_21327_, _21326_, _23786_);
  nor (_21328_, _21326_, _23786_);
  and (_21329_, _21231_, _21228_);
  nor (_21330_, _21329_, _21232_);
  and (_21331_, _21330_, _23782_);
  nor (_21332_, _21330_, _23782_);
  and (_21333_, _21226_, _21099_);
  nor (_21334_, _21333_, _21227_);
  nor (_21335_, _21334_, _23778_);
  and (_21336_, _21334_, _23778_);
  and (_21337_, _21224_, _21221_);
  nor (_21338_, _21337_, _21225_);
  nor (_21339_, _21338_, _23774_);
  and (_21340_, _21338_, _23774_);
  and (_21341_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21342_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_21343_, _21342_, _21341_);
  not (_21344_, _21343_);
  nand (_21345_, _21344_, _21216_);
  or (_21346_, _21344_, _21216_);
  and (_21347_, _21346_, _21345_);
  nor (_21348_, _21219_, _21217_);
  nor (_21349_, _21348_, _21220_);
  and (_21350_, _21349_, _23769_);
  nor (_21351_, _21349_, _23769_);
  or (_21352_, _21351_, _21350_);
  or (_21353_, _21352_, _21347_);
  or (_21354_, _21353_, _21340_);
  or (_21355_, _21354_, _21339_);
  or (_21356_, _21355_, _21336_);
  or (_21357_, _21356_, _21335_);
  or (_21358_, _21357_, _21332_);
  or (_21359_, _21358_, _21331_);
  or (_21360_, _21359_, _21328_);
  or (_21361_, _21360_, _21327_);
  or (_21362_, _21361_, _21324_);
  or (_21363_, _21362_, _21323_);
  or (_21364_, _21363_, _21320_);
  or (_21365_, _21364_, _21319_);
  or (_21366_, _21365_, _21314_);
  nor (_21367_, _21242_, _20916_);
  and (_21368_, _20918_, _23802_);
  nor (_21369_, _20918_, _23802_);
  nor (_21370_, _21369_, _21368_);
  not (_21371_, _21370_);
  nor (_21372_, _21371_, _21367_);
  and (_21373_, _21313_, _23798_);
  and (_21374_, _21371_, _21367_);
  or (_21375_, _21374_, _21373_);
  or (_21376_, _21375_, _21372_);
  or (_21377_, _21376_, _21366_);
  or (_21378_, _21377_, _21311_);
  or (_21379_, _21378_, _21306_);
  or (_21380_, _21379_, _21296_);
  or (_21381_, _21380_, _21291_);
  or (_21382_, _21381_, _21280_);
  or (_21383_, _21382_, _21279_);
  or (_21384_, _21383_, _21276_);
  and (_21385_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21386_, _21385_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_21387_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21388_, _21387_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_21389_, _21388_, _21386_);
  not (_21390_, _21389_);
  nor (_21391_, _21386_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21392_, _21386_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21393_, _21392_, _21391_);
  nand (_21394_, _21393_, _20813_);
  or (_21395_, _21393_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_21396_, _21395_, _21394_);
  and (_21397_, _21396_, _21390_);
  not (_21398_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_21399_, _21393_, _21398_);
  or (_21400_, _21393_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_21401_, _21400_, _21389_);
  and (_21402_, _21401_, _21399_);
  or (_21403_, _21402_, _21397_);
  or (_21404_, _21403_, _23769_);
  and (_21405_, _23774_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21406_, \oc8051_symbolic_cxrom1.regvalid [5], _23778_);
  and (_21407_, \oc8051_symbolic_cxrom1.regvalid [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21408_, _21407_, _21406_);
  and (_21409_, _21408_, _21405_);
  or (_21410_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21411_, \oc8051_symbolic_cxrom1.regvalid [1], _23778_);
  and (_21412_, _21411_, _21385_);
  and (_21413_, _21412_, _21410_);
  or (_21414_, _21413_, _21409_);
  nor (_21415_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21416_, _21415_, _23774_);
  nor (_21417_, _21416_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21418_, _21416_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21419_, _21418_, _21417_);
  and (_21420_, _21419_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_21421_, _21415_, _23774_);
  nor (_21422_, _21421_, _21416_);
  or (_21423_, _05018_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_21424_, _21423_, _21422_);
  or (_21425_, _21424_, _21420_);
  and (_21426_, _21425_, _23769_);
  nor (_21427_, _21419_, _05011_);
  and (_21428_, _21419_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_21429_, _21428_, _21427_);
  or (_21430_, _21429_, _21422_);
  and (_21431_, _21430_, _21426_);
  or (_21432_, _21431_, _21414_);
  and (_21433_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21434_, \oc8051_symbolic_cxrom1.regvalid [6], _23778_);
  or (_21435_, _21434_, _23774_);
  or (_21436_, _21435_, _21433_);
  or (_21437_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21438_, \oc8051_symbolic_cxrom1.regvalid [10], _23778_);
  and (_21439_, _21438_, _21437_);
  or (_21440_, _21439_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21441_, _21440_, _21436_);
  and (_21442_, _21441_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21443_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21444_, \oc8051_symbolic_cxrom1.regvalid [0], _23778_);
  or (_21445_, _21444_, _21443_);
  and (_21446_, _21445_, _23774_);
  and (_21447_, \oc8051_symbolic_cxrom1.regvalid [4], _23778_);
  and (_21448_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21449_, _21448_, _21447_);
  and (_21450_, _21449_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21451_, _21450_, _21446_);
  and (_21452_, _21451_, _23769_);
  or (_21453_, _21452_, _21442_);
  and (_21454_, _21453_, _23765_);
  and (_21455_, _21405_, _21449_);
  or (_21456_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21457_, \oc8051_symbolic_cxrom1.regvalid [0], _23778_);
  and (_21458_, _21457_, _21385_);
  and (_21459_, _21458_, _21456_);
  or (_21460_, _21459_, _21455_);
  and (_21461_, _21441_, _23769_);
  or (_21462_, _21461_, _21460_);
  and (_21463_, _21462_, _21454_);
  nand (_21464_, _21393_, _05024_);
  or (_21465_, _21393_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_21466_, _21465_, _21464_);
  and (_21467_, _21466_, _21390_);
  nand (_21468_, _21393_, _04986_);
  or (_21469_, _21393_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_21470_, _21469_, _21389_);
  and (_21471_, _21470_, _21468_);
  or (_21472_, _21471_, _21467_);
  or (_21473_, _21472_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21474_, _21473_, _21463_);
  and (_21475_, _21474_, _21432_);
  and (_21476_, _21475_, _21404_);
  or (_21477_, \oc8051_symbolic_cxrom1.regvalid [10], _23769_);
  or (_21478_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_21479_, _21478_, _21477_);
  nand (_21480_, _21479_, _21419_);
  or (_21481_, \oc8051_symbolic_cxrom1.regvalid [2], _23769_);
  or (_21482_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21483_, _21482_, _21481_);
  or (_21484_, _21483_, _21419_);
  and (_21485_, _21484_, _21480_);
  or (_21486_, _21485_, _21422_);
  nor (_21487_, _21393_, _05035_);
  and (_21488_, _21393_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_21489_, _21488_, _21487_);
  and (_21490_, _21489_, _21390_);
  or (_21491_, _21393_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_21492_, \oc8051_symbolic_cxrom1.regvalid [12], _23778_);
  and (_21493_, _21492_, _21389_);
  and (_21494_, _21493_, _21491_);
  or (_21495_, _21494_, _23769_);
  or (_21496_, _21495_, _21490_);
  nand (_21497_, \oc8051_symbolic_cxrom1.regvalid [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_21498_, _21497_, _21423_);
  or (_21499_, _21498_, _23774_);
  or (_21500_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21501_, \oc8051_symbolic_cxrom1.regvalid [11], _23778_);
  and (_21502_, _21501_, _21500_);
  or (_21503_, _21502_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21504_, _21503_, _21499_);
  and (_21505_, _21504_, _21387_);
  and (_21506_, _23769_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_21507_, _21408_, _23774_);
  or (_21508_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21509_, \oc8051_symbolic_cxrom1.regvalid [9], _23778_);
  and (_21510_, _21509_, _21508_);
  or (_21511_, _21510_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21512_, _21511_, _21507_);
  and (_21513_, _21512_, _21506_);
  or (_21514_, _21513_, _21505_);
  and (_21515_, _21504_, _23769_);
  or (_21516_, _21515_, _21414_);
  and (_21517_, _21516_, _21514_);
  and (_21518_, _21517_, _21496_);
  and (_21519_, _21518_, _21486_);
  or (_21520_, _21393_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_21521_, \oc8051_symbolic_cxrom1.regvalid [14], _23778_);
  and (_21522_, _21521_, _21520_);
  or (_21523_, _21522_, _21390_);
  nand (_21524_, _21393_, _20840_);
  or (_21525_, _21393_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_21526_, _21525_, _21524_);
  or (_21527_, _21526_, _21389_);
  and (_21528_, _21527_, _21523_);
  or (_21529_, _21528_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21530_, _21419_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_21531_, _21434_, _23769_);
  or (_21532_, _21531_, _21530_);
  and (_21533_, _21419_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_21534_, _21447_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_21535_, _21534_, _21533_);
  nand (_21536_, _21535_, _21532_);
  nand (_21537_, _21536_, _21422_);
  and (_21538_, _21537_, _21529_);
  and (_21539_, _21538_, _21519_);
  or (_21540_, _21539_, _21476_);
  nor (_21541_, _20782_, _23840_);
  and (_21542_, _20791_, _23835_);
  nor (_21543_, _21542_, _21541_);
  not (_21544_, _21543_);
  and (_21545_, _21541_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21546_, _21541_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21547_, _21546_, _21545_);
  and (_21548_, _21547_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_21549_, _21547_, _05011_);
  or (_21550_, _21549_, _21548_);
  and (_21551_, _21550_, _21544_);
  nand (_21552_, _21547_, _21398_);
  nor (_21553_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21554_, _21553_, _21544_);
  and (_21555_, _21554_, _21552_);
  or (_21556_, _21555_, _21551_);
  and (_21557_, _21556_, _20782_);
  and (_21558_, _21547_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_21559_, _21547_, _05474_);
  or (_21560_, _21559_, _21558_);
  and (_21561_, _21560_, _21544_);
  or (_21562_, _21547_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_21563_, _04986_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21564_, _21563_, _21544_);
  and (_21565_, _21564_, _21562_);
  or (_21566_, _21565_, _21561_);
  and (_21567_, _21566_, _20807_);
  or (_21568_, _21567_, _21557_);
  and (_21569_, _21547_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_21570_, _21547_, _05054_);
  or (_21571_, _21570_, _21569_);
  and (_21572_, _21571_, _21544_);
  nand (_21573_, _21547_, _05049_);
  nor (_21574_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21575_, _21574_, _21544_);
  and (_21576_, _21575_, _21573_);
  or (_21577_, _21576_, _21572_);
  and (_21578_, _21577_, _20821_);
  and (_21579_, _21547_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_21580_, _21547_, _05035_);
  or (_21581_, _21580_, _21579_);
  and (_21582_, _21581_, _21544_);
  or (_21583_, _21547_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_21584_, _05041_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21585_, _21584_, _21544_);
  and (_21586_, _21585_, _21583_);
  or (_21587_, _21586_, _21582_);
  and (_21588_, _21587_, _20834_);
  or (_21589_, _21588_, _21578_);
  or (_21590_, _21589_, _21568_);
  nor (_21591_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21592_, _21591_, _21584_);
  and (_21593_, _21592_, _20793_);
  nor (_21594_, _21593_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21595_, _05049_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21596_, _21595_);
  nor (_21597_, _21574_, _23840_);
  and (_21598_, _21597_, _21596_);
  and (_21599_, _20840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21600_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21601_, _21600_, _21599_);
  and (_21602_, _21601_, _23840_);
  nor (_21603_, _21602_, _21598_);
  nor (_21604_, _21603_, _23835_);
  nor (_21605_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21606_, _20827_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21607_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21608_, _21607_, _21606_);
  and (_21609_, _21608_, _21605_);
  nor (_21610_, _21609_, _21604_);
  and (_21611_, _21610_, _21594_);
  and (_21612_, _21398_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21613_, _21612_);
  nor (_21614_, _21553_, _23840_);
  and (_21615_, _21614_, _21613_);
  and (_21616_, _20813_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21617_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21618_, _21617_, _21616_);
  and (_21619_, _21618_, _23840_);
  nor (_21620_, _21619_, _21615_);
  nor (_21621_, _21620_, _23835_);
  nor (_21622_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_21623_, _05024_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21624_, _21623_, _21622_);
  and (_21625_, _21624_, _21605_);
  nor (_21626_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21627_, _21626_, _21563_);
  and (_21628_, _21627_, _20793_);
  or (_21629_, _21628_, _23830_);
  or (_21630_, _21629_, _21625_);
  nor (_21631_, _21630_, _21621_);
  nor (_21632_, _21631_, _21611_);
  nor (_21633_, _21603_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21634_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21635_, _21634_);
  not (_21636_, _20767_);
  and (_21637_, _05035_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21638_, _21637_, _21636_);
  and (_21639_, _21638_, _21635_);
  and (_21640_, _21592_, _20792_);
  or (_21641_, _21640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_21642_, _21641_, _21639_);
  nor (_21643_, _21642_, _21633_);
  nor (_21644_, _21620_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21645_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21646_, _21645_);
  and (_21647_, _05474_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21648_, _21647_, _21636_);
  and (_21649_, _21648_, _21646_);
  and (_21650_, _21627_, _20792_);
  or (_21651_, _21650_, _23830_);
  or (_21652_, _21651_, _21649_);
  nor (_21653_, _21652_, _21644_);
  nor (_21654_, _21653_, _21643_);
  not (_21655_, _23763_);
  nor (_21656_, _21655_, first_instr);
  and (_21657_, _21656_, _21654_);
  and (_21658_, _21657_, _21632_);
  nand (_21659_, _21658_, _21590_);
  nor (_21660_, _21659_, _20848_);
  and (_21661_, _21660_, _21540_);
  nor (_21662_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21663_, _06664_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21664_, _21663_, _21662_);
  and (_21665_, _21664_, _20792_);
  nor (_21666_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21667_, _06944_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21668_, _21667_, _21666_);
  and (_21669_, _21668_, _20793_);
  nor (_21670_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21671_, _06376_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21672_, _21671_, _21670_);
  and (_21673_, _21672_, _21605_);
  nor (_21674_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21675_, _07185_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21676_, _21675_, _21674_);
  and (_21677_, _21676_, _20767_);
  or (_21678_, _21677_, _21673_);
  or (_21679_, _21678_, _21669_);
  or (_21680_, _21679_, _21665_);
  and (_21681_, _21680_, _23844_);
  nor (_21682_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21683_, _07778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21684_, _21683_, _21682_);
  and (_21685_, _21684_, _20792_);
  nor (_21686_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21687_, _08052_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21688_, _21687_, _21686_);
  and (_21689_, _21688_, _20793_);
  nor (_21690_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21691_, _07520_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21692_, _21691_, _21690_);
  and (_21693_, _21692_, _21605_);
  nor (_21694_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21695_, _08319_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21696_, _21695_, _21694_);
  and (_21697_, _21696_, _20767_);
  or (_21698_, _21697_, _21693_);
  or (_21699_, _21698_, _21689_);
  or (_21700_, _21699_, _21685_);
  and (_21701_, _21700_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21702_, _21701_, _21681_);
  and (_21703_, _21702_, _21632_);
  nor (_21704_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21705_, _06642_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21706_, _21705_, _21704_);
  and (_21707_, _21706_, _20792_);
  nor (_21708_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21709_, _06929_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21710_, _21709_, _21708_);
  and (_21711_, _21710_, _20793_);
  nor (_21712_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21713_, _06353_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21714_, _21713_, _21712_);
  and (_21715_, _21714_, _21605_);
  nor (_21716_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21717_, _07157_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21718_, _21717_, _21716_);
  and (_21719_, _21718_, _20767_);
  or (_21720_, _21719_, _21715_);
  or (_21721_, _21720_, _21711_);
  or (_21722_, _21721_, _21707_);
  and (_21723_, _21722_, _23844_);
  nor (_21724_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21725_, _07758_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21726_, _21725_, _21724_);
  and (_21727_, _21726_, _20792_);
  nor (_21728_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21729_, _08025_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21730_, _21729_, _21728_);
  and (_21731_, _21730_, _20793_);
  nor (_21732_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21733_, _07498_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21734_, _21733_, _21732_);
  and (_21735_, _21734_, _21605_);
  nor (_21736_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21737_, _08305_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21738_, _21737_, _21736_);
  and (_21739_, _21738_, _20767_);
  or (_21740_, _21739_, _21735_);
  or (_21741_, _21740_, _21731_);
  or (_21742_, _21741_, _21727_);
  and (_21743_, _21742_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21744_, _21743_, _21723_);
  and (_21745_, _21744_, _21632_);
  nor (_21746_, _21745_, _21703_);
  nor (_21747_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21748_, _06703_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21749_, _21748_, _21747_);
  and (_21750_, _21749_, _20792_);
  nor (_21751_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21752_, _06972_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21753_, _21752_, _21751_);
  and (_21754_, _21753_, _20793_);
  nor (_21755_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21756_, _06404_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21757_, _21756_, _21755_);
  and (_21758_, _21757_, _21605_);
  nor (_21759_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21760_, _07218_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21761_, _21760_, _21759_);
  and (_21762_, _21761_, _20767_);
  or (_21763_, _21762_, _21758_);
  or (_21764_, _21763_, _21754_);
  or (_21765_, _21764_, _21750_);
  and (_21766_, _21765_, _23844_);
  nor (_21767_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21768_, _07806_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21769_, _21768_, _21767_);
  and (_21770_, _21769_, _20792_);
  nor (_21771_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21772_, _08077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21773_, _21772_, _21771_);
  and (_21774_, _21773_, _20793_);
  nor (_21775_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21776_, _07549_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21777_, _21776_, _21775_);
  and (_21778_, _21777_, _21605_);
  nor (_21779_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21780_, _08346_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21781_, _21780_, _21779_);
  and (_21782_, _21781_, _20767_);
  or (_21783_, _21782_, _21778_);
  or (_21784_, _21783_, _21774_);
  or (_21785_, _21784_, _21770_);
  and (_21786_, _21785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21787_, _21786_, _21766_);
  and (_21788_, _21787_, _21632_);
  nor (_21789_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21790_, _06686_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21791_, _21790_, _21789_);
  and (_21792_, _21791_, _20792_);
  nor (_21793_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21794_, _06958_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21795_, _21794_, _21793_);
  and (_21796_, _21795_, _20793_);
  nor (_21797_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21798_, _06391_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21799_, _21798_, _21797_);
  and (_21800_, _21799_, _21605_);
  nor (_21801_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21802_, _07200_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21803_, _21802_, _21801_);
  and (_21804_, _21803_, _20767_);
  or (_21805_, _21804_, _21800_);
  or (_21806_, _21805_, _21796_);
  or (_21807_, _21806_, _21792_);
  and (_21808_, _21807_, _23844_);
  nor (_21809_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21810_, _07791_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21811_, _21810_, _21809_);
  and (_21812_, _21811_, _20792_);
  nor (_21813_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21814_, _08065_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21815_, _21814_, _21813_);
  and (_21816_, _21815_, _20793_);
  nor (_21817_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21818_, _07531_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21819_, _21818_, _21817_);
  and (_21820_, _21819_, _21605_);
  nor (_21821_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21822_, _08333_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21823_, _21822_, _21821_);
  and (_21824_, _21823_, _20767_);
  or (_21825_, _21824_, _21820_);
  or (_21826_, _21825_, _21816_);
  or (_21827_, _21826_, _21812_);
  and (_21828_, _21827_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21829_, _21828_, _21808_);
  and (_21830_, _21829_, _21632_);
  nor (_21831_, _21830_, _21788_);
  and (_21832_, _21831_, _21746_);
  nor (_21833_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21834_, _05099_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21835_, _21834_, _21833_);
  and (_21836_, _21835_, _20793_);
  nor (_21837_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21838_, _05092_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21839_, _21838_, _21837_);
  and (_21840_, _21839_, _21605_);
  nor (_21841_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21842_, _05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21843_, _21842_, _21841_);
  and (_21844_, _21843_, _20767_);
  or (_21845_, _21844_, _21840_);
  nor (_21846_, _21845_, _21836_);
  nor (_21847_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21848_, _05111_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21849_, _21848_, _21847_);
  and (_21850_, _21849_, _20792_);
  nor (_21851_, _21850_, _23844_);
  and (_21852_, _21851_, _21846_);
  nor (_21853_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21854_, _05072_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21855_, _21854_, _21853_);
  and (_21856_, _21855_, _20767_);
  nor (_21857_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21858_, _05077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21859_, _21858_, _21857_);
  and (_21860_, _21859_, _20793_);
  nor (_21861_, _21860_, _21856_);
  nor (_21862_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21863_, _05083_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21864_, _21863_, _21862_);
  and (_21865_, _21864_, _20792_);
  nor (_21866_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21867_, _05065_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21868_, _21867_, _21866_);
  and (_21869_, _21868_, _21605_);
  nor (_21870_, _21869_, _21865_);
  and (_21871_, _21870_, _21861_);
  and (_21872_, _21871_, _23844_);
  nor (_21873_, _21872_, _21852_);
  and (_21874_, _21873_, _21632_);
  nor (_21875_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21876_, _07279_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21877_, _21876_, _21875_);
  and (_21878_, _21877_, _20767_);
  nor (_21879_, _21878_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21880_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21881_, _06447_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21882_, _21881_, _21880_);
  and (_21883_, _21882_, _21605_);
  not (_21884_, _21883_);
  nor (_21885_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21886_, _06745_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21887_, _21886_, _21885_);
  and (_21888_, _21887_, _20792_);
  nor (_21889_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21890_, _07013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21891_, _21890_, _21889_);
  and (_21892_, _21891_, _20793_);
  nor (_21893_, _21892_, _21888_);
  and (_21894_, _21893_, _21884_);
  and (_21895_, _21894_, _21879_);
  nor (_21896_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21897_, _08383_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21898_, _21897_, _21896_);
  and (_21899_, _21898_, _20767_);
  nor (_21900_, _21899_, _23844_);
  nor (_21901_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21902_, _07597_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21903_, _21902_, _21901_);
  and (_21904_, _21903_, _21605_);
  not (_21905_, _21904_);
  nor (_21906_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21907_, _07842_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21908_, _21907_, _21906_);
  and (_21909_, _21908_, _20792_);
  nor (_21910_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21911_, _08118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21912_, _21911_, _21910_);
  and (_21913_, _21912_, _20793_);
  nor (_21914_, _21913_, _21909_);
  and (_21915_, _21914_, _21905_);
  and (_21916_, _21915_, _21900_);
  nor (_21917_, _21916_, _21895_);
  and (_21918_, _21917_, _21632_);
  not (_21919_, _21918_);
  and (_21920_, _21919_, _21874_);
  nor (_21921_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21922_, _06419_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21923_, _21922_, _21921_);
  and (_21924_, _21923_, _21605_);
  nor (_21925_, _21924_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21926_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21927_, _06987_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21928_, _21927_, _21926_);
  and (_21929_, _21928_, _20793_);
  not (_21930_, _21929_);
  nor (_21931_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21932_, _06716_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21933_, _21932_, _21931_);
  and (_21934_, _21933_, _20792_);
  nor (_21935_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21936_, _07238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21937_, _21936_, _21935_);
  and (_21938_, _21937_, _20767_);
  nor (_21939_, _21938_, _21934_);
  and (_21940_, _21939_, _21930_);
  and (_21941_, _21940_, _21925_);
  nor (_21942_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21943_, _07561_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21944_, _21943_, _21942_);
  and (_21945_, _21944_, _21605_);
  nor (_21946_, _21945_, _23844_);
  nor (_21947_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21948_, _08089_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21949_, _21948_, _21947_);
  and (_21950_, _21949_, _20793_);
  not (_21951_, _21950_);
  nor (_21952_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21953_, _07818_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21954_, _21953_, _21952_);
  and (_21955_, _21954_, _20792_);
  nor (_21956_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21957_, _08359_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21958_, _21957_, _21956_);
  and (_21959_, _21958_, _20767_);
  nor (_21960_, _21959_, _21955_);
  and (_21961_, _21960_, _21951_);
  and (_21962_, _21961_, _21946_);
  nor (_21963_, _21962_, _21941_);
  and (_21964_, _21963_, _21632_);
  nor (_21965_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21966_, _06430_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21967_, _21966_, _21965_);
  and (_21968_, _21967_, _21605_);
  nor (_21969_, _21968_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21970_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21971_, _07000_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21972_, _21971_, _21970_);
  and (_21973_, _21972_, _20793_);
  not (_21974_, _21973_);
  nor (_21975_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21976_, _06728_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21977_, _21976_, _21975_);
  and (_21978_, _21977_, _20792_);
  nor (_21979_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21980_, _07257_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21981_, _21980_, _21979_);
  and (_21982_, _21981_, _20767_);
  nor (_21983_, _21982_, _21978_);
  and (_21984_, _21983_, _21974_);
  and (_21985_, _21984_, _21969_);
  nor (_21986_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21987_, _07581_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21988_, _21987_, _21986_);
  and (_21989_, _21988_, _21605_);
  nor (_21990_, _21989_, _23844_);
  nor (_21991_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21992_, _08103_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21993_, _21992_, _21991_);
  and (_21994_, _21993_, _20793_);
  not (_21995_, _21994_);
  nor (_21996_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21997_, _07830_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21998_, _21997_, _21996_);
  and (_21999_, _21998_, _20792_);
  nor (_22000_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22001_, _08370_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22002_, _22001_, _22000_);
  and (_22003_, _22002_, _20767_);
  nor (_22004_, _22003_, _21999_);
  and (_22005_, _22004_, _21995_);
  and (_22006_, _22005_, _21990_);
  nor (_22007_, _22006_, _21985_);
  and (_22008_, _22007_, _21632_);
  nor (_22009_, _22008_, _21964_);
  and (_22010_, _22009_, _21920_);
  and (_22011_, _22010_, _21832_);
  and (_22012_, _22011_, _21661_);
  and (_22013_, _22012_, _21384_);
  and (_22014_, _21726_, _21605_);
  and (_22015_, _21738_, _20793_);
  and (_22016_, _21734_, _20767_);
  and (_22017_, _21730_, _20792_);
  or (_22018_, _22017_, _22016_);
  or (_22019_, _22018_, _22015_);
  or (_22020_, _22019_, _22014_);
  and (_22021_, _22020_, _21057_);
  and (_22022_, _21706_, _21605_);
  and (_22023_, _21718_, _20793_);
  and (_22024_, _21714_, _20767_);
  and (_22025_, _21710_, _20792_);
  or (_22026_, _22025_, _22024_);
  or (_22027_, _22026_, _22023_);
  or (_22028_, _22027_, _22022_);
  and (_22029_, _22028_, _20787_);
  or (_22030_, _22029_, _22021_);
  and (_22031_, _22030_, _21654_);
  nand (_22032_, _22031_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_22033_, _22031_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_22034_, _22033_, _22032_);
  and (_22035_, _21696_, _20793_);
  and (_22036_, _21688_, _20792_);
  nor (_22037_, _22036_, _22035_);
  and (_22038_, _21684_, _21605_);
  and (_22039_, _21692_, _23844_);
  nor (_22040_, _22039_, _22038_);
  and (_22041_, _22040_, _22037_);
  nor (_22042_, _22041_, _20787_);
  and (_22043_, _21676_, _20793_);
  and (_22044_, _21668_, _20792_);
  nor (_22045_, _22044_, _22043_);
  and (_22046_, _21664_, _21605_);
  and (_22047_, _21672_, _20767_);
  nor (_22048_, _22047_, _22046_);
  and (_22049_, _22048_, _22045_);
  nor (_22050_, _22049_, _21057_);
  nor (_22051_, _22050_, _22042_);
  not (_22052_, _22051_);
  and (_22053_, _22052_, _21654_);
  and (_22054_, _22053_, _23769_);
  nor (_22055_, _22053_, _23769_);
  or (_22056_, _22055_, _22054_);
  or (_22057_, _22056_, _22034_);
  and (_22058_, _21795_, _20792_);
  or (_22059_, _22058_, _21057_);
  and (_22060_, _21799_, _20767_);
  and (_22061_, _21791_, _21605_);
  or (_22062_, _22061_, _22060_);
  and (_22063_, _21803_, _20793_);
  or (_22064_, _22063_, _22062_);
  or (_22065_, _22064_, _22059_);
  and (_22066_, _21815_, _20792_);
  or (_22067_, _22066_, _20787_);
  and (_22068_, _21819_, _20767_);
  and (_22069_, _21811_, _21605_);
  and (_22070_, _21823_, _20793_);
  or (_22071_, _22070_, _22069_);
  or (_22072_, _22071_, _22068_);
  or (_22073_, _22072_, _22067_);
  and (_22074_, _22073_, _22065_);
  and (_22075_, _22074_, _21654_);
  or (_22076_, _22075_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_22077_, _22075_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_22078_, _22077_, _22076_);
  and (_22079_, _21753_, _20792_);
  or (_22080_, _22079_, _21057_);
  and (_22081_, _21757_, _20767_);
  and (_22082_, _21749_, _21605_);
  or (_22083_, _22082_, _22081_);
  and (_22084_, _21761_, _20793_);
  or (_22085_, _22084_, _22083_);
  or (_22086_, _22085_, _22080_);
  and (_22087_, _21773_, _20792_);
  and (_22088_, _21781_, _20793_);
  and (_22089_, _21777_, _20767_);
  or (_22090_, _22089_, _22088_);
  or (_22091_, _22090_, _22087_);
  and (_22092_, _21769_, _21605_);
  or (_22093_, _22092_, _20787_);
  or (_22094_, _22093_, _22091_);
  and (_22095_, _22094_, _22086_);
  and (_22096_, _22095_, _21654_);
  nand (_22097_, _22096_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22098_, _22096_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22099_, _22098_, _22097_);
  or (_22100_, _22099_, _22078_);
  or (_22101_, _22100_, _22057_);
  and (_22102_, _21855_, _20793_);
  and (_22103_, _21868_, _20767_);
  and (_22104_, _21859_, _20792_);
  or (_22105_, _22104_, _22103_);
  nor (_22106_, _22105_, _22102_);
  and (_22107_, _21864_, _21605_);
  nor (_22108_, _22107_, _21057_);
  and (_22109_, _22108_, _22106_);
  and (_22110_, _21843_, _20793_);
  and (_22111_, _21835_, _20792_);
  nor (_22112_, _22111_, _22110_);
  and (_22113_, _21839_, _20767_);
  and (_22114_, _21849_, _21605_);
  nor (_22115_, _22114_, _22113_);
  and (_22116_, _22115_, _22112_);
  and (_22117_, _22116_, _21057_);
  nor (_22118_, _22117_, _22109_);
  and (_22119_, _22118_, _21654_);
  nand (_22120_, _22119_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_22121_, _22119_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_22122_, _22121_, _22120_);
  and (_22123_, _21891_, _20792_);
  or (_22124_, _22123_, _21057_);
  and (_22125_, _21882_, _20767_);
  and (_22126_, _21887_, _21605_);
  or (_22127_, _22126_, _22125_);
  and (_22128_, _21877_, _20793_);
  or (_22129_, _22128_, _22127_);
  or (_22130_, _22129_, _22124_);
  and (_22131_, _21912_, _20792_);
  or (_22132_, _22131_, _20787_);
  and (_22133_, _21903_, _20767_);
  and (_22134_, _21908_, _21605_);
  and (_22135_, _21898_, _20793_);
  or (_22136_, _22135_, _22134_);
  or (_22137_, _22136_, _22133_);
  or (_22138_, _22137_, _22132_);
  and (_22139_, _22138_, _22130_);
  and (_22140_, _22139_, _21654_);
  and (_22141_, _22140_, _23790_);
  nor (_22142_, _22140_, _23790_);
  or (_22143_, _22142_, _22141_);
  or (_22144_, _22143_, _22122_);
  and (_22145_, _22002_, _20793_);
  and (_22146_, _21993_, _20792_);
  nor (_22147_, _22146_, _22145_);
  and (_22148_, _21998_, _21605_);
  and (_22149_, _21988_, _23844_);
  nor (_22150_, _22149_, _22148_);
  and (_22151_, _22150_, _22147_);
  nor (_22152_, _22151_, _20787_);
  and (_22153_, _21981_, _20793_);
  and (_22154_, _21972_, _20792_);
  nor (_22155_, _22154_, _22153_);
  and (_22156_, _21977_, _21605_);
  and (_22157_, _21967_, _20767_);
  nor (_22158_, _22157_, _22156_);
  and (_22159_, _22158_, _22155_);
  nor (_22160_, _22159_, _21057_);
  nor (_22161_, _22160_, _22152_);
  not (_22162_, _22161_);
  and (_22163_, _22162_, _21654_);
  nor (_22164_, _22163_, _23786_);
  and (_22165_, _22163_, _23786_);
  or (_22166_, _22165_, _22164_);
  and (_22167_, _21928_, _20792_);
  or (_22168_, _22167_, _21057_);
  and (_22169_, _21923_, _20767_);
  and (_22170_, _21933_, _21605_);
  or (_22171_, _22170_, _22169_);
  and (_22172_, _21937_, _20793_);
  or (_22173_, _22172_, _22171_);
  or (_22174_, _22173_, _22168_);
  and (_22175_, _21949_, _20792_);
  and (_22176_, _21958_, _20793_);
  and (_22177_, _21944_, _20767_);
  or (_22178_, _22177_, _22176_);
  or (_22179_, _22178_, _22175_);
  and (_22180_, _21954_, _21605_);
  or (_22181_, _22180_, _20787_);
  or (_22182_, _22181_, _22179_);
  and (_22183_, _22182_, _22174_);
  and (_22184_, _22183_, _21654_);
  nor (_22185_, _22184_, _23782_);
  and (_22186_, _22184_, _23782_);
  or (_22187_, _22186_, _22185_);
  or (_22188_, _22187_, _22166_);
  or (_22189_, _22188_, _22144_);
  or (_22190_, _22189_, _22101_);
  or (_22191_, _21177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_22192_, _21177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_22193_, _22192_, _22191_);
  nor (_22194_, _21216_, _23798_);
  and (_22195_, _21216_, _23798_);
  or (_22196_, _22195_, _22194_);
  or (_22197_, _22196_, _22193_);
  or (_22198_, _21095_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_22199_, _21095_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_22200_, _22199_, _22198_);
  and (_22201_, _21138_, _23806_);
  nor (_22202_, _21138_, _23806_);
  or (_22203_, _22202_, _22201_);
  or (_22204_, _22203_, _22200_);
  or (_22205_, _22204_, _22197_);
  or (_22206_, _21011_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_22207_, _21011_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22208_, _22207_, _22206_);
  and (_22209_, _21053_, _23816_);
  nor (_22210_, _21053_, _23816_);
  or (_22211_, _22210_, _22209_);
  or (_22212_, _22211_, _22208_);
  or (_22213_, _20887_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_22214_, _20887_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_22215_, _22214_, _22213_);
  and (_22216_, _20966_, _23824_);
  nor (_22217_, _20966_, _23824_);
  or (_22218_, _22217_, _22216_);
  or (_22219_, _22218_, _22215_);
  or (_22220_, _22219_, _22212_);
  or (_22221_, _22220_, _22205_);
  or (_22222_, _22221_, _22190_);
  not (_22223_, _22008_);
  not (_22224_, _21745_);
  and (_22225_, _21831_, _22224_);
  and (_22226_, _22225_, _21703_);
  and (_22227_, _22226_, _22223_);
  nor (_22228_, _21918_, _21874_);
  and (_22229_, _22228_, _22227_);
  and (_22230_, _22229_, _22222_);
  not (_22231_, _21964_);
  nor (_22232_, _21787_, _21702_);
  and (_22233_, _22232_, _21830_);
  and (_22234_, _22233_, _21745_);
  and (_22235_, _22234_, _22231_);
  not (_22236_, _21874_);
  and (_22237_, _21830_, _21703_);
  and (_22238_, _22237_, _21964_);
  and (_22239_, _22238_, _22008_);
  and (_22240_, _21830_, _22224_);
  and (_22241_, _22240_, _22232_);
  and (_22242_, _22008_, _21788_);
  and (_22243_, _22242_, _21964_);
  or (_22244_, _22243_, _22241_);
  or (_22245_, _22244_, _22226_);
  or (_22246_, _22245_, _22239_);
  and (_22247_, _22246_, _22236_);
  or (_22248_, _22247_, _22235_);
  and (_22249_, _22248_, _21918_);
  not (_22250_, _22007_);
  and (_22251_, _22250_, _21918_);
  and (_22252_, _22251_, _22225_);
  and (_22253_, _22007_, _21918_);
  and (_22254_, _22253_, _22234_);
  or (_22255_, _22254_, _22252_);
  or (_22256_, _22255_, _22227_);
  and (_22257_, _22256_, _21874_);
  not (_22258_, _21917_);
  and (_22259_, _22008_, _22258_);
  and (_22260_, _22259_, _22233_);
  and (_22261_, _22234_, _22223_);
  or (_22262_, _22261_, _22260_);
  and (_22263_, _22262_, _22236_);
  and (_22264_, _22223_, _21920_);
  and (_22265_, _22233_, _21964_);
  and (_22266_, _22265_, _22264_);
  and (_22267_, _22008_, _22225_);
  not (_22268_, _21788_);
  nor (_22269_, _21963_, _22268_);
  and (_22270_, _22237_, _22231_);
  or (_22271_, _22270_, _22269_);
  or (_22272_, _22271_, _22267_);
  and (_22273_, _22272_, _21920_);
  or (_22274_, _22273_, _22266_);
  or (_22275_, _22274_, _22263_);
  or (_22276_, _22275_, _22257_);
  or (_22277_, _22276_, _22249_);
  nor (_22278_, _20893_, _23816_);
  and (_22279_, _20893_, _23816_);
  or (_22280_, _22279_, _22278_);
  or (_22281_, _22280_, _21284_);
  nor (_22282_, _20781_, _23824_);
  and (_22283_, _20781_, _23824_);
  or (_22284_, _22283_, _22282_);
  or (_22285_, _22284_, _21269_);
  or (_22286_, _22285_, _22281_);
  or (_22287_, _20905_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_22288_, _20905_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_22289_, _22288_, _22287_);
  and (_22290_, _20928_, _23790_);
  nor (_22291_, _20794_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_22292_, _20794_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_22293_, _22292_, _22291_);
  nor (_22294_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_22295_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_22296_, _22295_, _22294_);
  not (_22297_, _22296_);
  and (_22298_, _22297_, _20768_);
  or (_22299_, _22298_, _22293_);
  and (_22300_, _20787_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_22301_, _20787_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22302_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_22303_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_22304_, _22303_, _22302_);
  nand (_22305_, _22304_, _21343_);
  nor (_22306_, _22297_, _20768_);
  or (_22307_, _22306_, _22305_);
  or (_22308_, _22307_, _22301_);
  or (_22309_, _22308_, _22300_);
  or (_22310_, _22309_, _22299_);
  nor (_22311_, _20928_, _23790_);
  or (_22312_, _22311_, _22310_);
  or (_22313_, _22312_, _22290_);
  or (_22314_, _20915_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_22315_, _20915_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_22316_, _22315_, _22314_);
  nor (_22317_, _20973_, _23786_);
  and (_22318_, _20973_, _23786_);
  or (_22319_, _22318_, _22317_);
  nor (_22320_, _20922_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_22321_, _20922_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_22322_, _22321_, _22320_);
  or (_22323_, _22322_, _22319_);
  or (_22324_, _22323_, _22316_);
  or (_22325_, _22324_, _22313_);
  nor (_22326_, _20912_, _23802_);
  and (_22327_, _20912_, _23802_);
  or (_22328_, _22327_, _22326_);
  or (_22329_, _22328_, _21299_);
  or (_22330_, _22329_, _22325_);
  or (_22331_, _22330_, _22289_);
  or (_22332_, _22331_, _22286_);
  and (_22333_, _22332_, _22277_);
  and (_22334_, _22260_, _22231_);
  and (_22335_, _22240_, _22268_);
  and (_22336_, _22008_, _22224_);
  or (_22337_, _22336_, _22242_);
  or (_22338_, _22337_, _22335_);
  and (_22339_, _22338_, _21918_);
  or (_22340_, _22339_, _22334_);
  and (_22341_, _22340_, _21874_);
  and (_22342_, _21745_, _21703_);
  and (_22343_, _22342_, _21831_);
  and (_22344_, _22241_, _22009_);
  or (_22345_, _22344_, _22343_);
  and (_22346_, _22345_, _21919_);
  and (_22347_, _22269_, _21918_);
  or (_22348_, _22237_, _21788_);
  and (_22349_, _22348_, _22228_);
  or (_22350_, _22349_, _22347_);
  nor (_22351_, _22008_, _21788_);
  and (_22352_, _22351_, _22238_);
  and (_22353_, _22250_, _21788_);
  and (_22354_, _22258_, _21964_);
  or (_22355_, _22354_, _22236_);
  and (_22356_, _22355_, _22353_);
  or (_22357_, _22356_, _22352_);
  or (_22358_, _22357_, _22350_);
  nand (_22359_, _22342_, _22268_);
  nor (_22360_, _22359_, _22236_);
  or (_22361_, _22360_, _22270_);
  and (_22362_, _22361_, _21918_);
  and (_22363_, _22009_, _21746_);
  and (_22364_, _22240_, _22223_);
  or (_22365_, _22364_, _22363_);
  and (_22366_, _22365_, _22228_);
  or (_22367_, _22366_, _22362_);
  or (_22368_, _22367_, _22358_);
  or (_22369_, _22368_, _22346_);
  or (_22370_, _22369_, _22341_);
  and (_22371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _23830_);
  and (_22372_, _20890_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22373_, _22372_, _22371_);
  and (_22374_, _22373_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_22375_, _22373_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_22376_, _23867_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_22377_, _20912_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22378_, _22377_, _22376_);
  nor (_22379_, _22378_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_22380_, _22378_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_22381_, _22380_, _22379_);
  or (_22382_, _22381_, _22375_);
  or (_22383_, _22382_, _22374_);
  and (_22384_, _20779_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_22385_, _20778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22386_, _22385_, _23885_);
  nor (_22387_, _22386_, _22384_);
  nand (_22388_, _22387_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_22389_, _22387_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_22390_, _22389_, _22388_);
  and (_22391_, _20768_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22392_, _22391_, _20771_);
  and (_22393_, _22392_, _20775_);
  and (_22394_, _22393_, _23878_);
  nor (_22395_, _22393_, _23878_);
  or (_22396_, _22395_, _22394_);
  nand (_22397_, _22396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_22398_, _22396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_22399_, _22398_, _22397_);
  not (_22400_, _22392_);
  nor (_22401_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_22402_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_22403_, _22402_, _22401_);
  nor (_22404_, _22403_, _22400_);
  and (_22405_, _22403_, _22400_);
  or (_22406_, _22405_, _22404_);
  nor (_22407_, _20796_, _23774_);
  and (_22408_, _20796_, _23774_);
  or (_22409_, _22408_, _22407_);
  or (_22410_, _22409_, _22406_);
  and (_22411_, _20919_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22412_, _22411_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22413_, _22412_, _22392_);
  nor (_22414_, _22413_, _23794_);
  nand (_22415_, _22304_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_22416_, _22304_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22417_, _22416_, _22415_);
  nor (_22418_, _22391_, _22297_);
  and (_22419_, _22391_, _22297_);
  or (_22420_, _22419_, _21343_);
  or (_22421_, _22420_, _22418_);
  or (_22422_, _22421_, _22417_);
  or (_22423_, _22422_, _22414_);
  or (_22424_, _22423_, _22410_);
  nor (_22425_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_22426_, _22425_, _22411_);
  nor (_22427_, _22426_, _20927_);
  and (_22428_, _22427_, _23790_);
  nor (_22429_, _22427_, _23790_);
  or (_22430_, _22429_, _22428_);
  or (_22431_, _22430_, _22424_);
  or (_22432_, _23851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_22433_, _20973_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22434_, _22433_, _22432_);
  nor (_22435_, _22434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_22436_, _20789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22437_, _20789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22438_, _22437_, _22436_);
  and (_22439_, _22413_, _23794_);
  or (_22440_, _22439_, _22438_);
  or (_22441_, _22440_, _22435_);
  or (_22442_, _22441_, _22431_);
  or (_22443_, _22442_, _22399_);
  not (_22444_, _20904_);
  nor (_22445_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22446_, _22392_, _20774_);
  nor (_22447_, _22446_, _22445_);
  and (_22448_, _22447_, _22444_);
  and (_22449_, _22448_, _23806_);
  nor (_22450_, _22448_, _23806_);
  or (_22451_, _22450_, _22449_);
  nor (_22452_, _22446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_22453_, _22446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_22454_, _22453_, _22452_);
  and (_22455_, _22454_, _23811_);
  nor (_22456_, _22454_, _23811_);
  and (_22457_, _22434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_22458_, _22457_, _22456_);
  or (_22459_, _22458_, _22455_);
  or (_22460_, _22459_, _22451_);
  or (_22461_, _22460_, _22443_);
  or (_22462_, _22461_, _22390_);
  nor (_22463_, _22384_, _09922_);
  and (_22464_, _22384_, _09922_);
  or (_22465_, _22464_, _22463_);
  nor (_22466_, _22465_, _20455_);
  and (_22467_, _22465_, _20455_);
  or (_22468_, _22467_, _22466_);
  or (_22469_, _22468_, _22462_);
  or (_22470_, _22469_, _22383_);
  and (_22471_, _22470_, _22370_);
  and (_22472_, _21964_, _21832_);
  or (_22473_, _22472_, _22235_);
  and (_22474_, _22473_, _22264_);
  and (_22475_, _22254_, _21963_);
  nand (_22476_, _22007_, _21963_);
  and (_22477_, _22476_, _21918_);
  and (_22478_, _22477_, _22343_);
  or (_22479_, _22478_, _22475_);
  and (_22480_, _22479_, _22236_);
  or (_22481_, _22480_, _22474_);
  and (_22482_, _21545_, _20771_);
  and (_22483_, _22482_, _20774_);
  and (_22484_, _22483_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_22485_, _22484_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_22486_, _22485_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_22487_, _22486_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_22488_, _22487_, _21265_);
  nor (_22489_, _22487_, _21265_);
  nor (_22490_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22491_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_22492_, _22491_, _22490_);
  nor (_22493_, _22492_, _22485_);
  and (_22494_, _22492_, _22485_);
  and (_22495_, _22482_, _20773_);
  and (_22496_, _22482_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22497_, _22496_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_22498_, _22497_, _22495_);
  nor (_22499_, _22498_, _23802_);
  and (_22500_, _22498_, _23802_);
  or (_22501_, _22500_, _22499_);
  and (_22502_, _21545_, _20770_);
  and (_22503_, _21545_, _20769_);
  nor (_22504_, _22503_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_22505_, _22504_, _22502_);
  nor (_22506_, _22505_, _23790_);
  or (_22507_, _22506_, _22501_);
  or (_22508_, _22507_, _22494_);
  or (_22509_, _22508_, _22493_);
  or (_22510_, _22509_, _22489_);
  or (_22511_, _22510_, _22488_);
  nor (_22512_, _22486_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_22513_, _22512_, _22487_);
  nor (_22514_, _22513_, _23824_);
  and (_22515_, _22513_, _23824_);
  nor (_22516_, _22484_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_22517_, _22516_, _22485_);
  and (_22518_, _22517_, _23816_);
  nor (_22519_, _22517_, _23816_);
  or (_22520_, _22519_, _22518_);
  nor (_22521_, _22502_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22522_, _22521_, _22482_);
  and (_22523_, _22522_, _23794_);
  nor (_22524_, _22495_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_22525_, _22524_, _22483_);
  nor (_22526_, _22525_, _23806_);
  nor (_22527_, _22522_, _23794_);
  or (_22528_, _22527_, _22526_);
  or (_22529_, _22528_, _22523_);
  and (_22530_, _22505_, _23790_);
  or (_22531_, _21547_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_22532_, _21547_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22533_, _22532_, _22531_);
  or (_22534_, _22296_, _21545_);
  nand (_22535_, _22296_, _21545_);
  and (_22536_, _22535_, _22534_);
  nand (_22537_, _22417_, _21344_);
  and (_22538_, _21543_, _23774_);
  nor (_22539_, _21543_, _23774_);
  or (_22540_, _22539_, _22538_);
  or (_22541_, _22540_, _22537_);
  or (_22542_, _22541_, _22536_);
  or (_22543_, _22542_, _22533_);
  or (_22544_, _22543_, _22530_);
  nor (_22545_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_22546_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_22547_, _22546_, _22545_);
  nor (_22548_, _22547_, _22483_);
  and (_22549_, _22547_, _22483_);
  or (_22550_, _22549_, _22548_);
  or (_22551_, _22550_, _22544_);
  and (_22552_, _22525_, _23806_);
  nor (_22553_, _22482_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22554_, _22553_, _22496_);
  nor (_22555_, _22554_, _23798_);
  and (_22556_, _21545_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_22557_, _22556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_22558_, _22557_, _22503_);
  and (_22559_, _22558_, _23786_);
  or (_22560_, _22559_, _22555_);
  and (_22561_, _22554_, _23798_);
  nor (_22562_, _22558_, _23786_);
  or (_22563_, _22562_, _22561_);
  or (_22564_, _22563_, _22560_);
  or (_22565_, _22564_, _22552_);
  or (_22566_, _22565_, _22551_);
  or (_22567_, _22566_, _22529_);
  or (_22568_, _22567_, _22520_);
  or (_22569_, _22568_, _22515_);
  or (_22570_, _22569_, _22514_);
  or (_22571_, _22570_, _22511_);
  and (_22572_, _22571_, _22481_);
  or (_22573_, _22572_, _22471_);
  or (_22574_, _22573_, _22333_);
  or (_22575_, _22574_, _22230_);
  and (_22576_, _22575_, _21661_);
  and (_22577_, _22008_, _23798_);
  nor (_22578_, _22008_, _23798_);
  or (_22579_, _22578_, _22577_);
  nor (_22580_, _21918_, _23802_);
  and (_22581_, _21918_, _23802_);
  or (_22582_, _22581_, _22580_);
  or (_22583_, _22582_, _22579_);
  nor (_22584_, _21874_, _23806_);
  and (_22585_, _21874_, _23806_);
  or (_22586_, _22585_, _22584_);
  or (_22587_, _22586_, _21299_);
  or (_22588_, _22587_, _22583_);
  or (_22589_, _22588_, _22286_);
  or (_22590_, _21177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_22591_, _21177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22592_, _22591_, _22590_);
  and (_22593_, _21216_, _23765_);
  nor (_22594_, _21216_, _23765_);
  or (_22595_, _22594_, _22593_);
  or (_22596_, _22595_, _22592_);
  or (_22597_, _21095_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_22598_, _21095_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22599_, _22598_, _22597_);
  nor (_22600_, _21138_, _23774_);
  and (_22601_, _21138_, _23774_);
  or (_22602_, _22601_, _22600_);
  or (_22603_, _22602_, _22599_);
  or (_22604_, _22603_, _22596_);
  or (_22605_, _21011_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_22606_, _21011_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_22607_, _22606_, _22605_);
  nor (_22608_, _21053_, _23782_);
  and (_22609_, _21053_, _23782_);
  or (_22610_, _22609_, _22608_);
  or (_22611_, _22610_, _22607_);
  nor (_22612_, _20887_, _23794_);
  and (_22613_, _20887_, _23794_);
  or (_22614_, _22613_, _22612_);
  and (_22615_, _20966_, _23790_);
  nor (_22616_, _20966_, _23790_);
  or (_22617_, _22616_, _22615_);
  or (_22618_, _22617_, _22614_);
  or (_22619_, _22618_, _22611_);
  or (_22620_, _22619_, _22604_);
  or (_22621_, _22620_, _22589_);
  nor (_22622_, _22224_, _21702_);
  and (_22623_, _22622_, _21831_);
  and (_22624_, _22623_, _21661_);
  and (_22625_, _22624_, _22621_);
  or (_22626_, _22625_, _22576_);
  or (property_invalid, _22626_, _22013_);
  and (_22627_, _16219_, _23715_);
  and (_22628_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or (_12142_, _22628_, _22627_);
  and (_22629_, _21655_, first_instr);
  or (_00000_, _22629_, rst);
  and (_22630_, _16219_, _23693_);
  and (_22631_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or (_12148_, _22631_, _22630_);
  and (_22632_, _02798_, _23900_);
  and (_22633_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_12201_, _22633_, _22632_);
  and (_22634_, _16219_, _24027_);
  and (_22635_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or (_12203_, _22635_, _22634_);
  and (_22636_, _16219_, _23983_);
  and (_22637_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or (_12216_, _22637_, _22636_);
  and (_22638_, _10547_, _23693_);
  and (_22639_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or (_27009_, _22639_, _22638_);
  and (_22640_, _10514_, _23920_);
  and (_22641_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_12220_, _22641_, _22640_);
  and (_22642_, _10514_, _23751_);
  and (_22643_, _10516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_26977_, _22643_, _22642_);
  and (_22644_, _02350_, _24027_);
  and (_22645_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_12259_, _22645_, _22644_);
  and (_22646_, _10547_, _23715_);
  and (_22647_, _10549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or (_12261_, _22647_, _22646_);
  and (_22648_, _15246_, _24053_);
  and (_22649_, _15248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_12269_, _22649_, _22648_);
  and (_22650_, _02350_, _23983_);
  and (_22651_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_12273_, _22651_, _22650_);
  and (_22652_, _10536_, _23900_);
  and (_22653_, _10538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or (_12278_, _22653_, _22652_);
  and (_22654_, _04767_, _23983_);
  and (_22655_, _04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_12285_, _22655_, _22654_);
  and (_22656_, _10695_, _23920_);
  and (_22657_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_12297_, _22657_, _22656_);
  and (_22658_, _01936_, _23900_);
  and (_22659_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_12299_, _22659_, _22658_);
  and (_22660_, _10695_, _23751_);
  and (_22661_, _10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_27029_, _22661_, _22660_);
  and (_22662_, _01936_, _23715_);
  and (_22663_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_12313_, _22663_, _22662_);
  and (_22664_, _02326_, _23983_);
  and (_22665_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or (_12319_, _22665_, _22664_);
  and (_22666_, _01936_, _23920_);
  and (_22667_, _01938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_12326_, _22667_, _22666_);
  and (_22668_, _02798_, _24053_);
  and (_22669_, _02800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_12338_, _22669_, _22668_);
  and (_22670_, _25482_, _23920_);
  and (_22671_, _25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_12340_, _22671_, _22670_);
  and (_22672_, _16219_, _24053_);
  and (_22673_, _16221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or (_12342_, _22673_, _22672_);
  and (_22674_, _25198_, _23751_);
  and (_22675_, _25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or (_12346_, _22675_, _22674_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _26814_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _26814_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _26814_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _26814_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _26814_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _26814_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _26814_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _26814_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _26830_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _26812_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _26812_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _26812_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _26812_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _26812_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _26812_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _26812_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _26812_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _26812_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _26812_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _26812_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _26812_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _26812_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _26812_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _26812_[15]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _26821_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _26821_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _26821_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _26821_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _26821_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _26821_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _26821_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _26821_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _26822_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _26822_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _26822_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _26822_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _26822_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _26822_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _26822_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _26822_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _26823_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _26823_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _26823_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _26823_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _26823_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _26823_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _26823_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _26823_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _26824_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _26824_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _26824_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _26813_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _26824_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _26824_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _26824_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _26824_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _26825_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _26825_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _26825_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _26825_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _26825_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _26825_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _26825_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _26825_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _26826_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _26826_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _26826_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _26826_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _26826_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _26826_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _26826_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _26826_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _26827_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _26827_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _26827_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _26827_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _26827_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _26827_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _26827_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _26827_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _26828_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _26828_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _26828_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _26828_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _26828_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _26828_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _26828_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _26828_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _26829_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _26829_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _26829_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _26829_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _26829_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _26829_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _26829_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _26829_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _26815_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _26815_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _26815_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _26815_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _26815_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _26815_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _26815_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _26815_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _26816_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _26816_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _26816_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _26816_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _26816_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _26816_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _26816_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _26816_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _26817_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _26817_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _26817_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _26817_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _26817_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _26817_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _26817_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _26817_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _26818_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _26818_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _26818_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _26818_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _26818_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _26818_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _26818_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _26818_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _26819_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _26819_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _26819_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _26819_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _26819_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _26819_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _26819_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _26819_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _26820_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _26820_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _26820_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _26820_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _26820_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _26820_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _26820_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _26820_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _05495_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _05488_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _05493_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _05490_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _05503_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _11453_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _05531_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00732_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _05548_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _05542_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _05545_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _05565_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _05558_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _05562_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _05572_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _11359_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11716_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _11199_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11659_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11639_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11641_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11661_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11670_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11643_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11645_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _11663_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11647_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11649_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11665_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11674_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11653_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11655_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _26831_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _26831_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _26831_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _26831_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _26831_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _26831_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _26831_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _26831_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _26858_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _26858_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _26858_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _26858_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _26858_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _26858_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _26858_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _26858_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _26868_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _26868_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _26868_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _26868_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _26868_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _26868_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _26868_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _26868_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _26838_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _26838_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _26839_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _26839_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _26839_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _26840_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _26840_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _26840_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _26841_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _26841_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _26842_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _26842_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _26842_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _26842_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _26843_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _26843_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _26844_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _26832_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _26832_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _26832_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _26833_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _26833_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _26833_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _26834_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _26834_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _26835_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _26835_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _26835_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _26835_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _26835_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _26835_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _26835_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _26835_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _26836_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _26837_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _26837_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _26883_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _26845_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _26845_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _26845_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _26845_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _26845_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _26845_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _26845_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _26845_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _26846_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _26846_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _26846_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _26846_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _26846_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _26846_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _26846_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _26846_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _26847_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _26847_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _26847_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _26847_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _26847_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _26847_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _26847_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _26847_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _26848_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _26848_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _26848_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _26848_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _26848_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _26848_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _26848_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _26848_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _26849_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _26849_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _26849_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _26849_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _26849_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _26849_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _26849_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _26849_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _26850_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _26850_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _26850_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _26850_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _26850_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _26850_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _26850_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _26850_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _26851_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _26851_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _26851_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _26851_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _26851_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _26851_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _26851_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _26851_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _26852_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _26852_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _26852_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _26852_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _26852_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _26852_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _26852_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _26852_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _26856_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _26856_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _26856_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _26856_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _26856_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _26853_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _26853_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _26853_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _26853_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _26853_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _26853_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _26853_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _26853_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _26853_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _26853_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _26853_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _26853_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _26853_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _26853_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _26853_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _26853_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _26854_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26854_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26854_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _26854_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _26854_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _26854_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _26854_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _26854_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _26854_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _26854_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _26854_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26854_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _26854_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _26854_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _26854_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _26854_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _26874_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _26874_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _26874_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _26874_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _26874_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _26874_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _26874_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _26874_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _26874_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _26874_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _26874_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _26874_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _26874_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _26874_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _26874_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _26874_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _26874_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _26874_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _26874_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _26874_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _26874_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _26874_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _26874_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _26874_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _26874_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _26874_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _26874_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _26874_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _26874_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _26874_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _26874_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _26874_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _26855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _26857_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _26857_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _26857_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _26857_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _26857_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _26857_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _26857_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _26857_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _26859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _26860_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _26861_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _26861_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _26861_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _26861_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _26861_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _26861_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _26861_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _26861_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _26861_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _26861_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _26861_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _26861_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _26861_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _26861_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _26861_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _26861_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _26862_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _26862_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _26862_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _26862_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _26862_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _26862_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _26862_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _26862_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _26862_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _26862_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _26862_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _26862_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _26862_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _26862_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _26862_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _26862_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _26863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _26865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _26864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _26866_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _26866_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _26866_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _26866_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _26866_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _26866_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _26866_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _26866_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _26867_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26867_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _26867_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _26869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _26870_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _26870_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _26870_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _26870_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _26870_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _26870_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _26870_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _26870_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _26871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _26872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _26873_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _26873_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _26873_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _26873_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _26875_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _26875_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _26875_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _26875_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _26875_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _26875_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _26875_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _26875_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _26875_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _26875_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _26875_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _26875_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _26875_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _26875_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _26875_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _26875_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _26875_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _26875_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _26875_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _26875_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _26875_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _26875_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _26875_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _26875_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _26875_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _26875_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _26875_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _26875_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _26875_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _26875_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _26875_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _26875_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _26876_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _26877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _26878_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _26879_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _26879_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _26879_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _26879_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _26880_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _26881_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26882_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26882_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26882_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26882_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26882_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26882_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26882_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _26882_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _26884_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _26884_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _26884_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _04737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _05794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _05777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _26943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _05861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _05857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _05845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _08554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _13221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _11829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _26934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _26935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _26936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _05901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _09187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _26937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _26917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _26918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _26919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _26920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _26921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _26922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _22680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _11727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _22699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _26899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _22708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _22707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _26900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _22684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _22683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _22690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _26957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _06040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _04531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _06092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _06083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _09521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _00142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _22730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _22709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _27317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _27318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _22714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _22713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _22711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _27319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _27320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _14057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _11170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _27156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _15507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _15748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _11145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _15790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _27157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _15283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _27136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _27137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _15465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _13813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _11176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _13864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _13976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _11154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _14974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _27120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _15046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _15235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _11149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _27121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _15250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _09268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _10216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _09380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _09369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _09045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _08991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _08989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _10231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _10621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _07595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _09473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _27216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _09633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _09594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _08039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _09235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _27213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _11538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _11500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _10157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _07751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _10281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _27214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _27215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _09895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _07805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _22737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _27212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _10143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _07667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _10135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _11324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _09848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _03266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _01943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _07673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _01708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _09859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _26029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _27211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _01416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _27209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _01782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _01677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _27210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _22858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _24794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _23227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _10126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _00364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _01039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _00705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _07682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _09812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _26791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _07679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _07395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _06270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _10116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _27205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _27206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _27207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _23556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _27208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _09646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _09484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _10114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _11541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _27202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _07765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _03505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _03317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _08812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _07643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _05506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _27201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _23457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _11472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _11109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _10100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _08707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _27199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _10087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _09073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _09083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _09085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _10097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _27200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _10676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _27311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _10680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _09171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _10694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _27312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _09165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _27313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _27309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _27310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _09013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _10633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _09173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _10653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _09010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _10660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _09025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _09265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _10393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _09022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _10423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _10535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _09019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _10555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _10339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _27308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _09280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _10344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _10355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _09034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _10373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _09032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _10232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _10256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _09104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _09293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _10262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _10301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _27307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _10325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _09231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _10163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _10179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _09110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _09283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _10185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _10228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _09108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _09157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _09864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _09155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _09883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _09251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _09296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _10133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _10159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _27304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _09114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _09309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _09326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _09305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _09162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _27305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _27306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _02490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _09433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _10944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _07678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _27273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _07738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _10954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _27274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _27298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _27299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _10068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _27300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _09118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _10093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _10098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _10104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _10627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _07441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _26893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _26894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _10885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _07266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _10893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _07264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _10401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _07350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _09917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _07353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _10493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _10571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _07341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _26892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _10791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _10798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _26890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _10800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _07277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _10804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _26891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _09920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _10750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _07403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _10763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _07288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _10767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _10786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _10789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _07282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _25935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _09311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _06371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _02308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _26910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _22925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _06662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _26911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _26905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _26906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _26907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _26908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _26909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _09474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _06652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _06374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _07206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _26902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _07363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _11178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _11187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _26903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _07176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _26904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _05305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _02169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _05389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _27160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _05004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _05000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _02180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _05171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _05905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _24587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _05608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _05539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _05703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _05690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _24584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _05333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _02131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _25286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _05852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _05843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _27159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _05789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _05945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _05942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _27158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _06604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _24600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _06064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _06046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _06038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _06129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _06166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _06774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _06766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _02108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _25296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _06556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _06550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _06538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _06650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _02102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _06898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _27153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _27154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _02095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _06673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _27155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _06761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _07023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _07039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _07031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _24614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _25553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _06854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _06852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _27152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _27149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _27150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _07099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _07227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _07163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _27151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _06971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _06965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _07337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _07299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _07292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _02065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _07374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _27147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _02061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _27148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _02042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _27146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _07480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _07477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _07448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _02057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _07544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _07533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _07767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _08055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _27143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _08036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _27144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _07603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _27145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _07716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _03991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _10890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _02078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _27271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _10917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _27272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _02837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _02787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _09834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _24656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _08406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _08403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _27141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _08934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _27142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _25366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _09313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _09291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _09387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _24780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _25616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _09249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _09167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _27140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _05767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _24786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _00520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _27138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _04294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _24783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _00418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _27139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _24792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _10559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _10332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _00379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _10783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _00375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _25629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _00490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _01989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _25371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _27132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _07664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _09015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _27133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _27134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _27135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _10492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _27131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _24692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _10037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _10014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _01993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _10236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _10194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _10778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _01973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _10912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _27130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _24701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _10336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _10348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _01985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _24713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _11022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _27129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _10998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _11159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _11130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _01956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _10762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _11836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _01930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _27126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _27127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _27128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _01950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _11373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _11404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _12338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _24734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _11864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _27125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _12201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _01912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _25391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _11617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _05614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _09208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _23042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _10773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _01884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _25669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _12259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _12273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _12621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _27267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _05231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _27268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _27269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _27270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _04331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _04257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _08649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _27124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _07596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _07233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _11076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _01853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _25498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _01968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _22689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _00936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _23382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _24760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _25598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _09623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _09591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _01845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _10826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _27259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _27260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _11269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _11227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _10991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _09808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _27261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _10506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _10419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _10313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _27265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _10993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _27266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _11983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _11020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _27122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _11861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _24771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _27123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _02804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _10769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _09777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _01763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _05279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _02830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _03129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _09245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _11570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _25130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _13792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _24776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _02678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _05195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _27118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _27119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _02673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _05256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _02834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _05272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _27254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _09539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _27255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _07695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _11680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _11667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _10735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _11851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _10725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _08817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _08963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _10744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _27256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _27257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _10741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _27258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _02987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _24194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _10664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _07700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _22736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _10679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _22722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _22720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _27248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _27249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _27250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _08729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _27251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _00105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _00164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _07540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _11621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _27061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _11389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _24327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _24334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _11637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _27062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _11633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _06185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _27246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _22729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _27247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _26159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _22733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _07546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _22686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _24645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _26885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _11619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _24496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _24493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _24491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _24465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _24547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _11678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _23684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _27220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _27221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _23477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _23473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _23592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _23574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _23916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _23908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _23720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _24007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _24001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _23956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _27203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _27204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _24208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _24291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _11651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _27177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _24075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _24070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _11657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _27178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _22769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _27284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _22936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _22921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _27285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _27286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _27287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _11692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _23049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _23027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _23141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _23203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _27262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _11689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _27263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _27264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _27236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _23329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _23339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _23334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _27237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _27238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _23410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _27239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _22767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _27301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _22715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _22721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _22716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _22735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _27302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _27303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _04976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _05095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _02692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _02969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _05121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _02690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _05147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _27117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _02854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _04013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _04132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _02703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _02972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _04199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _04956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _02698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _02859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _03187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _03245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _02713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _27116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _03193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _03254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _04011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _01593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _02868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _01623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _01649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _27114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _02979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _27115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _02965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _02743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _01398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _02875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _01507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _01540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _02729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _27113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _01576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _01329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _02757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _01334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _02878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _01354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _01392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _02747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _02993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _22698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _02812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _07586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _27111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _07608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _04693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _27112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _03045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _01277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _02881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _03177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _22911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _02824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _22718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _02946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _27110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _02774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _27103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _02887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _01184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _02770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _01190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _27104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _01257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _23829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _00919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _02784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _03041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _00944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _02781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _00954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _02890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _02915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _27101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _23762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _02793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _27102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _23807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _23826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _02788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _05446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _05640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _26115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _27099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _05551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _26085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _03581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _27100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _05469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _25770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _05360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _25772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _25760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _26141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _26015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _26020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _05612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _27096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _05600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _05373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _27097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _27098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _05497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _05465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _04958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _03876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _27095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _04978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _03866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _04980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _04997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _03850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _04140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _04885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _04894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _03899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _04212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _04898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _27094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _04933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _03947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _27092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _04831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _03932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _27093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _04145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _04855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _04878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _27089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _04764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _03969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _27090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _04776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _27091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _04780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _04153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _04687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _04005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _04701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _03995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _04703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _04157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _27088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _04739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _04597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _04620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _04026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _04626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _04161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _04638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _04664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _04675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _04122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _04314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _27085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _04112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _27086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _04108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _27087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _04245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _27083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _04540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _04562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _27084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _04034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _04299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _04309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _04119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _27077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _04239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _27078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _27079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _04068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _27080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _27081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _27082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _27071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _27072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _27073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _27074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _04084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _27075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _04181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _27076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _27068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _26251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _26248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _26233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _05522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _26011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _27069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _27070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _27064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _26280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _27065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _26316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _27066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _27067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _05461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _26194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _25679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _25793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _25788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _25783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _05382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _00445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _00437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _26299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _25819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _25834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _05378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _27063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _25950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _25927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _05370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _25699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _02948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _27060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _03472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _03464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _03439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _03579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _03545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _05603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _03144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _27059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _03291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _03281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _00779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _00537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _00525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _02955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _04987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _11331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _05315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _27057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _05386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _05366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _27058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _03577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _10712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _10704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _10688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _27054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _07012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _27055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _04990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _27056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _03591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _27051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _27052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _27053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _10875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _10861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _10529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _10369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _27046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _27047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _27048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _11124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _11061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _27049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _27050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _11842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _27044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _06973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _23491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _23438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _04909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _27045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _04936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _22719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _03722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _27043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _26000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _04907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _01690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _01696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _04903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _10924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _07061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _03248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _02294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _02374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _02299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _04226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _03744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _03409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _09142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _09137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _03257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _27041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _05290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _05259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _27042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _07335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _27038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _27039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _09464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _09447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _04862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _08886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _08938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _04882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _09607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _09571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _10557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _10530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _27037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _03264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _09275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _09363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _23018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _03272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _10855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _27036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _11522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _11497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _11492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _03269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _27035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _04603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _03542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _04804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _19899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _19933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _22738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _16505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _09092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _07606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _04791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _10810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _04784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _03726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _23358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _22771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _09149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _09970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _10027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _09147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _10034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _27297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _10041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _09241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _10947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _27296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _10935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _04897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _09902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _09935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _09151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _09940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _11039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _27294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _11018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _11000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _10903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _10895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _27295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _02537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _27292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _10700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _10715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _10732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _08116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _10739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _27293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _11030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _10638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _08125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _08925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _10645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _10665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _08123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _27291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _10691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _10508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _10572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _08132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _08927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _10582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _10607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _08129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _10626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _10368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _10386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _08136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _27289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _08973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _10389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _10468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _27290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _08420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _10321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _10340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _08142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _08930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _10346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _10359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _08139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _10197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _08150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _10217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _27288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _10258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _08148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _10264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _10302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _09874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _27283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _09885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _08920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _10142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _10161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _08154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _10169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _10124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _27281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _08398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _09781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _09307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _08399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _27282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _09846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _08912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _10076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _10095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _08162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _27280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _08160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _10105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _10121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _10029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _08169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _10039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _27279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _10050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _08914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _10063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _08166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _10929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _27278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _09909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _09938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _08172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _09943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _09964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _08917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _08689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _10949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _27275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _27276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _27277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _07186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _06914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _06887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _01828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _01710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _10299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _07719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _25073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _23857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _23517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _00516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _10066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _20019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _27197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _00125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _10073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _22726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _10072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _27198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _10287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _02635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _03348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _02961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _10269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _01263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _01581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _01706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _08604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _07654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _08790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _10056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _09009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _07649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _08051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _22688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _27218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _06483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _27219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _06311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _10254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _02459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _02449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _02433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _27194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _09979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _07579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _10845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _27195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _10016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _07784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _27196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _09134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _07182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _27217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _07070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _07045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _08884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _07503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _04713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _27191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _09966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _27192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _09962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _27193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _24311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _24260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _10011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _22677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _27190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _09933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _07801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _06089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _09955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _06668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _06647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _27185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _27186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _11078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _27187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _27188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _27189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _14209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _01899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _27179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _11090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _27180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _11088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _27181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _27182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _27183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _27184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _11103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _27172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _11190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _27173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _27174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _11095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _27175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _27176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _18277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _11113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _27170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _11192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _18497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _20227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _11107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _27171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _17511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _27167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _17562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _11194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _17583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _17655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _27168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _27169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _27164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _16112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _11132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _27165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _27166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _16999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _17181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _11121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _11141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _27162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _15881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _15952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _11138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _16003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _11134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _27163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _27008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _05244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _27009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _12261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _05735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _27010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _05642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _05638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _27105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _14652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _14743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _27106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _27107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _27108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _11156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _27109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _10898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _27315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _02563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _10951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _10938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _10956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _27316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _02600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _24695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _27016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _24499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _24558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _24552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _27017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _03693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _24409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _03536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _24306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _27018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _27019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _03691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _27020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _07594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _27021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _24256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _26984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _24073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _26985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _24125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _26986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _26987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _26988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _07565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _07572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _07611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _07657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _07641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _07613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _06280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _06537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _07475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _07468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _06796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _07508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _07514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _07510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _07368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _07707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _07696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _07692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _07688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _07763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _07748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _07744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _07742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _11417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _11572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _11611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _06749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _06465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _05848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _06624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _06366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _10737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _27314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _11028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _11007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _11036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _11011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _11014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _05277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _27252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _09659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _10701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _11480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _27253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _07535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _00629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _12319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _25724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _27244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _07499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _25070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _23838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _23834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _27245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _07702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _27241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _01182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _27242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _01165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _01377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _01337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _27243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _10623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _05568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _10540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _08156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _08050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _10518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _05192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _05211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _05200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _05066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _04974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _10587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _01402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _27240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _10608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _02398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _02342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _05331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _05302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _10560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _07705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _03519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _04003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _03822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _10596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _27231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _10380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _11173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _07562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _27232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _27233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _10388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _10858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _10391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _09708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _09689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _09675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _10408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _10362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _27235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _07710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _07559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _08029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _08110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _10668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _10659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _10613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _10753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _27234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _27225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _27226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _27227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _27228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _27229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _12340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _11406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _27230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _07662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _07575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _11849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _11845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _11875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _11868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _07570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _11004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _05472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _12346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _14118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _14469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _11166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _14520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _11163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _14591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _05237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _05203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _05427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _05440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _12278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _05420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _05476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _05483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _27028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _27029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _05666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _05669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _27030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _12297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _05528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _05520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _05583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _27040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _05560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _12313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _12299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _12326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _22732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _05216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _05297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _26977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _26978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _26979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _05342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _12220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _26980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _05158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _08685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _08702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _03284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _10460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _06875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _23773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _09200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _27034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _22731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _05292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _00421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _27031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _09190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _03286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _03729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _08617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _08577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _08593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _22724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _22725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _22727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _27032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _27033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _08854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _01424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _25563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _25675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _08667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _08663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _23369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _04720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _07161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _10835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _22734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _03320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _13520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _06078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _07332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _22772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _06193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _04696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _11866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _10284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _22728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _23674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _02442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _22687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _03304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _03308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _01561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _07344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _04984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _02511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _20200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _25555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _24430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _08950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _03081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _02806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _27027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _03328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _09128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _09828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _08412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _27025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _25009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _23070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _27026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _00032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _26760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _09923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _22697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _03965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _03910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _27023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _03372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _27024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _00968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _02107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _01850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _24766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _03553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _25602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _25588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _27014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _27015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _03575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _24607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _08895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _04951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _27022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _04613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _06564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _06151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _03381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _02819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _11248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _04575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _12219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _12004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _04567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _27007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _09661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _04584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _27011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _10593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _04580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _03663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _27012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _27013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _25377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _24739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _17634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _03437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _12910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _12759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _04559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _13885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _13601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _03434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _22679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _22678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _22676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _27005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _15769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _15486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _15265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _27006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _03457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _22681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _22682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _22691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _27001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _27002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _27003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _27004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _22777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _22770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _22934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _03475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _22761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _26995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _22766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _03470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _22712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _22710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _26996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _22717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _26997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _26998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _26999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _27000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _26992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _26993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _23486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _03480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _23113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _23072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _23320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _26994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _26972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _26973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _26974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _05712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _26975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _05707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _26976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _05954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _23947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _23962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _23619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _26989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _23646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _26990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _23430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _26991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _05701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _26981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _26982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _05695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _26983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _05940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _00510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _24187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _05975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _04307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _05729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _26969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _05964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _26970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _26971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _05722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _05753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _06099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _04276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _05750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _04279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _05981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _26968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _04302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _04217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _05764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _06101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _04221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _26967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _05760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _04248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _05757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _06002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _26964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _04168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _05774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _04184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _26965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _26966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _04193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _26963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _06009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _04115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _04126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _05800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _06110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _04129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _04148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _05928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _03863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _03868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _26961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _26962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _03799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _06176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _04103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _05865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _04037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _26959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _04043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _04048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _05855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _06119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _04079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _26960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _04086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _04099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _05839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _06114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _03833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _05931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _03966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _05879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _03972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _06056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _03984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _04009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _26958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _06125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _08026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _03889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _05899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _03901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _06067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _03915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _03937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _05884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _03678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _06902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _26954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _26955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _06899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _26956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _07154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _07153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _26951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _04946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _04972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _06879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _04743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _04732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _04723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _06884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _04798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _26952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _04552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _04522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _26953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _04659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _04633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _06888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _05106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _05078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _05060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _06877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _05152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _05175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _06211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _26950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _05554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _06218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _05299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _05284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _05268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _05379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _05353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _05348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _26947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _05717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _06857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _05525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _26948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _26949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _06866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _05574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _05986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _05972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _06050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _06075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _06062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _06848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _05829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _26945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _05875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _05903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _05892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _26946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _06523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _05654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _05649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _06859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _06127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _06161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _06153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _06526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _06520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _06481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _06248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _26944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _06731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _26942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _06528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _06565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _06559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _06640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _06638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _06622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _06843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _26941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _06837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _06841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _06693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _06683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _06677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _06744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _26940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _06267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _06535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _07017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _06992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _06978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _07035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _06829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _06893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _06890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _06839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _06948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _06835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _06433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _06793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _06787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _07231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _07310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _07306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _07295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _06806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _07065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _07074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _06826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _07360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _26938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _07407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _07405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _26939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _06436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _07229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _07243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _08414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _06784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _08024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _07803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _06790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _08041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _08047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _08044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _06781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _09131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _09169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _06780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _08394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _08392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _08389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _08386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _09317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _09321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _09319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _09951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _09911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _26933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _09029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _08979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _06759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _10630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _10618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _06763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _26928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _26929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _26930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _26931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _10296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _10374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _10371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _10357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _06293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _10091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _26932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _10201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _27161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _25549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _25722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _04810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _04789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _04781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _04930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _04910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _06757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _11136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _11126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _11099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _06460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _10870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _10863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _10971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _11197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _26925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _26926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _11363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _11336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _26927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _11065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _11043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _06382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _06634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _05438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _26923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _03981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _04297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _04290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _26924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _02852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _02808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _06375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _06895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _06660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _06620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _07248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _06601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _06333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _11833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _11724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _11685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _11855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _11853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _06746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _11469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _12342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _06734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _12148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _12142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _12082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _06742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _12203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _12216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _06697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _26915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _05581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _26916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _06701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _06477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _22685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _10156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _02002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _06340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _00033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _06729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _10873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _06708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _06546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _12285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _06685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _11721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _11566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _06695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _02990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _06346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _10614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _26914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _06682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _26913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _06680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _06480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _22693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _22723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _06687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _10397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _12269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _06665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _26912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _07591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _06671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _10832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _10867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _06359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _11045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _07371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _11086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _11097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _07224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _07446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _11111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _26901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _11002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _07375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _11009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _11024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _07236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _07450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _07493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _11032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _07252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _10960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _07387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _10968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _10983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _07246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _07454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _10988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _26888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _10686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _26889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _07473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _10696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _10707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _07409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _10748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _27222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _25839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _07577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _27223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _22706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _16477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _27224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _22768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _07259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _26895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _26896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _26897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _07256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _26898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _10941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _07486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _11058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _05451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _05580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _10979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _05397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _10981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _10640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _26887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _02665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _10878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _02706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _26886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _10925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _05034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _10927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _04829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _27321_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _06407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _10234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _27321_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _08982_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _27322_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _27323_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _27323_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _27323_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _27323_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _27324_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _27325_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _27326_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _27326_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _27326_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _27326_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _27326_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _27326_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _27326_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _27326_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10438_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10484_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10350_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _07452_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _07460_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _07458_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _07466_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _07464_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _07462_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _07470_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _10165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _10021_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _10147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _10082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _10048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _10151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _10149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _09919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09993_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _10182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _10167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _10023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _10146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _10119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _10089_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _09928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _05970_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _22701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _12309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _12420_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _12399_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _12358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _12333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _05984_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _11627_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _11357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _11462_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _11499_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _22703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _11355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _11871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _22702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _11365_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _10854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _11290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _11430_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _11415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _11440_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _11423_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _10467_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _10451_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _10435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _11456_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _09879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _09763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _09861_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _09826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _09790_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _22704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _10212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _11450_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _09351_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _09331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _09302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _09255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _22705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _09573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _09536_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _11444_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _06272_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _23500_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _15135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _14995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _15120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _15106_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _15092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _10794_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _15324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _06283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _23815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _24593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _24744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _24800_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _12105_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _10806_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _12092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _12090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _12088_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _12086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _12094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _12078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _12076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _10818_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _11609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _11607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _11552_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _11591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _11872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _11554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _11605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _10816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10202_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10394_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10377_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _10174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _07651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _09915_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _09789_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _09974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _09958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _09819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _09841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _09862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _07647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _07889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _03412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _04685_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _11459_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _10366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _04679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _06454_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _10839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _10635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _07761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _04690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _06986_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _23069_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _00001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _07159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _07273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _07250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _05533_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _11840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _11183_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _05792_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _05762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _05715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _04716_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _06170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _06770_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _06441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _23931_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _02645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _02389_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _04726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _04706_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _04357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _04241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _04028_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _11736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _04785_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _09477_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _09373_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _04729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _00565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _22846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _26609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _26173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _03200_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01000_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _07439_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _07420_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _07417_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _07414_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _07412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _04031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _07063_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _07385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _07380_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _07378_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _04088_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _01214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _23609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _07308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _07348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _07345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _04101_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _07275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _07271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _07269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _07261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _07220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _07217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _07214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _07211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _07209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _07204_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _04131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _07150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _07143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _04139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _07180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _07165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _07178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _07173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _23066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _23081_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _23078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _23075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _22788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _22929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _22763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _22764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _22765_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _22830_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _01523_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _26220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _26218_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _01598_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _26237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _26235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _22909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _01596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _22833_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _22847_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _22985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _01521_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _22695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _22696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _23022_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _22694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _23052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _23001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _23031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _01547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _26184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _26162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _26181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _01603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _22893_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _22916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _22919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _26206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _22758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _22743_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _22744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _22751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _22757_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _22750_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _22756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _22741_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _26203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _22748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _22755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _22739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _22740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _22762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _22747_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _22754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _22752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _22759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _22745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _22753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _22760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _22746_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _22692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01519_);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
