
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire [15:0] _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire [7:0] _28169_;
  wire [7:0] _28170_;
  wire [7:0] _28171_;
  wire [7:0] _28172_;
  wire [7:0] _28173_;
  wire [7:0] _28174_;
  wire [7:0] _28175_;
  wire [7:0] _28176_;
  wire [7:0] _28177_;
  wire [7:0] _28178_;
  wire [7:0] _28179_;
  wire [7:0] _28180_;
  wire _28181_;
  wire [7:0] _28182_;
  wire [2:0] _28183_;
  wire [2:0] _28184_;
  wire [1:0] _28185_;
  wire [7:0] _28186_;
  wire _28187_;
  wire [1:0] _28188_;
  wire [1:0] _28189_;
  wire [2:0] _28190_;
  wire [2:0] _28191_;
  wire [1:0] _28192_;
  wire [3:0] _28193_;
  wire [1:0] _28194_;
  wire _28195_;
  wire [7:0] _28196_;
  wire [7:0] _28197_;
  wire [7:0] _28198_;
  wire [7:0] _28199_;
  wire [7:0] _28200_;
  wire [7:0] _28201_;
  wire [7:0] _28202_;
  wire [7:0] _28203_;
  wire [15:0] _28204_;
  wire [15:0] _28205_;
  wire _28206_;
  wire [4:0] _28207_;
  wire [7:0] _28208_;
  wire _28209_;
  wire _28210_;
  wire [15:0] _28211_;
  wire [15:0] _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire [7:0] _28216_;
  wire [2:0] _28217_;
  wire [7:0] _28218_;
  wire [7:0] _28219_;
  wire _28220_;
  wire [7:0] _28221_;
  wire _28222_;
  wire _28223_;
  wire [3:0] _28224_;
  wire [31:0] _28225_;
  wire [31:0] _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire [15:0] _28230_;
  wire _28231_;
  wire _28232_;
  wire [7:0] _28233_;
  wire _28234_;
  wire [2:0] _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire [3:0] _28378_;
  wire _28379_;
  wire _28380_;
  wire [7:0] _28381_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _28382_ (_23870_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _28383_ (_23871_, \oc8051_top_1.oc8051_decoder1.wr , _23870_);
  not _28384_ (_23872_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nor _28385_ (_23873_, _23872_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _28386_ (_23874_, _23873_);
  nor _28387_ (_23875_, _23874_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not _28388_ (_23876_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _28389_ (_23877_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _28390_ (_23878_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  not _28391_ (_23879_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  not _28392_ (_23880_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _28393_ (_23881_, _23880_, _23879_);
  not _28394_ (_23882_, _23881_);
  nor _28395_ (_23883_, _23882_, _23878_);
  nand _28396_ (_23884_, _23883_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _28397_ (_23885_, _23884_, _23877_);
  nand _28398_ (_23886_, _23885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _28399_ (_23887_, _23886_, _23876_);
  nor _28400_ (_23888_, _23887_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  not _28401_ (_23889_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not _28402_ (_23890_, _23875_);
  nor _28403_ (_23891_, _23890_, _23889_);
  nand _28404_ (_23892_, _23887_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand _28405_ (_23893_, _23892_, _23891_);
  nor _28406_ (_23894_, _23893_, _23888_);
  nor _28407_ (_23895_, _23874_, _23889_);
  nand _28408_ (_23896_, _23895_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not _28409_ (_23897_, _23896_);
  not _28410_ (_23898_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _28411_ (_23899_, _23889_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _28412_ (_23900_, _23899_, _23872_);
  nor _28413_ (_23901_, _23900_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not _28414_ (_23902_, _23901_);
  nor _28415_ (_23903_, _23902_, _23898_);
  nor _28416_ (_23904_, _23903_, _23897_);
  nor _28417_ (_23905_, _23890_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  nand _28418_ (_23906_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not _28419_ (_23907_, _23906_);
  not _28420_ (_23908_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  not _28421_ (_23909_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor _28422_ (_23910_, _23900_, _23909_);
  not _28423_ (_23911_, _23910_);
  nor _28424_ (_23912_, _23911_, _23908_);
  nor _28425_ (_23913_, _23912_, _23907_);
  nand _28426_ (_23914_, _23913_, _23904_);
  nor _28427_ (_23915_, _23914_, _23894_);
  nor _28428_ (_23916_, _23915_, _23875_);
  nor _28429_ (_23917_, _23916_, _23871_);
  not _28430_ (_23918_, _23917_);
  nor _28431_ (_23919_, _23883_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nand _28432_ (_23920_, _23884_, _23891_);
  nor _28433_ (_23921_, _23920_, _23919_);
  not _28434_ (_23922_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _28435_ (_23923_, _23902_, _23922_);
  nand _28436_ (_23924_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _23870_);
  nor _28437_ (_23925_, _23899_, _23873_);
  nand _28438_ (_23926_, _23925_, _23924_);
  not _28439_ (_23927_, _23926_);
  nand _28440_ (_23928_, _23927_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  not _28441_ (_23929_, _23928_);
  nor _28442_ (_23931_, _23929_, _23923_);
  not _28443_ (_23932_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nor _28444_ (_23933_, _23911_, _23932_);
  nand _28445_ (_23934_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  not _28446_ (_23935_, _23934_);
  nor _28447_ (_23936_, _23935_, _23933_);
  nand _28448_ (_23937_, _23936_, _23931_);
  nor _28449_ (_23938_, _23937_, _23921_);
  not _28450_ (_23939_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not _28451_ (_23940_, _23915_);
  nor _28452_ (_23941_, _23940_, _23939_);
  not _28453_ (_23942_, _23941_);
  nor _28454_ (_23943_, _23942_, _23938_);
  nand _28455_ (_23944_, _23910_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not _28456_ (_23945_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _28457_ (_23946_, _23902_, _23945_);
  not _28458_ (_23948_, _23946_);
  nand _28459_ (_23950_, _23948_, _23944_);
  nand _28460_ (_23951_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not _28461_ (_23952_, _23891_);
  nor _28462_ (_23953_, _23952_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  not _28463_ (_23954_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _28464_ (_23955_, _23926_, _23954_);
  nor _28465_ (_23956_, _23955_, _23953_);
  nand _28466_ (_23957_, _23956_, _23951_);
  nor _28467_ (_23958_, _23957_, _23950_);
  nor _28468_ (_23959_, _23958_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28469_ (_23960_, _23959_, _23943_);
  nor _28470_ (_23961_, _23960_, _23918_);
  not _28471_ (_23962_, _23961_);
  nand _28472_ (_23963_, _23884_, _23877_);
  nand _28473_ (_23964_, _23963_, _23891_);
  nor _28474_ (_23965_, _23964_, _23885_);
  not _28475_ (_23966_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor _28476_ (_23967_, _23911_, _23966_);
  nor _28477_ (_23968_, _23967_, _23965_);
  nand _28478_ (_23969_, _23927_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  not _28479_ (_23970_, _23969_);
  not _28480_ (_23971_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _28481_ (_23972_, _23902_, _23971_);
  nor _28482_ (_23973_, _23972_, _23970_);
  not _28483_ (_23974_, _23973_);
  nand _28484_ (_23975_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nand _28485_ (_23976_, _23975_, _23896_);
  nor _28486_ (_23977_, _23976_, _23974_);
  nand _28487_ (_23978_, _23977_, _23968_);
  not _28488_ (_23979_, _23978_);
  nor _28489_ (_23980_, _23979_, _23942_);
  nor _28490_ (_23981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _28491_ (_23982_, _23981_, _23881_);
  nand _28492_ (_23984_, _23982_, _23891_);
  nand _28493_ (_23985_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nand _28494_ (_23986_, _23985_, _23984_);
  not _28495_ (_23987_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor _28496_ (_23988_, _23902_, _23987_);
  not _28497_ (_23989_, _23988_);
  not _28498_ (_23990_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nor _28499_ (_23991_, _23911_, _23990_);
  nand _28500_ (_23992_, _23927_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  not _28501_ (_23993_, _23992_);
  nor _28502_ (_23994_, _23993_, _23991_);
  nand _28503_ (_23995_, _23994_, _23989_);
  nor _28504_ (_23996_, _23995_, _23986_);
  nor _28505_ (_23997_, _23996_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28506_ (_23998_, _23997_, _23980_);
  nor _28507_ (_23999_, _23998_, _23918_);
  nor _28508_ (_24000_, _23999_, _23962_);
  not _28509_ (_24001_, _24000_);
  nand _28510_ (_24002_, _23886_, _23876_);
  nand _28511_ (_24003_, _24002_, _23891_);
  nor _28512_ (_24004_, _24003_, _23887_);
  not _28513_ (_24005_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _28514_ (_24006_, _23902_, _24005_);
  nor _28515_ (_24007_, _24006_, _23897_);
  nand _28516_ (_24009_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  not _28517_ (_24010_, _24009_);
  not _28518_ (_24012_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor _28519_ (_24013_, _23911_, _24012_);
  nor _28520_ (_24014_, _24013_, _24010_);
  nand _28521_ (_24015_, _24014_, _24007_);
  nor _28522_ (_24016_, _24015_, _24004_);
  nor _28523_ (_24017_, _24016_, _23942_);
  nor _28524_ (_24018_, _23941_, _23938_);
  nor _28525_ (_24019_, _24018_, _24017_);
  nor _28526_ (_24020_, _24019_, _23918_);
  not _28527_ (_24021_, _24020_);
  nor _28528_ (_24023_, _23885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand _28529_ (_24024_, _23886_, _23891_);
  nor _28530_ (_24025_, _24024_, _24023_);
  not _28531_ (_24026_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _28532_ (_24027_, _23902_, _24026_);
  nor _28533_ (_24028_, _24027_, _23897_);
  nand _28534_ (_24029_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  not _28535_ (_24030_, _24029_);
  not _28536_ (_24031_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor _28537_ (_24032_, _23911_, _24031_);
  nor _28538_ (_24033_, _24032_, _24030_);
  nand _28539_ (_24034_, _24033_, _24028_);
  nor _28540_ (_24035_, _24034_, _24025_);
  nor _28541_ (_24036_, _24035_, _23942_);
  nor _28542_ (_24037_, _23881_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _28543_ (_24038_, _24037_, _23883_);
  nand _28544_ (_24039_, _24038_, _23891_);
  nand _28545_ (_24040_, _23905_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nand _28546_ (_24041_, _24040_, _24039_);
  not _28547_ (_24042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor _28548_ (_24043_, _23902_, _24042_);
  not _28549_ (_24044_, _24043_);
  not _28550_ (_24045_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  nor _28551_ (_24046_, _23911_, _24045_);
  nand _28552_ (_24047_, _23927_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  not _28553_ (_24048_, _24047_);
  nor _28554_ (_24049_, _24048_, _24046_);
  nand _28555_ (_24050_, _24049_, _24044_);
  nor _28556_ (_24051_, _24050_, _24041_);
  nor _28557_ (_24052_, _24051_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28558_ (_24053_, _24052_, _24036_);
  nor _28559_ (_24054_, _24053_, _23918_);
  not _28560_ (_24055_, _24054_);
  nor _28561_ (_24056_, _24055_, _24021_);
  not _28562_ (_24057_, _24056_);
  nor _28563_ (_24058_, _24057_, _24001_);
  not _28564_ (_24059_, _24058_);
  not _28565_ (_24060_, _24035_);
  nor _28566_ (_24061_, _24060_, _23941_);
  nor _28567_ (_24062_, _24061_, _23918_);
  not _28568_ (_24063_, _24062_);
  nor _28569_ (_24064_, _23979_, _23941_);
  not _28570_ (_24065_, _24064_);
  nor _28571_ (_24066_, _24065_, _23918_);
  nor _28572_ (_24067_, _24066_, _24063_);
  not _28573_ (_24068_, _24067_);
  not _28574_ (_24069_, _24016_);
  nor _28575_ (_24070_, _24069_, _23915_);
  not _28576_ (_24071_, _24070_);
  nor _28577_ (_24072_, _24071_, _24068_);
  not _28578_ (_24073_, _24072_);
  nor _28579_ (_24074_, _24073_, _24059_);
  not _28580_ (_24075_, _24074_);
  nand _28581_ (_24076_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  not _28582_ (_24077_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  nor _28583_ (_24078_, \oc8051_top_1.oc8051_sfr1.wait_data , _24077_);
  not _28584_ (_24079_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  nor _28585_ (_24080_, _24079_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _28586_ (_24081_, _24080_, _24078_);
  not _28587_ (_24082_, _24081_);
  not _28588_ (_24083_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  nor _28589_ (_24084_, _24083_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _28590_ (_24085_, _24084_);
  nor _28591_ (_24086_, _24085_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not _28592_ (_24087_, _24086_);
  nor _28593_ (_24088_, _24087_, _24082_);
  not _28594_ (_24089_, _24088_);
  not _28595_ (_24090_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _28596_ (_24091_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nor _28597_ (_24092_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _24091_);
  nand _28598_ (_24093_, _24092_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor _28599_ (_24094_, _24093_, _24090_);
  not _28600_ (_24095_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _28601_ (_24096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _28602_ (_24097_, _24096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor _28603_ (_24098_, _24097_, _24095_);
  nor _28604_ (_24099_, _24098_, _24094_);
  not _28605_ (_24100_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _28606_ (_24102_, _24092_, _24100_);
  nor _28607_ (_24103_, _24102_, _23898_);
  nor _28608_ (_24104_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _28609_ (_24105_, _24104_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nor _28610_ (_24106_, _24105_, _23908_);
  nor _28611_ (_24108_, _24106_, _24103_);
  nand _28612_ (_24109_, _24108_, _24099_);
  not _28613_ (_24110_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _28614_ (_24111_, _24104_, _24110_);
  not _28615_ (_24112_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  nand _28616_ (_24113_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _24112_);
  nor _28617_ (_24114_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not _28618_ (_24115_, _24114_);
  not _28619_ (_24116_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nand _28620_ (_24117_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , _24116_);
  nand _28621_ (_24118_, _24117_, _24115_);
  nand _28622_ (_24119_, _24118_, _24113_);
  nor _28623_ (_24120_, _24113_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  not _28624_ (_24121_, _24120_);
  nand _28625_ (_24122_, _24121_, _24119_);
  nor _28626_ (_24123_, _24122_, _24111_);
  not _28627_ (_24124_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _28628_ (_24125_, _24110_, _24091_);
  nand _28629_ (_24126_, _24125_, _24100_);
  nor _28630_ (_24127_, _24126_, _24124_);
  nand _28631_ (_24128_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nor _28632_ (_24129_, _24128_, _24100_);
  nand _28633_ (_24130_, _24129_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  not _28634_ (_24131_, _24130_);
  nor _28635_ (_24132_, _24131_, _24127_);
  not _28636_ (_24133_, _24132_);
  nor _28637_ (_24135_, _24133_, _24123_);
  not _28638_ (_24136_, _24135_);
  nor _28639_ (_24137_, _24136_, _24109_);
  nor _28640_ (_24138_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not _28641_ (_24139_, _24138_);
  nor _28642_ (_24140_, _24139_, _24122_);
  nand _28643_ (_24142_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor _28644_ (_24143_, _24142_, _23898_);
  not _28645_ (_24144_, _24143_);
  not _28646_ (_24145_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor _28647_ (_24146_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], _24145_);
  nand _28648_ (_24147_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand _28649_ (_24148_, _24147_, _24144_);
  nor _28650_ (_24149_, _24148_, _24140_);
  nor _28651_ (_24150_, _24149_, _24137_);
  not _28652_ (_24151_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _28653_ (_24152_, _24097_, _24151_);
  not _28654_ (_24153_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _28655_ (_24154_, _24093_, _24153_);
  nor _28656_ (_24155_, _24154_, _24152_);
  nor _28657_ (_24156_, _24128_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _28658_ (_24157_, _24156_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not _28659_ (_24158_, _24157_);
  nor _28660_ (_24159_, _24105_, _24031_);
  nor _28661_ (_24160_, _24159_, _24158_);
  nand _28662_ (_24161_, _24160_, _24155_);
  not _28663_ (_24162_, _24111_);
  not _28664_ (_24163_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor _28665_ (_24164_, _24163_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  nor _28666_ (_24165_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  not _28667_ (_24166_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor _28668_ (_24167_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _24166_);
  nor _28669_ (_24169_, _24167_, _24165_);
  nor _28670_ (_24170_, _24169_, _24164_);
  nor _28671_ (_24171_, _24113_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor _28672_ (_24172_, _24171_, _24170_);
  nand _28673_ (_24173_, _24172_, _24162_);
  nor _28674_ (_24174_, _24102_, _24026_);
  nand _28675_ (_24175_, _24129_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  not _28676_ (_24176_, _24175_);
  nor _28677_ (_24177_, _24176_, _24174_);
  nand _28678_ (_24178_, _24177_, _24173_);
  nor _28679_ (_24179_, _24178_, _24161_);
  not _28680_ (_24180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nand _28681_ (_24181_, _24166_, _24180_);
  not _28682_ (_24182_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5]);
  nand _28683_ (_24183_, _24182_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nand _28684_ (_24184_, _24183_, _24181_);
  nand _28685_ (_24185_, _24184_, _24113_);
  not _28686_ (_24186_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _28687_ (_24187_, _24164_, _24186_);
  nand _28688_ (_24188_, _24187_, _24185_);
  nor _28689_ (_24189_, _24188_, _24139_);
  nor _28690_ (_24190_, _24142_, _24026_);
  not _28691_ (_24191_, _24190_);
  nand _28692_ (_24192_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _28693_ (_24193_, _24192_, _24191_);
  nor _28694_ (_24194_, _24193_, _24189_);
  nor _28695_ (_24195_, _24194_, _24179_);
  not _28696_ (_24196_, _24179_);
  nand _28697_ (_24197_, _24172_, _24138_);
  not _28698_ (_24198_, _24193_);
  nand _28699_ (_24199_, _24198_, _24197_);
  nor _28700_ (_24200_, _24199_, _24196_);
  nor _28701_ (_24201_, _24200_, _24195_);
  not _28702_ (_24202_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _28703_ (_24203_, _24093_, _24202_);
  not _28704_ (_24204_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _28705_ (_24205_, _24097_, _24204_);
  nor _28706_ (_24206_, _24205_, _24203_);
  nor _28707_ (_24207_, _24102_, _23971_);
  nor _28708_ (_24208_, _24105_, _23966_);
  nor _28709_ (_24209_, _24208_, _24207_);
  nand _28710_ (_24210_, _24209_, _24206_);
  nor _28711_ (_24211_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor _28712_ (_24212_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _24166_);
  nor _28713_ (_24213_, _24212_, _24211_);
  nor _28714_ (_24214_, _24213_, _24164_);
  nor _28715_ (_24215_, _24113_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor _28716_ (_24216_, _24215_, _24214_);
  nand _28717_ (_24217_, _24216_, _24162_);
  nand _28718_ (_24218_, _24156_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _28719_ (_24220_, _24129_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nand _28720_ (_24221_, _24220_, _24218_);
  not _28721_ (_24222_, _24221_);
  nand _28722_ (_24223_, _24222_, _24217_);
  nor _28723_ (_24224_, _24223_, _24210_);
  not _28724_ (_24225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nand _28725_ (_24226_, _24166_, _24225_);
  not _28726_ (_24227_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4]);
  nand _28727_ (_24228_, _24227_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nand _28728_ (_24229_, _24228_, _24226_);
  nand _28729_ (_24230_, _24229_, _24113_);
  not _28730_ (_24231_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _28731_ (_24232_, _24164_, _24231_);
  nand _28732_ (_24234_, _24232_, _24230_);
  nor _28733_ (_24235_, _24234_, _24139_);
  nor _28734_ (_24236_, _24142_, _23971_);
  not _28735_ (_24237_, _24236_);
  nand _28736_ (_24239_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _28737_ (_24240_, _24239_, _24237_);
  nor _28738_ (_24241_, _24240_, _24235_);
  nor _28739_ (_24242_, _24241_, _24224_);
  not _28740_ (_24243_, _24224_);
  nand _28741_ (_24244_, _24216_, _24138_);
  not _28742_ (_24245_, _24240_);
  nand _28743_ (_24247_, _24245_, _24244_);
  nor _28744_ (_24248_, _24247_, _24243_);
  nor _28745_ (_24249_, _24248_, _24242_);
  not _28746_ (_24250_, _24249_);
  not _28747_ (_24251_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _28748_ (_24252_, _24093_, _24251_);
  not _28749_ (_24253_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _28750_ (_24254_, _24097_, _24253_);
  nor _28751_ (_24255_, _24254_, _24252_);
  nor _28752_ (_24256_, _24102_, _23922_);
  nor _28753_ (_24257_, _24105_, _23932_);
  nor _28754_ (_24258_, _24257_, _24256_);
  nand _28755_ (_24259_, _24258_, _24255_);
  not _28756_ (_24260_, _24259_);
  not _28757_ (_24261_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nor _28758_ (_24262_, _24113_, _24261_);
  not _28759_ (_24263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nand _28760_ (_24264_, _24166_, _24263_);
  not _28761_ (_24265_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3]);
  nand _28762_ (_24266_, _24265_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nand _28763_ (_24267_, _24266_, _24264_);
  nor _28764_ (_24268_, _24267_, _24164_);
  nor _28765_ (_24269_, _24268_, _24262_);
  nor _28766_ (_24270_, _24269_, _24111_);
  not _28767_ (_24271_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _28768_ (_24272_, _24126_, _24271_);
  nand _28769_ (_24273_, _24129_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not _28770_ (_24274_, _24273_);
  nor _28771_ (_24275_, _24274_, _24272_);
  not _28772_ (_24276_, _24275_);
  nor _28773_ (_24277_, _24276_, _24270_);
  nand _28774_ (_24278_, _24277_, _24260_);
  not _28775_ (_24279_, _24278_);
  nor _28776_ (_24280_, _24269_, _24139_);
  nor _28777_ (_24281_, _24142_, _23922_);
  not _28778_ (_24282_, _24281_);
  nand _28779_ (_24283_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand _28780_ (_24284_, _24283_, _24282_);
  nor _28781_ (_24285_, _24284_, _24280_);
  nor _28782_ (_24286_, _24285_, _24279_);
  nand _28783_ (_24287_, _24164_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nor _28784_ (_24288_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor _28785_ (_24289_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _24166_);
  nor _28786_ (_24290_, _24289_, _24288_);
  nand _28787_ (_24292_, _24290_, _24113_);
  nand _28788_ (_24293_, _24292_, _24287_);
  nand _28789_ (_24294_, _24293_, _24138_);
  not _28790_ (_24295_, _24284_);
  nand _28791_ (_24296_, _24295_, _24294_);
  nor _28792_ (_24297_, _24296_, _24278_);
  nor _28793_ (_24298_, _24297_, _24286_);
  not _28794_ (_24299_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand _28795_ (_24300_, _24125_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor _28796_ (_24301_, _24300_, _24299_);
  not _28797_ (_24302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _28798_ (_24303_, _24126_, _24302_);
  nor _28799_ (_24304_, _24303_, _24301_);
  not _28800_ (_24305_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _28801_ (_24306_, _24093_, _24305_);
  not _28802_ (_24308_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _28803_ (_24309_, _24097_, _24308_);
  nor _28804_ (_24310_, _24309_, _24306_);
  nand _28805_ (_24311_, _24310_, _24304_);
  nor _28806_ (_24312_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  nor _28807_ (_24313_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _24166_);
  nor _28808_ (_24314_, _24313_, _24312_);
  nor _28809_ (_24315_, _24314_, _24164_);
  nor _28810_ (_24316_, _24113_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nor _28811_ (_24317_, _24316_, _24315_);
  nand _28812_ (_24318_, _24317_, _24162_);
  nor _28813_ (_24319_, _24102_, _24042_);
  nor _28814_ (_24320_, _24105_, _24045_);
  nor _28815_ (_24321_, _24320_, _24319_);
  nand _28816_ (_24322_, _24321_, _24318_);
  nor _28817_ (_24323_, _24322_, _24311_);
  not _28818_ (_24324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  nand _28819_ (_24325_, _24166_, _24324_);
  not _28820_ (_24326_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2]);
  nand _28821_ (_24327_, _24326_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nand _28822_ (_24328_, _24327_, _24325_);
  nand _28823_ (_24329_, _24328_, _24113_);
  not _28824_ (_24330_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _28825_ (_24331_, _24164_, _24330_);
  nand _28826_ (_24332_, _24331_, _24329_);
  nor _28827_ (_24333_, _24332_, _24139_);
  nor _28828_ (_24334_, _24142_, _24042_);
  not _28829_ (_24335_, _24334_);
  nand _28830_ (_24336_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand _28831_ (_24337_, _24336_, _24335_);
  nor _28832_ (_24338_, _24337_, _24333_);
  nor _28833_ (_24339_, _24338_, _24323_);
  nand _28834_ (_24340_, _24110_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nor _28835_ (_24342_, _24340_, _24100_);
  nand _28836_ (_24343_, _24342_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _28837_ (_24344_, _24340_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _28838_ (_24345_, _24344_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand _28839_ (_24346_, _24345_, _24343_);
  nor _28840_ (_24347_, _24320_, _24309_);
  nand _28841_ (_24348_, _24347_, _24304_);
  nor _28842_ (_24349_, _24348_, _24346_);
  nand _28843_ (_24350_, _24349_, _24318_);
  nand _28844_ (_24351_, _24317_, _24138_);
  not _28845_ (_24352_, _24337_);
  nand _28846_ (_24353_, _24352_, _24351_);
  nor _28847_ (_24354_, _24353_, _24350_);
  nor _28848_ (_24355_, _24354_, _24339_);
  not _28849_ (_24356_, _24355_);
  nor _28850_ (_24357_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor _28851_ (_24358_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _24166_);
  nor _28852_ (_24359_, _24358_, _24357_);
  nor _28853_ (_24360_, _24359_, _24164_);
  nor _28854_ (_24361_, _24113_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nor _28855_ (_24362_, _24361_, _24360_);
  nand _28856_ (_24363_, _24362_, _24162_);
  not _28857_ (_24364_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _28858_ (_24365_, _24093_, _24364_);
  not _28859_ (_24366_, _24365_);
  nor _28860_ (_24367_, _24102_, _23987_);
  not _28861_ (_24368_, _24367_);
  nand _28862_ (_24369_, _24368_, _24366_);
  nand _28863_ (_24370_, _24156_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand _28864_ (_24371_, _24129_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand _28865_ (_24372_, _24371_, _24370_);
  not _28866_ (_24373_, _24372_);
  not _28867_ (_24374_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _28868_ (_24375_, _24097_, _24374_);
  nor _28869_ (_24376_, _24105_, _23990_);
  nor _28870_ (_24377_, _24376_, _24375_);
  nand _28871_ (_24378_, _24377_, _24373_);
  nor _28872_ (_24379_, _24378_, _24369_);
  nand _28873_ (_24380_, _24379_, _24363_);
  not _28874_ (_24381_, _24380_);
  not _28875_ (_24382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nand _28876_ (_24383_, _24166_, _24382_);
  not _28877_ (_24384_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1]);
  nand _28878_ (_24385_, _24384_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nand _28879_ (_24386_, _24385_, _24383_);
  nand _28880_ (_24387_, _24386_, _24113_);
  not _28881_ (_24388_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _28882_ (_24389_, _24164_, _24388_);
  nand _28883_ (_24390_, _24389_, _24387_);
  nor _28884_ (_24391_, _24390_, _24139_);
  nor _28885_ (_24392_, _24142_, _23987_);
  not _28886_ (_24393_, _24392_);
  nand _28887_ (_24394_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand _28888_ (_24395_, _24394_, _24393_);
  nor _28889_ (_24396_, _24395_, _24391_);
  nor _28890_ (_24397_, _24396_, _24381_);
  not _28891_ (_24398_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _28892_ (_24400_, _24097_, _24398_);
  not _28893_ (_24401_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _28894_ (_24402_, _24093_, _24401_);
  nor _28895_ (_24403_, _24402_, _24400_);
  not _28896_ (_24404_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _28897_ (_24405_, _24126_, _24404_);
  not _28898_ (_24406_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor _28899_ (_24407_, _24105_, _24406_);
  nor _28900_ (_24408_, _24407_, _24405_);
  nand _28901_ (_24409_, _24408_, _24403_);
  not _28902_ (_24410_, _24409_);
  not _28903_ (_24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nand _28904_ (_24412_, _24166_, _24411_);
  not _28905_ (_24413_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0]);
  nand _28906_ (_24414_, _24413_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nand _28907_ (_24415_, _24414_, _24412_);
  nand _28908_ (_24416_, _24415_, _24113_);
  not _28909_ (_24417_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _28910_ (_24418_, _24164_, _24417_);
  nand _28911_ (_24419_, _24418_, _24416_);
  nor _28912_ (_24420_, _24419_, _24111_);
  nor _28913_ (_24421_, _24102_, _23945_);
  nand _28914_ (_24422_, _24129_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not _28915_ (_24423_, _24422_);
  nor _28916_ (_24424_, _24423_, _24421_);
  not _28917_ (_24425_, _24424_);
  nor _28918_ (_24426_, _24425_, _24420_);
  nand _28919_ (_24427_, _24426_, _24410_);
  not _28920_ (_24428_, _24427_);
  nor _28921_ (_24429_, _24419_, _24139_);
  nor _28922_ (_24430_, _24142_, _23945_);
  not _28923_ (_24431_, _24430_);
  nand _28924_ (_24432_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nand _28925_ (_24433_, _24432_, _24431_);
  nor _28926_ (_24434_, _24433_, _24429_);
  nor _28927_ (_24435_, _24434_, _24428_);
  not _28928_ (_24436_, _24435_);
  nand _28929_ (_24437_, _24362_, _24138_);
  not _28930_ (_24438_, _24395_);
  nand _28931_ (_24439_, _24438_, _24437_);
  nor _28932_ (_24440_, _24439_, _24380_);
  nor _28933_ (_24441_, _24440_, _24397_);
  not _28934_ (_24442_, _24441_);
  nor _28935_ (_24443_, _24442_, _24436_);
  nor _28936_ (_24444_, _24443_, _24397_);
  nor _28937_ (_24445_, _24444_, _24356_);
  nor _28938_ (_24446_, _24445_, _24339_);
  nor _28939_ (_24447_, _24446_, _24298_);
  nand _28940_ (_24448_, _24446_, _24298_);
  not _28941_ (_24449_, _24448_);
  nor _28942_ (_24450_, _24449_, _24447_);
  nor _28943_ (_24451_, _24113_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not _28944_ (_24452_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not _28945_ (_24453_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor _28946_ (_24454_, _24453_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  not _28947_ (_24455_, _24454_);
  nor _28948_ (_24456_, _24455_, _24184_);
  nor _28949_ (_24457_, _24456_, _24452_);
  not _28950_ (_24458_, _24457_);
  nor _28951_ (_24459_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  not _28952_ (_24460_, _24459_);
  nor _28953_ (_24461_, _24460_, _24229_);
  not _28954_ (_24462_, _24461_);
  nand _28955_ (_24463_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nor _28956_ (_24464_, _24463_, _24118_);
  nor _28957_ (_24465_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  not _28958_ (_24466_, _24465_);
  not _28959_ (_24467_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6]);
  nand _28960_ (_24468_, _24467_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nand _28961_ (_24469_, _24468_, _24466_);
  nand _28962_ (_24470_, _24453_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nor _28963_ (_24471_, _24470_, _24469_);
  nor _28964_ (_24472_, _24471_, _24464_);
  nand _28965_ (_24473_, _24472_, _24462_);
  nor _28966_ (_24474_, _24473_, _24458_);
  nor _28967_ (_24475_, _24455_, _24386_);
  nor _28968_ (_24476_, _24475_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not _28969_ (_24477_, _24476_);
  nor _28970_ (_24478_, _24470_, _24328_);
  not _28971_ (_24479_, _24478_);
  nor _28972_ (_24480_, _24463_, _24267_);
  nor _28973_ (_24481_, _24460_, _24415_);
  nor _28974_ (_24482_, _24481_, _24480_);
  nand _28975_ (_24483_, _24482_, _24479_);
  nor _28976_ (_24484_, _24483_, _24477_);
  nor _28977_ (_24485_, _24484_, _24474_);
  nor _28978_ (_24486_, _24485_, _24164_);
  nor _28979_ (_24488_, _24486_, _24451_);
  not _28980_ (_24489_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not _28981_ (_24490_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _28982_ (_24491_, _24490_, _24489_);
  nor _28983_ (_24492_, _24491_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _28984_ (_24493_, _24492_);
  nand _28985_ (_24494_, _24493_, _24488_);
  nor _28986_ (_24495_, _24492_, _24489_);
  not _28987_ (_24496_, _24495_);
  nand _28988_ (_24497_, _24496_, _24494_);
  not _28989_ (_24498_, _24497_);
  nor _28990_ (_24499_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor _28991_ (_24500_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _24166_);
  nor _28992_ (_24501_, _24500_, _24499_);
  nor _28993_ (_24502_, _24501_, _24164_);
  nor _28994_ (_24504_, _24113_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nor _28995_ (_24505_, _24504_, _24502_);
  nand _28996_ (_24506_, _24505_, _24138_);
  not _28997_ (_24507_, _24433_);
  nand _28998_ (_24508_, _24507_, _24506_);
  nor _28999_ (_24509_, _24508_, _24427_);
  nor _29000_ (_24510_, _24509_, _24435_);
  not _29001_ (_24511_, _24510_);
  nor _29002_ (_24512_, _24511_, _24498_);
  not _29003_ (_24513_, _24512_);
  nor _29004_ (_24514_, _24513_, _24442_);
  nand _29005_ (_24515_, _24444_, _24356_);
  not _29006_ (_24516_, _24515_);
  nor _29007_ (_24517_, _24516_, _24445_);
  nand _29008_ (_24518_, _24517_, _24514_);
  nor _29009_ (_24519_, _24518_, _24450_);
  nor _29010_ (_24520_, _24446_, _24297_);
  nor _29011_ (_24521_, _24520_, _24286_);
  not _29012_ (_24522_, _24521_);
  nor _29013_ (_24523_, _24522_, _24519_);
  nor _29014_ (_24524_, _24523_, _24250_);
  nand _29015_ (_24525_, _24524_, _24201_);
  not _29016_ (_24527_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _29017_ (_24528_, _24093_, _24527_);
  not _29018_ (_24529_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _29019_ (_24530_, _24097_, _24529_);
  nor _29020_ (_24531_, _24530_, _24528_);
  nor _29021_ (_24532_, _24102_, _24005_);
  nor _29022_ (_24533_, _24105_, _24012_);
  nor _29023_ (_24534_, _24533_, _24532_);
  nand _29024_ (_24535_, _24534_, _24531_);
  nand _29025_ (_24536_, _24469_, _24113_);
  nor _29026_ (_24537_, _24113_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  not _29027_ (_24538_, _24537_);
  nand _29028_ (_24539_, _24538_, _24536_);
  nor _29029_ (_24540_, _24539_, _24111_);
  not _29030_ (_24541_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _29031_ (_24542_, _24126_, _24541_);
  nand _29032_ (_24543_, _24129_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  not _29033_ (_24544_, _24543_);
  nor _29034_ (_24545_, _24544_, _24542_);
  not _29035_ (_24546_, _24545_);
  nor _29036_ (_24547_, _24546_, _24540_);
  not _29037_ (_24548_, _24547_);
  nor _29038_ (_24549_, _24548_, _24535_);
  nor _29039_ (_24550_, _24539_, _24139_);
  nor _29040_ (_24551_, _24142_, _24005_);
  not _29041_ (_24552_, _24551_);
  nand _29042_ (_24553_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _29043_ (_24554_, _24553_, _24552_);
  nor _29044_ (_24555_, _24554_, _24550_);
  nor _29045_ (_24556_, _24555_, _24549_);
  not _29046_ (_24557_, _24549_);
  not _29047_ (_24558_, _24555_);
  nor _29048_ (_24559_, _24558_, _24557_);
  nor _29049_ (_24560_, _24559_, _24556_);
  not _29050_ (_24561_, _24560_);
  not _29051_ (_24562_, _24201_);
  not _29052_ (_24563_, _24242_);
  nor _29053_ (_24564_, _24563_, _24562_);
  nor _29054_ (_24565_, _24564_, _24195_);
  nor _29055_ (_24566_, _24565_, _24561_);
  not _29056_ (_24567_, _24566_);
  nand _29057_ (_24568_, _24565_, _24561_);
  nand _29058_ (_24569_, _24568_, _24567_);
  nor _29059_ (_24570_, _24569_, _24525_);
  nor _29060_ (_24571_, _24566_, _24556_);
  not _29061_ (_24573_, _24571_);
  nor _29062_ (_24574_, _24573_, _24570_);
  not _29063_ (_24575_, _24137_);
  not _29064_ (_24576_, _24149_);
  nor _29065_ (_24577_, _24576_, _24575_);
  nor _29066_ (_24578_, _24577_, _24150_);
  not _29067_ (_24579_, _24578_);
  nor _29068_ (_24580_, _24579_, _24574_);
  nor _29069_ (_24581_, _24580_, _24150_);
  nor _29070_ (_24582_, _24581_, _24089_);
  not _29071_ (_24583_, _24582_);
  not _29072_ (_24584_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  nor _29073_ (_24585_, _24584_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29074_ (_24586_, _24585_);
  nor _29075_ (_24588_, _24586_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  not _29076_ (_24589_, _24588_);
  nor _29077_ (_24590_, _24589_, _24082_);
  not _29078_ (_24591_, _24590_);
  nor _29079_ (_24592_, _24149_, _24575_);
  nor _29080_ (_24593_, _24558_, _24549_);
  nor _29081_ (_24594_, _24199_, _24179_);
  nor _29082_ (_24595_, _24241_, _24243_);
  nor _29083_ (_24597_, _24595_, _24201_);
  nor _29084_ (_24599_, _24597_, _24594_);
  nor _29085_ (_24600_, _24599_, _24560_);
  nor _29086_ (_24601_, _24600_, _24593_);
  nand _29087_ (_24602_, _24599_, _24560_);
  not _29088_ (_24603_, _24602_);
  nor _29089_ (_24604_, _24603_, _24600_);
  nand _29090_ (_24605_, _24595_, _24201_);
  not _29091_ (_24606_, _24605_);
  nor _29092_ (_24607_, _24606_, _24597_);
  nor _29093_ (_24609_, _24434_, _24427_);
  nor _29094_ (_24610_, _24609_, _24441_);
  nor _29095_ (_24611_, _24439_, _24381_);
  nor _29096_ (_24612_, _24611_, _24610_);
  nor _29097_ (_24613_, _24612_, _24355_);
  nor _29098_ (_24614_, _24353_, _24323_);
  nor _29099_ (_24616_, _24614_, _24613_);
  nor _29100_ (_24617_, _24616_, _24298_);
  not _29101_ (_24618_, _24298_);
  not _29102_ (_24619_, _24616_);
  nor _29103_ (_24620_, _24619_, _24618_);
  nor _29104_ (_24621_, _24620_, _24617_);
  nand _29105_ (_24622_, _24612_, _24355_);
  not _29106_ (_24623_, _24622_);
  nor _29107_ (_24624_, _24623_, _24613_);
  nand _29108_ (_24625_, _24609_, _24441_);
  not _29109_ (_24626_, _24625_);
  nor _29110_ (_24627_, _24626_, _24610_);
  nor _29111_ (_24628_, _24510_, _24498_);
  not _29112_ (_24629_, _24628_);
  nor _29113_ (_24630_, _24629_, _24627_);
  not _29114_ (_24631_, _24630_);
  nor _29115_ (_24632_, _24631_, _24624_);
  not _29116_ (_24633_, _24632_);
  nor _29117_ (_24634_, _24633_, _24621_);
  nor _29118_ (_24635_, _24296_, _24279_);
  nor _29119_ (_24636_, _24285_, _24278_);
  nor _29120_ (_24637_, _24616_, _24636_);
  nor _29121_ (_24638_, _24637_, _24635_);
  nor _29122_ (_24639_, _24638_, _24634_);
  nor _29123_ (_24640_, _24639_, _24249_);
  not _29124_ (_24641_, _24640_);
  nor _29125_ (_24642_, _24641_, _24607_);
  not _29126_ (_24643_, _24642_);
  nor _29127_ (_24644_, _24643_, _24604_);
  nor _29128_ (_24645_, _24644_, _24601_);
  nor _29129_ (_24646_, _24645_, _24578_);
  nor _29130_ (_24647_, _24646_, _24592_);
  nor _29131_ (_24648_, _24647_, _24591_);
  nand _29132_ (_24649_, _24080_, _24077_);
  nor _29133_ (_24650_, _24649_, _24087_);
  not _29134_ (_24651_, _24650_);
  nor _29135_ (_24653_, _24557_, _24196_);
  nor _29136_ (_24654_, _24653_, _24137_);
  nor _29137_ (_24655_, _24654_, _24498_);
  nor _29138_ (_24656_, _24380_, _24350_);
  nor _29139_ (_24657_, _24656_, _24279_);
  not _29140_ (_24658_, _24654_);
  nor _29141_ (_24659_, _24658_, _24497_);
  nor _29142_ (_24661_, _24659_, _24657_);
  not _29143_ (_24663_, _24661_);
  nor _29144_ (_24664_, _24663_, _24655_);
  nor _29145_ (_24665_, _24664_, _24651_);
  nor _29146_ (_24666_, _24585_, _24084_);
  not _29147_ (_24667_, _24666_);
  nor _29148_ (_24668_, _24667_, _24082_);
  nor _29149_ (_24669_, _24668_, _24498_);
  nor _29150_ (_24670_, _24649_, _24589_);
  nor _29151_ (_24671_, _24670_, _24497_);
  nor _29152_ (_24672_, _24671_, _24669_);
  nor _29153_ (_24673_, _24495_, _24488_);
  not _29154_ (_24674_, _24078_);
  nor _29155_ (_24675_, _24674_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  not _29156_ (_24676_, _24675_);
  nor _29157_ (_24677_, _24676_, _24087_);
  not _29158_ (_24678_, _24494_);
  nor _29159_ (_24679_, _24676_, _24667_);
  not _29160_ (_24680_, _24679_);
  nor _29161_ (_24681_, _24680_, _24678_);
  nor _29162_ (_24682_, _24681_, _24677_);
  nor _29163_ (_24683_, _24682_, _24673_);
  not _29164_ (_24684_, _24488_);
  nor _29165_ (_24685_, _24493_, _24684_);
  nor _29166_ (_24686_, _24676_, _24589_);
  nor _29167_ (_24687_, _24586_, _24083_);
  not _29168_ (_24688_, _24687_);
  nor _29169_ (_24689_, _24688_, _24649_);
  not _29170_ (_24690_, _24689_);
  nor _29171_ (_24691_, _24690_, _24684_);
  nor _29172_ (_24692_, _24691_, _24686_);
  nor _29173_ (_24693_, _24692_, _24685_);
  nor _29174_ (_24694_, _24498_, _24488_);
  nor _29175_ (_24695_, _24674_, _24079_);
  not _29176_ (_24696_, _24695_);
  nor _29177_ (_24697_, _24696_, _24667_);
  nand _29178_ (_24698_, _24697_, _24694_);
  nor _29179_ (_24699_, _24676_, _24688_);
  not _29180_ (_24700_, _24699_);
  nor _29181_ (_24701_, _24700_, _24137_);
  nor _29182_ (_24702_, _24696_, _24087_);
  not _29183_ (_24703_, _24702_);
  nor _29184_ (_24704_, _24703_, _24428_);
  nor _29185_ (_24705_, _24704_, _24701_);
  nand _29186_ (_24706_, _24705_, _24698_);
  nor _29187_ (_24707_, _24706_, _24693_);
  not _29188_ (_24708_, _24707_);
  nor _29189_ (_24709_, _24708_, _24683_);
  not _29190_ (_24710_, _24709_);
  nor _29191_ (_24711_, _24710_, _24672_);
  not _29192_ (_24712_, _24711_);
  nor _29193_ (_24713_, _24712_, _24665_);
  not _29194_ (_24714_, _24713_);
  nor _29195_ (_24715_, _24714_, _24648_);
  nand _29196_ (_24716_, _24715_, _24583_);
  not _29197_ (_24717_, _24716_);
  not _29198_ (_24718_, _24463_);
  nor _29199_ (_24719_, _24452_, _23939_);
  nand _29200_ (_24721_, _24719_, _24718_);
  nor _29201_ (_24722_, _24721_, _24717_);
  nor _29202_ (_24723_, _24427_, _24380_);
  nand _29203_ (_24724_, _24723_, _24323_);
  nor _29204_ (_24725_, _24724_, _24278_);
  not _29205_ (_24726_, _24725_);
  nor _29206_ (_24727_, _24726_, _24243_);
  nand _29207_ (_24728_, _24727_, _24179_);
  nor _29208_ (_24729_, _24728_, _24557_);
  nor _29209_ (_24730_, _24729_, _24498_);
  nand _29210_ (_24731_, _24427_, _24380_);
  nor _29211_ (_24732_, _24731_, _24323_);
  nand _29212_ (_24733_, _24732_, _24278_);
  nor _29213_ (_24734_, _24733_, _24224_);
  not _29214_ (_24735_, _24734_);
  nor _29215_ (_24736_, _24735_, _24179_);
  nand _29216_ (_24737_, _24736_, _24557_);
  nand _29217_ (_24738_, _24737_, _24498_);
  not _29218_ (_24739_, _24738_);
  nor _29219_ (_24740_, _24739_, _24730_);
  nor _29220_ (_24741_, _24740_, _24575_);
  nor _29221_ (_24742_, _24696_, _24589_);
  not _29222_ (_24743_, _24742_);
  not _29223_ (_24744_, _24740_);
  nor _29224_ (_24745_, _24744_, _24137_);
  nor _29225_ (_24746_, _24745_, _24743_);
  not _29226_ (_24747_, _24746_);
  nor _29227_ (_24748_, _24747_, _24741_);
  nor _29228_ (_24749_, _24498_, _24576_);
  nor _29229_ (_24750_, _24696_, _24688_);
  not _29230_ (_24751_, _24750_);
  nor _29231_ (_24752_, _24497_, _24575_);
  nor _29232_ (_24753_, _24752_, _24751_);
  not _29233_ (_24754_, _24753_);
  nor _29234_ (_24755_, _24754_, _24749_);
  nor _29235_ (_24756_, _24755_, _24748_);
  nor _29236_ (_24757_, _24680_, _24579_);
  not _29237_ (_24758_, _24677_);
  nor _29238_ (_24759_, _24758_, _24577_);
  nor _29239_ (_24760_, _24759_, _24757_);
  not _29240_ (_24761_, _24150_);
  nor _29241_ (_24762_, _24690_, _24761_);
  not _29242_ (_24763_, _24670_);
  nor _29243_ (_24764_, _24763_, _24575_);
  nor _29244_ (_24765_, _24764_, _24762_);
  nand _29245_ (_24766_, _24765_, _24760_);
  nor _29246_ (_24767_, _24667_, _24649_);
  not _29247_ (_24768_, _24767_);
  nor _29248_ (_24769_, _24087_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  nor _29249_ (_24770_, _24688_, _24082_);
  nor _29250_ (_24771_, _24770_, _24769_);
  nand _29251_ (_24772_, _24771_, _24768_);
  nor _29252_ (_24773_, _24696_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not _29253_ (_24774_, _24773_);
  nor _29254_ (_24775_, _24676_, _24586_);
  nor _29255_ (_24776_, _24775_, _24668_);
  nand _29256_ (_24777_, _24776_, _24774_);
  nor _29257_ (_24778_, _24777_, _24772_);
  nor _29258_ (_24779_, _24778_, _24137_);
  nor _29259_ (_24780_, _24779_, _24766_);
  nand _29260_ (_24782_, _24780_, _24756_);
  nand _29261_ (_24783_, _24782_, _23939_);
  nand _29262_ (_24784_, _24718_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor _29263_ (_24785_, _24118_, _23939_);
  nand _29264_ (_24786_, _24785_, _24784_);
  nand _29265_ (_24787_, _24786_, _24783_);
  nor _29266_ (_24788_, _24787_, _24722_);
  nor _29267_ (_24789_, _24788_, _23918_);
  nand _29268_ (_24790_, _24789_, _24074_);
  nand _29269_ (_09169_, _24790_, _24076_);
  not _29270_ (_24791_, _23999_);
  nor _29271_ (_24792_, _24791_, _23961_);
  not _29272_ (_24793_, _24792_);
  nor _29273_ (_24794_, _24793_, _24057_);
  not _29274_ (_24795_, _24794_);
  nor _29275_ (_24796_, _24795_, _24073_);
  not _29276_ (_24797_, _24796_);
  nand _29277_ (_24798_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  nor _29278_ (_24799_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], _23939_);
  not _29279_ (_24801_, _24799_);
  nor _29280_ (_24802_, _24801_, _24460_);
  not _29281_ (_24803_, _24802_);
  nor _29282_ (_24804_, _24803_, _24717_);
  nor _29283_ (_24805_, _24758_, _24509_);
  nor _29284_ (_24806_, _24680_, _24511_);
  nor _29285_ (_24807_, _24806_, _24805_);
  not _29286_ (_24808_, _24807_);
  nor _29287_ (_24809_, _24690_, _24436_);
  nor _29288_ (_24810_, _24763_, _24427_);
  nor _29289_ (_24811_, _24810_, _24809_);
  nor _29290_ (_24813_, _24751_, _24434_);
  nor _29291_ (_24814_, _24743_, _24427_);
  nor _29292_ (_24815_, _24814_, _24813_);
  not _29293_ (_24816_, _24815_);
  nor _29294_ (_24817_, _24778_, _24428_);
  nor _29295_ (_24818_, _24817_, _24816_);
  nand _29296_ (_24819_, _24818_, _24811_);
  nor _29297_ (_24820_, _24819_, _24808_);
  not _29298_ (_24821_, _24820_);
  nor _29299_ (_24822_, _24821_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _29300_ (_24823_, _24501_, _23939_);
  nor _29301_ (_24824_, _24823_, _24802_);
  not _29302_ (_24826_, _24824_);
  nor _29303_ (_24827_, _24826_, _24822_);
  nor _29304_ (_24829_, _24827_, _24804_);
  nor _29305_ (_24830_, _24829_, _23918_);
  nand _29306_ (_24831_, _24830_, _24796_);
  nand _29307_ (_16578_, _24831_, _24798_);
  nor _29308_ (_24832_, _24060_, _23979_);
  not _29309_ (_24833_, _24832_);
  nor _29310_ (_24835_, _24069_, _23940_);
  not _29311_ (_24836_, _24835_);
  nor _29312_ (_24837_, _24836_, _24833_);
  not _29313_ (_24838_, _24837_);
  nand _29314_ (_24839_, _24051_, _23996_);
  nor _29315_ (_24840_, _24839_, _23958_);
  not _29316_ (_24842_, _24840_);
  nor _29317_ (_24843_, _24842_, _23938_);
  not _29318_ (_24845_, _24843_);
  nor _29319_ (_24846_, _24845_, _24838_);
  not _29320_ (_24848_, _24846_);
  nor _29321_ (_24849_, _23871_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not _29322_ (_24850_, _24849_);
  nor _29323_ (_24852_, _24850_, _24848_);
  nand _29324_ (_24853_, _24852_, _24830_);
  not _29325_ (_24855_, _24852_);
  nand _29326_ (_24856_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nand _29327_ (_23481_, _24856_, _24853_);
  not _29328_ (_24858_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _29329_ (_24859_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nand _29330_ (_24860_, _24859_, _24858_);
  nor _29331_ (_24861_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  not _29332_ (_24862_, _24861_);
  nor _29333_ (_24863_, _24862_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29334_ (_24864_, _24863_);
  nor _29335_ (_24865_, _24864_, _24860_);
  nand _29336_ (_24866_, _24865_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  nor _29337_ (_24867_, _24866_, _24095_);
  not _29338_ (_24868_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _29339_ (_24869_, _24866_);
  nor _29340_ (_24870_, _24869_, _24868_);
  nor _29341_ (_24871_, _24870_, _24867_);
  nor _29342_ (_28204_[15], _24871_, rst);
  nor _29343_ (_24872_, _24866_, _24868_);
  not _29344_ (_24873_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _29345_ (_24874_, _24869_, _24873_);
  nor _29346_ (_24876_, _24874_, _24872_);
  nor _29347_ (_28205_[15], _24876_, rst);
  nor _29348_ (_24877_, _24054_, _24020_);
  not _29349_ (_24878_, _24877_);
  nor _29350_ (_24881_, _24878_, _24793_);
  not _29351_ (_24882_, _24881_);
  nor _29352_ (_24883_, _24065_, _24063_);
  not _29353_ (_24884_, _24883_);
  nand _29354_ (_24885_, _24069_, _23942_);
  nor _29355_ (_24886_, _24885_, _23918_);
  nand _29356_ (_24887_, _24886_, _23915_);
  nor _29357_ (_24888_, _24887_, _24884_);
  not _29358_ (_24889_, _24888_);
  nor _29359_ (_24890_, _24889_, _24882_);
  nand _29360_ (_24891_, _24719_, _24454_);
  nor _29361_ (_24892_, _24891_, _24717_);
  nor _29362_ (_24893_, _24498_, _24194_);
  nor _29363_ (_24894_, _24497_, _24179_);
  nor _29364_ (_24895_, _24894_, _24893_);
  nor _29365_ (_24896_, _24895_, _24751_);
  nor _29366_ (_24897_, _24727_, _24498_);
  nand _29367_ (_24898_, _24735_, _24498_);
  not _29368_ (_24899_, _24898_);
  nor _29369_ (_24900_, _24899_, _24897_);
  not _29370_ (_24902_, _24900_);
  nor _29371_ (_24903_, _24902_, _24179_);
  nor _29372_ (_24904_, _24900_, _24196_);
  nor _29373_ (_24905_, _24904_, _24743_);
  not _29374_ (_24906_, _24905_);
  nor _29375_ (_24907_, _24906_, _24903_);
  nor _29376_ (_24908_, _24907_, _24896_);
  nor _29377_ (_24909_, _24680_, _24562_);
  nor _29378_ (_24910_, _24758_, _24200_);
  nor _29379_ (_24911_, _24910_, _24909_);
  nand _29380_ (_24912_, _24689_, _24195_);
  not _29381_ (_24913_, _24912_);
  nor _29382_ (_24914_, _24763_, _24196_);
  nor _29383_ (_24916_, _24914_, _24913_);
  nand _29384_ (_24917_, _24916_, _24911_);
  nor _29385_ (_24918_, _24778_, _24179_);
  nor _29386_ (_24919_, _24918_, _24917_);
  nand _29387_ (_24920_, _24919_, _24908_);
  nand _29388_ (_24921_, _24920_, _23939_);
  nand _29389_ (_24922_, _24454_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor _29390_ (_24923_, _24184_, _23939_);
  nand _29391_ (_24924_, _24923_, _24922_);
  nand _29392_ (_24925_, _24924_, _24921_);
  nor _29393_ (_24926_, _24925_, _24892_);
  nor _29394_ (_24927_, _24926_, _23918_);
  nand _29395_ (_24928_, _24927_, _24890_);
  not _29396_ (_24929_, _24890_);
  nand _29397_ (_24930_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  nand _29398_ (_23753_, _24930_, _24928_);
  nand _29399_ (_24931_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _29400_ (_24933_, _24931_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _29401_ (_24934_, _24933_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not _29402_ (_24935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not _29403_ (_24936_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not _29404_ (_24938_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _29405_ (_24939_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _24938_);
  nand _29406_ (_24940_, _24939_, _24936_);
  nor _29407_ (_24941_, _24940_, _24935_);
  not _29408_ (_24942_, _24941_);
  nand _29409_ (_24944_, _24942_, _24934_);
  not _29410_ (_24945_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _29411_ (_24946_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _29412_ (_24947_, _24946_, _24936_);
  not _29413_ (_24949_, _24947_);
  nor _29414_ (_24950_, _24949_, _24945_);
  not _29415_ (_24951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand _29416_ (_24953_, _24946_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _29417_ (_24954_, _24953_, _24951_);
  nor _29418_ (_24955_, _24954_, _24950_);
  not _29419_ (_24956_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _29420_ (_24957_, _24946_, _24936_);
  nor _29421_ (_24958_, _24957_, _24956_);
  not _29422_ (_24959_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  not _29423_ (_24960_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _29424_ (_24961_, _24960_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _29425_ (_24962_, _24961_, _24936_);
  nor _29426_ (_24963_, _24962_, _24959_);
  nor _29427_ (_24964_, _24963_, _24958_);
  nand _29428_ (_24965_, _24964_, _24955_);
  nor _29429_ (_24966_, _24965_, _24944_);
  nor _29430_ (_24968_, _24966_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _29431_ (_24969_, _24968_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _29432_ (_24970_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _29433_ (_24971_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _24970_);
  nor _29434_ (_24972_, _24971_, _24969_);
  not _29435_ (_24973_, _24972_);
  nor _29436_ (_28182_[6], _24973_, rst);
  nor _29437_ (_24975_, _23999_, _23961_);
  not _29438_ (_24976_, _24975_);
  nor _29439_ (_24977_, _24976_, _24057_);
  not _29440_ (_24978_, _24977_);
  not _29441_ (_24979_, _24066_);
  nor _29442_ (_24981_, _24979_, _24062_);
  not _29443_ (_24982_, _24981_);
  nor _29444_ (_24983_, _24887_, _24982_);
  not _29445_ (_24984_, _24983_);
  nor _29446_ (_24985_, _24984_, _24978_);
  nand _29447_ (_24986_, _24985_, _24789_);
  not _29448_ (_24987_, _24985_);
  nand _29449_ (_24988_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nand _29450_ (_24720_, _24988_, _24986_);
  nor _29451_ (_24989_, _23918_, _23915_);
  nor _29452_ (_24990_, _24886_, _24989_);
  not _29453_ (_24991_, _24990_);
  nor _29454_ (_24992_, _24991_, _24982_);
  not _29455_ (_24993_, _24992_);
  nor _29456_ (_24994_, _24054_, _24021_);
  not _29457_ (_24995_, _24994_);
  nor _29458_ (_24996_, _24791_, _23962_);
  not _29459_ (_24997_, _24996_);
  nor _29460_ (_24998_, _24997_, _24995_);
  not _29461_ (_24999_, _24998_);
  nor _29462_ (_25000_, _24999_, _24993_);
  not _29463_ (_25001_, _24719_);
  nor _29464_ (_25002_, _25001_, _24460_);
  nand _29465_ (_25003_, _25002_, _24716_);
  nor _29466_ (_25004_, _24497_, _24224_);
  nor _29467_ (_25005_, _24498_, _24241_);
  nor _29468_ (_25006_, _25005_, _25004_);
  nor _29469_ (_25007_, _25006_, _24751_);
  not _29470_ (_25008_, _24733_);
  nor _29471_ (_25009_, _25008_, _24497_);
  nor _29472_ (_25010_, _24725_, _24498_);
  nor _29473_ (_25011_, _25010_, _25009_);
  nor _29474_ (_25012_, _25011_, _24243_);
  nand _29475_ (_25013_, _25011_, _24243_);
  nand _29476_ (_25014_, _25013_, _24742_);
  nor _29477_ (_25015_, _25014_, _25012_);
  nor _29478_ (_25017_, _25015_, _25007_);
  nor _29479_ (_25018_, _24680_, _24250_);
  nor _29480_ (_25020_, _24758_, _24248_);
  nor _29481_ (_25021_, _25020_, _25018_);
  nor _29482_ (_25022_, _24690_, _24563_);
  nor _29483_ (_25023_, _24763_, _24243_);
  nor _29484_ (_25024_, _25023_, _25022_);
  nand _29485_ (_25025_, _25024_, _25021_);
  nor _29486_ (_25026_, _24778_, _24224_);
  nor _29487_ (_25027_, _25026_, _25025_);
  nand _29488_ (_25028_, _25027_, _25017_);
  not _29489_ (_25029_, _25028_);
  nor _29490_ (_25030_, _25029_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _29491_ (_25031_, _24460_, _24452_);
  nor _29492_ (_25032_, _24229_, _23939_);
  not _29493_ (_25033_, _25032_);
  nor _29494_ (_25034_, _25033_, _25031_);
  nor _29495_ (_25036_, _25034_, _25030_);
  nand _29496_ (_25037_, _25036_, _25003_);
  not _29497_ (_25038_, _25037_);
  nor _29498_ (_25039_, _25038_, _23918_);
  nand _29499_ (_25040_, _25039_, _25000_);
  not _29500_ (_25042_, _25000_);
  nand _29501_ (_25043_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nand _29502_ (_24781_, _25043_, _25040_);
  nor _29503_ (_25044_, _24055_, _24020_);
  not _29504_ (_25045_, _25044_);
  nor _29505_ (_25046_, _25045_, _24793_);
  not _29506_ (_25047_, _25046_);
  nor _29507_ (_25048_, _24016_, _23915_);
  not _29508_ (_25049_, _25048_);
  nor _29509_ (_25050_, _25049_, _24068_);
  not _29510_ (_25051_, _25050_);
  nor _29511_ (_25052_, _25051_, _25047_);
  not _29512_ (_25053_, _25052_);
  nand _29513_ (_25054_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  nand _29514_ (_25055_, _25052_, _24789_);
  nand _29515_ (_24812_, _25055_, _25054_);
  nor _29516_ (_25056_, _24995_, _24793_);
  not _29517_ (_25057_, _25056_);
  nor _29518_ (_25058_, _24884_, _24991_);
  not _29519_ (_25059_, _25058_);
  nor _29520_ (_25061_, _25059_, _25057_);
  nand _29521_ (_25062_, _24799_, _24454_);
  nor _29522_ (_25063_, _25062_, _24717_);
  nor _29523_ (_25065_, _24751_, _24396_);
  not _29524_ (_25066_, _25065_);
  not _29525_ (_25067_, _24731_);
  nor _29526_ (_25068_, _24723_, _25067_);
  not _29527_ (_25069_, _25068_);
  nor _29528_ (_25070_, _25069_, _24498_);
  nor _29529_ (_25071_, _25068_, _24497_);
  nor _29530_ (_25072_, _25071_, _25070_);
  nand _29531_ (_25073_, _25072_, _24742_);
  nand _29532_ (_25074_, _25073_, _25066_);
  nor _29533_ (_25075_, _24778_, _24381_);
  not _29534_ (_25076_, _25075_);
  nor _29535_ (_25078_, _24680_, _24442_);
  nor _29536_ (_25079_, _24758_, _24440_);
  not _29537_ (_25080_, _25079_);
  nand _29538_ (_25081_, _24689_, _24397_);
  not _29539_ (_25082_, _25081_);
  nor _29540_ (_25083_, _24763_, _24380_);
  nor _29541_ (_25084_, _25083_, _25082_);
  nand _29542_ (_25085_, _25084_, _25080_);
  nor _29543_ (_25086_, _25085_, _25078_);
  nand _29544_ (_25087_, _25086_, _25076_);
  nor _29545_ (_25088_, _25087_, _25074_);
  not _29546_ (_25089_, _25088_);
  nand _29547_ (_25091_, _25089_, _23939_);
  nand _29548_ (_25092_, _24799_, _24453_);
  nor _29549_ (_25093_, _24801_, _24463_);
  nor _29550_ (_25094_, _25093_, _24719_);
  nand _29551_ (_25095_, _25094_, _25092_);
  nand _29552_ (_25096_, _25095_, _24359_);
  nand _29553_ (_25097_, _25096_, _25091_);
  nor _29554_ (_25098_, _25097_, _25063_);
  nor _29555_ (_25099_, _25098_, _23918_);
  nand _29556_ (_25101_, _25099_, _25061_);
  not _29557_ (_25102_, _25061_);
  nand _29558_ (_25103_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  nand _29559_ (_24847_, _25103_, _25101_);
  nand _29560_ (_25104_, _25039_, _24890_);
  nand _29561_ (_25106_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nand _29562_ (_24879_, _25106_, _25104_);
  nand _29563_ (_25107_, _25061_, _24830_);
  nand _29564_ (_25108_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  nand _29565_ (_24901_, _25108_, _25107_);
  nand _29566_ (_25109_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nor _29567_ (_25110_, _25001_, _24470_);
  nand _29568_ (_25111_, _25110_, _24716_);
  nor _29569_ (_25112_, _24736_, _24557_);
  nor _29570_ (_25113_, _25112_, _24738_);
  not _29571_ (_25114_, _24729_);
  nand _29572_ (_25115_, _24728_, _24557_);
  nand _29573_ (_25116_, _25115_, _25114_);
  nand _29574_ (_25118_, _25116_, _24497_);
  not _29575_ (_25119_, _25118_);
  nor _29576_ (_25121_, _25119_, _25113_);
  nor _29577_ (_25122_, _25121_, _24743_);
  nor _29578_ (_25123_, _24555_, _24498_);
  nor _29579_ (_25125_, _24549_, _24497_);
  nor _29580_ (_25126_, _25125_, _25123_);
  nor _29581_ (_25127_, _25126_, _24751_);
  nor _29582_ (_25128_, _25127_, _25122_);
  nor _29583_ (_25129_, _24680_, _24561_);
  nor _29584_ (_25130_, _24758_, _24559_);
  nor _29585_ (_25131_, _25130_, _25129_);
  nand _29586_ (_25132_, _24689_, _24556_);
  not _29587_ (_25133_, _25132_);
  nor _29588_ (_25134_, _24763_, _24557_);
  nor _29589_ (_25135_, _25134_, _25133_);
  nand _29590_ (_25136_, _25135_, _25131_);
  nor _29591_ (_25137_, _24778_, _24549_);
  nor _29592_ (_25138_, _25137_, _25136_);
  nand _29593_ (_25139_, _25138_, _25128_);
  not _29594_ (_25140_, _25139_);
  nor _29595_ (_25141_, _25140_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _29596_ (_25143_, _24470_, _24452_);
  nor _29597_ (_25144_, _24469_, _23939_);
  not _29598_ (_25145_, _25144_);
  nor _29599_ (_25146_, _25145_, _25143_);
  nor _29600_ (_25147_, _25146_, _25141_);
  nand _29601_ (_25148_, _25147_, _25111_);
  not _29602_ (_25149_, _25148_);
  nor _29603_ (_25150_, _25149_, _23918_);
  nand _29604_ (_25151_, _25150_, _25052_);
  nand _29605_ (_24932_, _25151_, _25109_);
  nor _29606_ (_25152_, _24993_, _24795_);
  nand _29607_ (_25153_, _25152_, _25039_);
  not _29608_ (_25154_, _25152_);
  nand _29609_ (_25155_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nand _29610_ (_25328_, _25155_, _25153_);
  nor _29611_ (_25156_, _24066_, _24062_);
  not _29612_ (_25157_, _25156_);
  nor _29613_ (_25158_, _25157_, _24991_);
  not _29614_ (_25159_, _25158_);
  nor _29615_ (_25160_, _25159_, _24999_);
  nand _29616_ (_25161_, _25160_, _24789_);
  not _29617_ (_25162_, _25160_);
  nand _29618_ (_25163_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nand _29619_ (_25419_, _25163_, _25161_);
  nor _29620_ (_25164_, _24884_, _24071_);
  not _29621_ (_25165_, _25164_);
  nor _29622_ (_25166_, _25165_, _24882_);
  nand _29623_ (_25167_, _25166_, _24927_);
  not _29624_ (_25168_, _25166_);
  nand _29625_ (_25169_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  nand _29626_ (_25521_, _25169_, _25167_);
  nand _29627_ (_25170_, _25093_, _24716_);
  nor _29628_ (_25171_, _24680_, _24618_);
  nor _29629_ (_25172_, _24758_, _24297_);
  nor _29630_ (_25173_, _25172_, _25171_);
  nand _29631_ (_25174_, _24689_, _24286_);
  not _29632_ (_25175_, _25174_);
  nor _29633_ (_25176_, _24763_, _24278_);
  nor _29634_ (_25177_, _25176_, _25175_);
  nand _29635_ (_25178_, _25177_, _25173_);
  not _29636_ (_25179_, _25178_);
  nor _29637_ (_25180_, _24778_, _24279_);
  nor _29638_ (_25181_, _24732_, _24278_);
  not _29639_ (_25182_, _25181_);
  nand _29640_ (_25183_, _25182_, _25009_);
  nand _29641_ (_25185_, _24724_, _24278_);
  nand _29642_ (_25186_, _25185_, _24726_);
  nand _29643_ (_25187_, _25186_, _24497_);
  nand _29644_ (_25188_, _25187_, _25183_);
  nand _29645_ (_25189_, _25188_, _24742_);
  nor _29646_ (_25190_, _24751_, _24285_);
  not _29647_ (_25191_, _25190_);
  nand _29648_ (_25192_, _25191_, _25189_);
  nor _29649_ (_25193_, _25192_, _25180_);
  nand _29650_ (_25194_, _25193_, _25179_);
  not _29651_ (_25195_, _25194_);
  nor _29652_ (_25196_, _25195_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _29653_ (_25197_, _24463_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _29654_ (_25198_, _24290_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _29655_ (_25199_, _25198_, _25197_);
  nor _29656_ (_25200_, _25199_, _25196_);
  nand _29657_ (_25201_, _25200_, _25170_);
  not _29658_ (_25202_, _25201_);
  nor _29659_ (_25203_, _25202_, _23918_);
  nand _29660_ (_25204_, _25203_, _25160_);
  nand _29661_ (_25205_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand _29662_ (_25917_, _25205_, _25204_);
  nand _29663_ (_25206_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29664_ (_25207_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _29665_ (_25208_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _29666_ (_25209_, _24949_, _25208_);
  not _29667_ (_25210_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _29668_ (_25212_, _24940_, _25210_);
  nor _29669_ (_25213_, _25212_, _25209_);
  nand _29670_ (_25214_, _24933_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  not _29671_ (_25215_, _24962_);
  nand _29672_ (_25216_, _25215_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nand _29673_ (_25217_, _25216_, _25214_);
  not _29674_ (_25218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _29675_ (_25219_, _24957_, _25218_);
  not _29676_ (_25220_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _29677_ (_25222_, _24953_, _25220_);
  nor _29678_ (_25223_, _25222_, _25219_);
  not _29679_ (_25224_, _25223_);
  nor _29680_ (_25225_, _25224_, _25217_);
  nand _29681_ (_25226_, _25225_, _25213_);
  nand _29682_ (_25227_, _25226_, _25207_);
  nand _29683_ (_25228_, _25227_, _24970_);
  nor _29684_ (_25229_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _24970_);
  not _29685_ (_25230_, _25229_);
  nand _29686_ (_25231_, _25230_, _25228_);
  nand _29687_ (_25232_, _25231_, _24865_);
  nor _29688_ (_25233_, _24863_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _29689_ (_25234_, _25233_, _24860_);
  nand _29690_ (_25235_, _25234_, _25232_);
  not _29691_ (_25236_, _25235_);
  not _29692_ (_25237_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _29693_ (_25238_, _24949_, _25237_);
  not _29694_ (_25239_, _25238_);
  not _29695_ (_25240_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _29696_ (_25241_, _24953_, _25240_);
  not _29697_ (_25242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  not _29698_ (_25243_, _24933_);
  nor _29699_ (_25244_, _25243_, _25242_);
  nor _29700_ (_25245_, _25244_, _25241_);
  nand _29701_ (_25246_, _25245_, _25239_);
  not _29702_ (_25248_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _29703_ (_25249_, _24957_, _25248_);
  not _29704_ (_25250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _29705_ (_25251_, _24940_, _25250_);
  nor _29706_ (_25252_, _25251_, _25249_);
  not _29707_ (_25253_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _29708_ (_25254_, _24962_, _25253_);
  nor _29709_ (_25255_, _25254_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _29710_ (_25256_, _25255_, _25252_);
  nor _29711_ (_25258_, _25256_, _25246_);
  nand _29712_ (_25259_, _25258_, _24970_);
  nor _29713_ (_25260_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _24970_);
  not _29714_ (_25261_, _25260_);
  nand _29715_ (_25262_, _25261_, _25259_);
  nand _29716_ (_25263_, _25262_, _24865_);
  nor _29717_ (_25264_, _24863_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _29718_ (_25265_, _25264_, _24860_);
  nand _29719_ (_25266_, _25265_, _25263_);
  not _29720_ (_25267_, _25266_);
  not _29721_ (_25268_, _24865_);
  not _29722_ (_25269_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _29723_ (_25270_, _24957_, _25269_);
  not _29724_ (_25271_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _29725_ (_25272_, _24962_, _25271_);
  nor _29726_ (_25273_, _25272_, _25270_);
  not _29727_ (_25274_, _25273_);
  nand _29728_ (_25275_, _24947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  not _29729_ (_25276_, _25275_);
  not _29730_ (_25277_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _29731_ (_25278_, _24953_, _25277_);
  nor _29732_ (_25279_, _25278_, _25276_);
  nand _29733_ (_25280_, _24933_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  not _29734_ (_25281_, _25280_);
  not _29735_ (_25282_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _29736_ (_25283_, _24940_, _25282_);
  nor _29737_ (_25284_, _25283_, _25281_);
  nand _29738_ (_25285_, _25284_, _25279_);
  nor _29739_ (_25286_, _25285_, _25274_);
  nor _29740_ (_25287_, _25286_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _29741_ (_25288_, _25287_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _29742_ (_25289_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _24970_);
  nor _29743_ (_25290_, _25289_, _25288_);
  nor _29744_ (_25291_, _25290_, _25268_);
  nor _29745_ (_25292_, _24863_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _29746_ (_25293_, _25292_, _24860_);
  not _29747_ (_25294_, _25293_);
  nor _29748_ (_25295_, _25294_, _25291_);
  nand _29749_ (_25296_, _25295_, _25267_);
  nor _29750_ (_25297_, _25296_, _25236_);
  not _29751_ (_25298_, _25297_);
  not _29752_ (_25299_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _29753_ (_25300_, _24949_, _25299_);
  not _29754_ (_25301_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _29755_ (_25303_, _24953_, _25301_);
  not _29756_ (_25304_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _29757_ (_25305_, _25243_, _25304_);
  nor _29758_ (_25306_, _25305_, _25303_);
  not _29759_ (_25307_, _25306_);
  nor _29760_ (_25308_, _25307_, _25300_);
  not _29761_ (_25309_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _29762_ (_25310_, _24957_, _25309_);
  not _29763_ (_25311_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _29764_ (_25312_, _24940_, _25311_);
  nor _29765_ (_25313_, _25312_, _25310_);
  not _29766_ (_25314_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _29767_ (_25315_, _24962_, _25314_);
  nor _29768_ (_25316_, _25315_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _29769_ (_25317_, _25316_, _25313_);
  not _29770_ (_25318_, _25317_);
  nand _29771_ (_25319_, _25318_, _25308_);
  nor _29772_ (_25320_, _25319_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _29773_ (_25321_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _24970_);
  nor _29774_ (_25322_, _25321_, _25320_);
  nor _29775_ (_25323_, _25322_, _25268_);
  nor _29776_ (_25324_, _24863_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _29777_ (_25325_, _25324_, _24860_);
  not _29778_ (_25326_, _25325_);
  nor _29779_ (_25327_, _25326_, _25323_);
  not _29780_ (_25329_, _25327_);
  not _29781_ (_25330_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _29782_ (_25331_, _24940_, _25330_);
  not _29783_ (_25332_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _29784_ (_25333_, _24962_, _25332_);
  nor _29785_ (_25334_, _25333_, _25331_);
  not _29786_ (_25335_, _25334_);
  not _29787_ (_25336_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _29788_ (_25337_, _24949_, _25336_);
  not _29789_ (_25338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _29790_ (_25339_, _24953_, _25338_);
  nor _29791_ (_25340_, _25339_, _25337_);
  not _29792_ (_25341_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _29793_ (_25342_, _24957_, _25341_);
  not _29794_ (_25343_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _29795_ (_25344_, _25243_, _25343_);
  nor _29796_ (_25345_, _25344_, _25342_);
  nand _29797_ (_25346_, _25345_, _25340_);
  nor _29798_ (_25347_, _25346_, _25335_);
  nor _29799_ (_25348_, _25347_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _29800_ (_25349_, _25348_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _29801_ (_25350_, _24970_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nor _29802_ (_25351_, _25350_, _25349_);
  nor _29803_ (_25352_, _25351_, _25268_);
  nor _29804_ (_25353_, _24863_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _29805_ (_25354_, _25353_, _24860_);
  not _29806_ (_25355_, _25354_);
  nor _29807_ (_25356_, _25355_, _25352_);
  nor _29808_ (_25357_, _24972_, _25268_);
  nor _29809_ (_25358_, _24863_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _29810_ (_25359_, _25358_, _24860_);
  not _29811_ (_25360_, _25359_);
  nor _29812_ (_25361_, _25360_, _25357_);
  not _29813_ (_25362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _29814_ (_25363_, _24962_, _25362_);
  not _29815_ (_25364_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _29816_ (_25365_, _24940_, _25364_);
  nor _29817_ (_25366_, _25365_, _25363_);
  not _29818_ (_25367_, _25366_);
  nand _29819_ (_25368_, _24947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not _29820_ (_25369_, _25368_);
  not _29821_ (_25370_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _29822_ (_25371_, _24953_, _25370_);
  nor _29823_ (_25372_, _25371_, _25369_);
  not _29824_ (_25373_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _29825_ (_25374_, _24957_, _25373_);
  nand _29826_ (_25375_, _24933_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not _29827_ (_25376_, _25375_);
  nor _29828_ (_25377_, _25376_, _25374_);
  nand _29829_ (_25378_, _25377_, _25372_);
  nor _29830_ (_25379_, _25378_, _25367_);
  nor _29831_ (_25380_, _25379_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _29832_ (_25381_, _25380_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _29833_ (_25382_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _24970_);
  nor _29834_ (_25383_, _25382_, _25381_);
  nor _29835_ (_25384_, _25383_, _25268_);
  nor _29836_ (_25385_, _24863_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _29837_ (_25386_, _25385_, _24860_);
  not _29838_ (_25387_, _25386_);
  nor _29839_ (_25388_, _25387_, _25384_);
  not _29840_ (_25389_, _25388_);
  nand _29841_ (_25390_, _25389_, _25361_);
  nor _29842_ (_25391_, _25390_, _25356_);
  not _29843_ (_25392_, _25391_);
  nor _29844_ (_25393_, _25392_, _25329_);
  nor _29845_ (_25394_, _25361_, _25356_);
  nand _29846_ (_25395_, _25394_, _25388_);
  not _29847_ (_25396_, _25395_);
  nor _29848_ (_25397_, _25396_, _25393_);
  nor _29849_ (_25398_, _25397_, _25298_);
  not _29850_ (_25399_, _25398_);
  not _29851_ (_25400_, _25356_);
  nand _29852_ (_25401_, _25388_, _25361_);
  nor _29853_ (_25402_, _25401_, _25400_);
  nand _29854_ (_25403_, _25402_, _25329_);
  nor _29855_ (_25404_, _25403_, _25298_);
  nor _29856_ (_25405_, _25327_, _25236_);
  nor _29857_ (_25406_, _25390_, _25296_);
  nand _29858_ (_25407_, _25406_, _25405_);
  nor _29859_ (_25408_, _25407_, _25356_);
  nor _29860_ (_25409_, _25408_, _25404_);
  nand _29861_ (_25410_, _25409_, _25399_);
  nor _29862_ (_25411_, _25298_, _25329_);
  not _29863_ (_25412_, _25411_);
  not _29864_ (_25413_, _25361_);
  nand _29865_ (_25414_, _25413_, _25356_);
  not _29866_ (_25415_, _25414_);
  nand _29867_ (_25416_, _25415_, _25389_);
  nor _29868_ (_25417_, _25416_, _25412_);
  nor _29869_ (_25418_, _25390_, _25400_);
  not _29870_ (_25420_, _25418_);
  nor _29871_ (_25421_, _25420_, _25298_);
  nor _29872_ (_25422_, _25421_, _25417_);
  nand _29873_ (_25423_, _25394_, _25389_);
  nor _29874_ (_25424_, _25423_, _25298_);
  nor _29875_ (_25425_, _25414_, _25389_);
  nand _29876_ (_25426_, _25425_, _25327_);
  nor _29877_ (_25427_, _25426_, _25298_);
  nor _29878_ (_25428_, _25427_, _25424_);
  nand _29879_ (_25430_, _25428_, _25422_);
  nor _29880_ (_25431_, _25430_, _25410_);
  not _29881_ (_25432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _29882_ (_25433_, _24962_, _25432_);
  not _29883_ (_25434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _29884_ (_25435_, _24940_, _25434_);
  nor _29885_ (_25436_, _25435_, _25433_);
  not _29886_ (_25437_, _25436_);
  nand _29887_ (_25438_, _24947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  not _29888_ (_25439_, _25438_);
  not _29889_ (_25440_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _29890_ (_25441_, _24953_, _25440_);
  nor _29891_ (_25442_, _25441_, _25439_);
  not _29892_ (_25443_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _29893_ (_25444_, _24957_, _25443_);
  nand _29894_ (_25445_, _24933_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not _29895_ (_25446_, _25445_);
  nor _29896_ (_25447_, _25446_, _25444_);
  nand _29897_ (_25448_, _25447_, _25442_);
  nor _29898_ (_25449_, _25448_, _25437_);
  nor _29899_ (_25450_, _25449_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _29900_ (_25451_, _25450_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _29901_ (_25452_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _24970_);
  nor _29902_ (_25453_, _25452_, _25451_);
  nor _29903_ (_25454_, _25453_, _25268_);
  nor _29904_ (_25455_, _24863_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _29905_ (_25456_, _25455_, _24860_);
  not _29906_ (_25457_, _25456_);
  nor _29907_ (_25458_, _25457_, _25454_);
  not _29908_ (_25459_, _25458_);
  not _29909_ (_25460_, _25295_);
  nand _29910_ (_25461_, _25235_, _25460_);
  nor _29911_ (_25462_, _25461_, _25266_);
  not _29912_ (_25463_, _25462_);
  nor _29913_ (_25464_, _25463_, _25459_);
  not _29914_ (_25465_, _25464_);
  nand _29915_ (_25466_, _25425_, _25329_);
  nor _29916_ (_25467_, _25466_, _25465_);
  not _29917_ (_25468_, _25467_);
  nor _29918_ (_25469_, _25416_, _25329_);
  not _29919_ (_25470_, _25469_);
  nor _29920_ (_25471_, _25470_, _25465_);
  nor _29921_ (_25472_, _25401_, _25356_);
  not _29922_ (_25473_, _25472_);
  nor _29923_ (_25474_, _25329_, _25473_);
  not _29924_ (_25475_, _25474_);
  nor _29925_ (_25476_, _25465_, _25475_);
  nor _29926_ (_25477_, _25476_, _25471_);
  nand _29927_ (_25478_, _25477_, _25468_);
  nor _29928_ (_25479_, _25267_, _25458_);
  not _29929_ (_25480_, _25479_);
  nor _29930_ (_25481_, _25461_, _25480_);
  not _29931_ (_25482_, _25481_);
  nand _29932_ (_25483_, _25418_, _25327_);
  nor _29933_ (_25484_, _25483_, _25482_);
  nor _29934_ (_25485_, _25463_, _25458_);
  nand _29935_ (_25486_, _25485_, _25396_);
  not _29936_ (_25487_, _25486_);
  nor _29937_ (_25488_, _25487_, _25484_);
  nor _29938_ (_25489_, _25327_, _25473_);
  not _29939_ (_25490_, _25489_);
  nor _29940_ (_25491_, _25298_, _25490_);
  nor _29941_ (_25492_, _25416_, _25327_);
  not _29942_ (_25493_, _25492_);
  nor _29943_ (_25494_, _25493_, _25298_);
  nor _29944_ (_25495_, _25494_, _25491_);
  nand _29945_ (_25496_, _25495_, _25488_);
  nor _29946_ (_25497_, _25496_, _25478_);
  nand _29947_ (_25498_, _25497_, _25431_);
  nand _29948_ (_25499_, _24862_, _23870_);
  nand _29949_ (_25500_, _25499_, _25498_);
  not _29950_ (_25501_, \oc8051_top_1.oc8051_decoder1.state [1]);
  nor _29951_ (_25502_, _25501_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29952_ (_25503_, _25502_);
  nor _29953_ (_25504_, _25503_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not _29954_ (_25505_, _25504_);
  nor _29955_ (_25506_, _25482_, _25473_);
  not _29956_ (_25507_, _25506_);
  nor _29957_ (_25508_, _25507_, _25505_);
  not _29958_ (_25509_, _25485_);
  nor _29959_ (_25510_, _25395_, _25329_);
  not _29960_ (_25511_, _25510_);
  nor _29961_ (_25512_, _25511_, _25509_);
  nor _29962_ (_25513_, _25395_, _25327_);
  not _29963_ (_25514_, _25513_);
  nor _29964_ (_25515_, _25514_, _25509_);
  nor _29965_ (_25516_, _25515_, _25512_);
  not _29966_ (_25517_, \oc8051_top_1.oc8051_decoder1.state [0]);
  nor _29967_ (_25518_, _25503_, _25517_);
  not _29968_ (_25519_, _25518_);
  nor _29969_ (_25520_, _25519_, _25516_);
  nor _29970_ (_25522_, _25520_, _25508_);
  nand _29971_ (_25523_, _25522_, _25500_);
  nand _29972_ (_25524_, _25523_, _23870_);
  nand _29973_ (_25526_, _25524_, _25206_);
  not _29974_ (_25527_, _25526_);
  nand _29975_ (_25528_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29976_ (_25529_, _25528_);
  not _29977_ (_25530_, _25499_);
  nor _29978_ (_25531_, _25509_, _25466_);
  nor _29979_ (_25532_, _25483_, _25463_);
  nand _29980_ (_25533_, _25532_, _25459_);
  not _29981_ (_25534_, _25533_);
  nor _29982_ (_25535_, _25534_, _25531_);
  nor _29983_ (_25537_, _25511_, _25482_);
  nand _29984_ (_25538_, _25513_, _25481_);
  nor _29985_ (_25540_, _25423_, _25329_);
  nand _29986_ (_25541_, _25540_, _25481_);
  nand _29987_ (_25542_, _25541_, _25538_);
  nor _29988_ (_25544_, _25542_, _25537_);
  not _29989_ (_25545_, _25544_);
  nor _29990_ (_25546_, _25466_, _25235_);
  not _29991_ (_25547_, _25546_);
  nand _29992_ (_25548_, _25235_, _25295_);
  nand _29993_ (_25549_, _25266_, _25458_);
  nor _29994_ (_25550_, _25549_, _25548_);
  not _29995_ (_25551_, _25550_);
  nor _29996_ (_25552_, _25423_, _25327_);
  not _29997_ (_25553_, _25552_);
  nor _29998_ (_25554_, _25553_, _25551_);
  nand _29999_ (_25555_, _25462_, _25489_);
  not _30000_ (_25556_, _25555_);
  nor _30001_ (_25557_, _25556_, _25554_);
  nand _30002_ (_25558_, _25557_, _25547_);
  nor _30003_ (_25559_, _25558_, _25545_);
  nand _30004_ (_25560_, _25559_, _25535_);
  nor _30005_ (_25561_, _25392_, _25327_);
  nand _30006_ (_25562_, _25561_, _25550_);
  not _30007_ (_25563_, _25425_);
  nor _30008_ (_25564_, _25563_, _25482_);
  not _30009_ (_25565_, _25564_);
  nand _30010_ (_25566_, _25565_, _25562_);
  nand _30011_ (_25567_, _25485_, _25474_);
  nand _30012_ (_25568_, _25561_, _25462_);
  nand _30013_ (_25569_, _25568_, _25567_);
  nor _30014_ (_25570_, _25569_, _25566_);
  not _30015_ (_25571_, _25570_);
  not _30016_ (_25572_, _25540_);
  nor _30017_ (_25573_, _25551_, _25572_);
  nor _30018_ (_25574_, _25551_, _25483_);
  nor _30019_ (_25575_, _25574_, _25573_);
  nor _30020_ (_25576_, _25509_, _25426_);
  nand _30021_ (_25577_, _25418_, _25329_);
  nor _30022_ (_25578_, _25577_, _25509_);
  nor _30023_ (_25579_, _25578_, _25576_);
  nand _30024_ (_25580_, _25579_, _25575_);
  nor _30025_ (_25581_, _25580_, _25571_);
  nand _30026_ (_25582_, _25550_, _25489_);
  not _30027_ (_25583_, _25582_);
  nor _30028_ (_25584_, _25577_, _25551_);
  nor _30029_ (_25585_, _25584_, _25583_);
  nor _30030_ (_25586_, _25551_, _25397_);
  nand _30031_ (_25587_, _25485_, _25469_);
  nand _30032_ (_25588_, _25550_, _25492_);
  nand _30033_ (_25589_, _25588_, _25587_);
  nor _30034_ (_25590_, _25589_, _25586_);
  nand _30035_ (_25591_, _25590_, _25585_);
  nand _30036_ (_25592_, _25550_, _25469_);
  nor _30037_ (_25593_, _25551_, _25403_);
  not _30038_ (_25594_, _25593_);
  nand _30039_ (_25595_, _25594_, _25592_);
  not _30040_ (_25596_, _25426_);
  nand _30041_ (_25597_, _25550_, _25596_);
  not _30042_ (_25598_, _25466_);
  nand _30043_ (_25599_, _25598_, _25297_);
  nand _30044_ (_25600_, _25599_, _25597_);
  nor _30045_ (_25601_, _25600_, _25595_);
  nand _30046_ (_25602_, _25492_, _25485_);
  nand _30047_ (_25603_, _25462_, _25393_);
  nand _30048_ (_25604_, _25603_, _25602_);
  nand _30049_ (_25605_, _25418_, _25481_);
  nand _30050_ (_25606_, _25605_, _25486_);
  nor _30051_ (_25607_, _25606_, _25604_);
  nand _30052_ (_25608_, _25607_, _25601_);
  nor _30053_ (_25609_, _25608_, _25591_);
  nand _30054_ (_25610_, _25609_, _25581_);
  nor _30055_ (_25611_, _25610_, _25560_);
  nor _30056_ (_25612_, _25611_, _25530_);
  nor _30057_ (_25613_, _25519_, _25486_);
  not _30058_ (_25614_, _25613_);
  nor _30059_ (_25615_, _25392_, _25482_);
  not _30060_ (_25616_, _25615_);
  nor _30061_ (_25617_, _25616_, _25505_);
  nor _30062_ (_25618_, _25617_, _25508_);
  nand _30063_ (_25619_, _25618_, _25614_);
  nor _30064_ (_25620_, _25619_, _25612_);
  nor _30065_ (_25621_, _25620_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _30066_ (_25622_, _25621_, _25529_);
  nor _30067_ (_25623_, _25622_, _25527_);
  not _30068_ (_25624_, _25623_);
  not _30069_ (_25625_, _24782_);
  nor _30070_ (_25626_, _24060_, _23978_);
  nand _30071_ (_25627_, _25626_, _24070_);
  not _30072_ (_25628_, _25627_);
  nand _30073_ (_25629_, _24840_, _23938_);
  nor _30074_ (_25630_, _24850_, _23875_);
  not _30075_ (_25631_, _25630_);
  nor _30076_ (_25632_, _25631_, _25629_);
  nand _30077_ (_25633_, _25632_, _25628_);
  nor _30078_ (_25634_, _25633_, _25625_);
  not _30079_ (_25635_, _25633_);
  nor _30080_ (_25636_, _25635_, _23876_);
  not _30081_ (_25637_, _25636_);
  nand _30082_ (_25638_, _25635_, _25139_);
  nand _30083_ (_25639_, _25638_, _25637_);
  not _30084_ (_25640_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _30085_ (_25641_, _25635_, _25640_);
  not _30086_ (_25642_, _25641_);
  nand _30087_ (_25643_, _25635_, _24920_);
  nand _30088_ (_25644_, _25643_, _25642_);
  not _30089_ (_25645_, _25644_);
  nor _30090_ (_25646_, _25635_, _23877_);
  not _30091_ (_25647_, _25646_);
  nand _30092_ (_25648_, _25635_, _25028_);
  nand _30093_ (_25649_, _25648_, _25647_);
  nand _30094_ (_25650_, _25633_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  not _30095_ (_25651_, _25650_);
  nor _30096_ (_25652_, _25633_, _25195_);
  nor _30097_ (_25653_, _25652_, _25651_);
  nor _30098_ (_25654_, _25635_, _23878_);
  not _30099_ (_25655_, _25654_);
  nor _30100_ (_25656_, _24751_, _24338_);
  not _30101_ (_25657_, _24723_);
  nand _30102_ (_25658_, _25657_, _24497_);
  not _30103_ (_25659_, _25658_);
  nor _30104_ (_25660_, _25067_, _24497_);
  nor _30105_ (_25661_, _25660_, _25659_);
  nand _30106_ (_25662_, _25661_, _24350_);
  not _30107_ (_25663_, _25660_);
  nand _30108_ (_25664_, _25663_, _25658_);
  nand _30109_ (_25665_, _25664_, _24323_);
  nand _30110_ (_25666_, _25665_, _25662_);
  nor _30111_ (_25668_, _25666_, _24743_);
  nor _30112_ (_25669_, _25668_, _25656_);
  nor _30113_ (_25670_, _24680_, _24356_);
  nor _30114_ (_25671_, _24758_, _24354_);
  nor _30115_ (_25672_, _25671_, _25670_);
  nand _30116_ (_25673_, _24689_, _24339_);
  not _30117_ (_25674_, _25673_);
  nor _30118_ (_25675_, _24763_, _24350_);
  nor _30119_ (_25676_, _25675_, _25674_);
  nand _30120_ (_25677_, _25676_, _25672_);
  nor _30121_ (_25678_, _24778_, _24323_);
  nor _30122_ (_25679_, _25678_, _25677_);
  nand _30123_ (_25680_, _25679_, _25669_);
  nand _30124_ (_25681_, _25680_, _25635_);
  nand _30125_ (_25682_, _25681_, _25655_);
  nor _30126_ (_25683_, _25635_, _23880_);
  nor _30127_ (_25684_, _25633_, _25088_);
  nor _30128_ (_25685_, _25684_, _25683_);
  nor _30129_ (_25686_, _25635_, _23879_);
  nor _30130_ (_25687_, _25633_, _24820_);
  nor _30131_ (_25688_, _25687_, _25686_);
  nand _30132_ (_25689_, _25688_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  not _30133_ (_25690_, _25689_);
  nand _30134_ (_25691_, _25690_, _25685_);
  nor _30135_ (_25692_, _25691_, _25682_);
  nand _30136_ (_25693_, _25692_, _25653_);
  nor _30137_ (_25694_, _25693_, _25649_);
  nand _30138_ (_25695_, _25694_, _25645_);
  nor _30139_ (_25696_, _25695_, _25639_);
  nand _30140_ (_25697_, _25633_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _30141_ (_25698_, _25697_, _25696_);
  not _30142_ (_25699_, _25639_);
  not _30143_ (_25700_, _25649_);
  not _30144_ (_25701_, _25678_);
  nand _30145_ (_25702_, _25701_, _25669_);
  nor _30146_ (_25703_, _25702_, _25677_);
  nor _30147_ (_25704_, _25703_, _25633_);
  nor _30148_ (_25705_, _25704_, _25654_);
  nand _30149_ (_25706_, _25705_, _25653_);
  nor _30150_ (_25707_, _25706_, _25691_);
  nand _30151_ (_25708_, _25707_, _25700_);
  nor _30152_ (_25709_, _25708_, _25644_);
  nand _30153_ (_25710_, _25709_, _25699_);
  not _30154_ (_25711_, _25697_);
  nor _30155_ (_25712_, _25711_, _25710_);
  nor _30156_ (_25713_, _25712_, _25698_);
  nor _30157_ (_25714_, _25713_, _23891_);
  nor _30158_ (_25715_, _25714_, _23894_);
  nor _30159_ (_25716_, _25715_, _25635_);
  nor _30160_ (_25717_, _25716_, _25634_);
  nor _30161_ (_25718_, _25717_, _25624_);
  nand _30162_ (_25719_, _25622_, _25526_);
  not _30163_ (_25720_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  not _30164_ (_25721_, _23958_);
  nor _30165_ (_25722_, _24839_, _25721_);
  not _30166_ (_25723_, _25722_);
  not _30167_ (_25724_, _23938_);
  nor _30168_ (_25725_, _25631_, _25724_);
  not _30169_ (_25726_, _25725_);
  nor _30170_ (_25727_, _25726_, _25723_);
  nand _30171_ (_25728_, _25727_, _25048_);
  nor _30172_ (_25729_, _25728_, _24833_);
  nor _30173_ (_25730_, _25729_, _25720_);
  not _30174_ (_25731_, _25730_);
  nand _30175_ (_25732_, _25729_, _25028_);
  nand _30176_ (_25733_, _25732_, _25731_);
  not _30177_ (_25734_, _25733_);
  nor _30178_ (_25735_, _25734_, _23979_);
  nor _30179_ (_25736_, _25733_, _23978_);
  nor _30180_ (_25737_, _25736_, _25735_);
  not _30181_ (_25738_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _30182_ (_25739_, _25729_, _25738_);
  not _30183_ (_25740_, _25739_);
  nand _30184_ (_25741_, _25729_, _25194_);
  nand _30185_ (_25742_, _25741_, _25740_);
  not _30186_ (_25743_, _25742_);
  nor _30187_ (_25744_, _25743_, _23938_);
  nor _30188_ (_25745_, _25742_, _25724_);
  nor _30189_ (_25746_, _25745_, _25744_);
  nor _30190_ (_25747_, _25458_, _23958_);
  nor _30191_ (_25748_, _25459_, _25721_);
  nor _30192_ (_25749_, _25748_, _25747_);
  not _30193_ (_25750_, _24839_);
  nand _30194_ (_25751_, _24849_, _25750_);
  nor _30195_ (_25752_, _25751_, _24836_);
  nand _30196_ (_25753_, _25752_, _25749_);
  nor _30197_ (_25754_, _25753_, _24060_);
  not _30198_ (_25755_, _25754_);
  nor _30199_ (_25756_, _25755_, _25746_);
  not _30200_ (_25757_, _25756_);
  nor _30201_ (_25758_, _25757_, _25737_);
  not _30202_ (_25759_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _30203_ (_25760_, _25743_, _25458_);
  nand _30204_ (_25761_, _25760_, _25734_);
  nor _30205_ (_25762_, _25761_, _25759_);
  not _30206_ (_25764_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _30207_ (_25765_, _25742_, _25459_);
  nand _30208_ (_25766_, _25765_, _25734_);
  nor _30209_ (_25767_, _25766_, _25764_);
  nor _30210_ (_25768_, _25767_, _25762_);
  not _30211_ (_25769_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor _30212_ (_25770_, _25742_, _25458_);
  nand _30213_ (_25771_, _25770_, _25734_);
  nor _30214_ (_25772_, _25771_, _25769_);
  not _30215_ (_25773_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand _30216_ (_25774_, _25765_, _25733_);
  nor _30217_ (_25775_, _25774_, _25773_);
  nor _30218_ (_25776_, _25775_, _25772_);
  nand _30219_ (_25777_, _25776_, _25768_);
  not _30220_ (_25778_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nand _30221_ (_25779_, _25770_, _25733_);
  nor _30222_ (_25780_, _25779_, _25778_);
  not _30223_ (_25781_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _30224_ (_25782_, _25743_, _25459_);
  nand _30225_ (_25783_, _25782_, _25733_);
  nor _30226_ (_25784_, _25783_, _25781_);
  nor _30227_ (_25785_, _25784_, _25780_);
  not _30228_ (_25786_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand _30229_ (_25787_, _25760_, _25733_);
  nor _30230_ (_25788_, _25787_, _25786_);
  not _30231_ (_25789_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand _30232_ (_25790_, _25782_, _25734_);
  nor _30233_ (_25791_, _25790_, _25789_);
  nor _30234_ (_25792_, _25791_, _25788_);
  nand _30235_ (_25793_, _25792_, _25785_);
  nor _30236_ (_25794_, _25793_, _25777_);
  nor _30237_ (_25795_, _25794_, _25758_);
  nand _30238_ (_25796_, _25758_, _24782_);
  not _30239_ (_25797_, _25796_);
  nor _30240_ (_25798_, _25797_, _25795_);
  nor _30241_ (_25799_, _25798_, _25719_);
  nand _30242_ (_25800_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _30243_ (_25801_, _25800_);
  nor _30244_ (_25802_, _25548_, _25480_);
  not _30245_ (_25803_, _25802_);
  nor _30246_ (_25804_, _25803_, _25493_);
  nor _30247_ (_25805_, _25803_, _25466_);
  nor _30248_ (_25806_, _25805_, _25804_);
  nor _30249_ (_25807_, _25806_, _25499_);
  nor _30250_ (_25808_, _25615_, _25506_);
  nor _30251_ (_25809_, _25808_, _25505_);
  not _30252_ (_25810_, _25809_);
  not _30253_ (_25811_, _25806_);
  nor _30254_ (_25812_, _25811_, _25478_);
  nor _30255_ (_25813_, _25812_, _25530_);
  not _30256_ (_25814_, _25813_);
  nand _30257_ (_25815_, _25814_, _25810_);
  nor _30258_ (_25816_, _25815_, _25807_);
  nor _30259_ (_25817_, _25816_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _30260_ (_25818_, _25817_, _25801_);
  nor _30261_ (_25819_, _25622_, _25526_);
  nor _30262_ (_25820_, _24863_, _23898_);
  nor _30263_ (_25821_, _25243_, _25338_);
  nor _30264_ (_25822_, _24962_, _25343_);
  nor _30265_ (_25823_, _25822_, _25821_);
  not _30266_ (_25824_, _25823_);
  not _30267_ (_25825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _30268_ (_25826_, _24949_, _25825_);
  nor _30269_ (_25827_, _24957_, _25330_);
  nor _30270_ (_25828_, _25827_, _25826_);
  nor _30271_ (_25829_, _24953_, _25336_);
  nor _30272_ (_25830_, _24940_, _25332_);
  nor _30273_ (_25831_, _25830_, _25829_);
  nand _30274_ (_25832_, _25831_, _25828_);
  nor _30275_ (_25833_, _25832_, _25824_);
  nor _30276_ (_25834_, _24864_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _30277_ (_25835_, _25834_);
  nor _30278_ (_25836_, _25835_, _25833_);
  nor _30279_ (_25837_, _25836_, _25820_);
  not _30280_ (_25838_, _25837_);
  nand _30281_ (_25839_, _25838_, _25819_);
  nand _30282_ (_25840_, _25839_, _25818_);
  nor _30283_ (_25841_, _25840_, _25799_);
  not _30284_ (_25842_, _25841_);
  nor _30285_ (_25843_, _25842_, _25718_);
  nor _30286_ (_28206_, _25843_, rst);
  nor _30287_ (_28207_[4], _25734_, rst);
  nor _30288_ (_28208_[7], _25798_, rst);
  nor _30289_ (_25844_, _25517_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _30290_ (_25845_, _25617_, _25545_);
  nor _30291_ (_25846_, _25845_, _25844_);
  not _30292_ (_25847_, _25846_);
  nor _30293_ (_25848_, _25847_, _25809_);
  not _30294_ (_25849_, _25848_);
  not _30295_ (_25850_, _25818_);
  nor _30296_ (_25851_, _25850_, _25719_);
  not _30297_ (_25852_, _25851_);
  not _30298_ (_25853_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _30299_ (_25854_, _25783_, _25853_);
  not _30300_ (_25855_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor _30301_ (_25856_, _25787_, _25855_);
  nor _30302_ (_25857_, _25856_, _25854_);
  not _30303_ (_25858_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _30304_ (_25859_, _25771_, _25858_);
  not _30305_ (_25860_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _30306_ (_25861_, _25779_, _25860_);
  nor _30307_ (_25862_, _25861_, _25859_);
  nand _30308_ (_25863_, _25862_, _25857_);
  not _30309_ (_25864_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _30310_ (_25865_, _25766_, _25864_);
  not _30311_ (_25866_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _30312_ (_25867_, _25790_, _25866_);
  nor _30313_ (_25868_, _25867_, _25865_);
  not _30314_ (_25869_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _30315_ (_25870_, _25761_, _25869_);
  not _30316_ (_25871_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _30317_ (_25872_, _25774_, _25871_);
  nor _30318_ (_25873_, _25872_, _25870_);
  nand _30319_ (_25874_, _25873_, _25868_);
  nor _30320_ (_25876_, _25874_, _25863_);
  nor _30321_ (_25877_, _25876_, _25758_);
  not _30322_ (_25879_, _25758_);
  nor _30323_ (_25880_, _25879_, _25195_);
  nor _30324_ (_25881_, _25880_, _25877_);
  nor _30325_ (_25882_, _25881_, _25852_);
  nand _30326_ (_25883_, _25622_, _25527_);
  nor _30327_ (_25884_, _25883_, _25850_);
  nand _30328_ (_25885_, _25884_, _25742_);
  nand _30329_ (_25886_, _25818_, _25623_);
  nor _30330_ (_25887_, _25692_, _25653_);
  nor _30331_ (_25888_, _25887_, _25707_);
  nor _30332_ (_25889_, _25888_, _23891_);
  nor _30333_ (_25890_, _25889_, _23921_);
  nor _30334_ (_25891_, _25890_, _25635_);
  nor _30335_ (_25892_, _25891_, _25652_);
  nor _30336_ (_25893_, _25892_, _25886_);
  nand _30337_ (_25894_, _25819_, _25818_);
  nor _30338_ (_25895_, _24863_, _23922_);
  nor _30339_ (_25896_, _25243_, _25220_);
  not _30340_ (_25897_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _30341_ (_25898_, _24962_, _25897_);
  nor _30342_ (_25899_, _25898_, _25896_);
  not _30343_ (_25900_, _25899_);
  not _30344_ (_25901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _30345_ (_25902_, _24949_, _25901_);
  not _30346_ (_25903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _30347_ (_25904_, _24940_, _25903_);
  nor _30348_ (_25905_, _25904_, _25902_);
  nor _30349_ (_25906_, _24957_, _25210_);
  nor _30350_ (_25907_, _24953_, _25208_);
  nor _30351_ (_25908_, _25907_, _25906_);
  nand _30352_ (_25909_, _25908_, _25905_);
  nor _30353_ (_25910_, _25909_, _25900_);
  nor _30354_ (_25911_, _25910_, _25835_);
  nor _30355_ (_25912_, _25911_, _25895_);
  nor _30356_ (_25913_, _25912_, _25894_);
  nor _30357_ (_25914_, _25913_, _25893_);
  nand _30358_ (_25915_, _25914_, _25885_);
  nor _30359_ (_25916_, _25915_, _25882_);
  nor _30360_ (_25918_, _25916_, _23938_);
  not _30361_ (_25919_, _25916_);
  nor _30362_ (_25920_, _25919_, _25724_);
  nor _30363_ (_25921_, _25920_, _25918_);
  nor _30364_ (_25922_, _25843_, _23915_);
  nor _30365_ (_25923_, _25633_, _24782_);
  nor _30366_ (_25924_, _25635_, _23894_);
  not _30367_ (_25925_, _25924_);
  nor _30368_ (_25926_, _25925_, _25714_);
  nor _30369_ (_25927_, _25926_, _25923_);
  nand _30370_ (_25928_, _25927_, _25623_);
  nand _30371_ (_25929_, _25841_, _25928_);
  nor _30372_ (_25930_, _25929_, _23940_);
  nor _30373_ (_25931_, _25930_, _25922_);
  not _30374_ (_25932_, _25638_);
  nor _30375_ (_25933_, _25709_, _25699_);
  nor _30376_ (_25934_, _25933_, _25696_);
  nor _30377_ (_25935_, _25934_, _23891_);
  nor _30378_ (_25936_, _25935_, _24004_);
  nor _30379_ (_25937_, _25936_, _25635_);
  nor _30380_ (_25938_, _25937_, _25932_);
  nor _30381_ (_25939_, _25938_, _25886_);
  not _30382_ (_25940_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _30383_ (_25941_, _25779_, _25940_);
  not _30384_ (_25942_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor _30385_ (_25943_, _25774_, _25942_);
  nor _30386_ (_25944_, _25943_, _25941_);
  not _30387_ (_25945_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _30388_ (_25946_, _25783_, _25945_);
  not _30389_ (_25947_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _30390_ (_25948_, _25790_, _25947_);
  nor _30391_ (_25949_, _25948_, _25946_);
  nand _30392_ (_25950_, _25949_, _25944_);
  not _30393_ (_25951_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _30394_ (_25952_, _25766_, _25951_);
  not _30395_ (_25953_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor _30396_ (_25954_, _25771_, _25953_);
  nor _30397_ (_25955_, _25954_, _25952_);
  not _30398_ (_25956_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor _30399_ (_25957_, _25787_, _25956_);
  not _30400_ (_25958_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _30401_ (_25959_, _25761_, _25958_);
  nor _30402_ (_25960_, _25959_, _25957_);
  nand _30403_ (_25961_, _25960_, _25955_);
  nor _30404_ (_25962_, _25961_, _25950_);
  nor _30405_ (_25963_, _25962_, _25758_);
  nor _30406_ (_25964_, _25879_, _25140_);
  nor _30407_ (_25965_, _25964_, _25963_);
  nor _30408_ (_25966_, _25965_, _25852_);
  nand _30409_ (_25967_, _25850_, _25719_);
  not _30410_ (_25968_, _25967_);
  nor _30411_ (_25969_, _24863_, _24005_);
  nor _30412_ (_25970_, _25243_, _24951_);
  not _30413_ (_25971_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _30414_ (_25972_, _24962_, _25971_);
  nor _30415_ (_25973_, _25972_, _25970_);
  not _30416_ (_25974_, _25973_);
  not _30417_ (_25975_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _30418_ (_25976_, _24949_, _25975_);
  nor _30419_ (_25977_, _24940_, _24959_);
  nor _30420_ (_25978_, _25977_, _25976_);
  nor _30421_ (_25979_, _24957_, _24935_);
  nor _30422_ (_25980_, _24953_, _24945_);
  nor _30423_ (_25981_, _25980_, _25979_);
  nand _30424_ (_25982_, _25981_, _25978_);
  nor _30425_ (_25983_, _25982_, _25974_);
  nor _30426_ (_25984_, _25983_, _25835_);
  nor _30427_ (_25985_, _25984_, _25969_);
  nor _30428_ (_25986_, _25985_, _25894_);
  nor _30429_ (_25987_, _25986_, _25968_);
  not _30430_ (_25988_, _25987_);
  nor _30431_ (_25989_, _25988_, _25966_);
  not _30432_ (_25990_, _25989_);
  nor _30433_ (_25991_, _25990_, _25939_);
  nor _30434_ (_25992_, _25991_, _24016_);
  not _30435_ (_25993_, _25991_);
  nor _30436_ (_25994_, _25993_, _24069_);
  nor _30437_ (_25995_, _25994_, _25992_);
  nor _30438_ (_25996_, _25995_, _25931_);
  nor _30439_ (_25997_, _24863_, _23971_);
  nor _30440_ (_25998_, _25243_, _25301_);
  nor _30441_ (_25999_, _24962_, _25304_);
  nor _30442_ (_26000_, _25999_, _25998_);
  not _30443_ (_26001_, _26000_);
  not _30444_ (_26002_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _30445_ (_26003_, _24949_, _26002_);
  nor _30446_ (_26004_, _24940_, _25314_);
  nor _30447_ (_26005_, _26004_, _26003_);
  nor _30448_ (_26006_, _24957_, _25311_);
  nor _30449_ (_26007_, _24953_, _25299_);
  nor _30450_ (_26008_, _26007_, _26006_);
  nand _30451_ (_26009_, _26008_, _26005_);
  nor _30452_ (_26010_, _26009_, _26001_);
  nor _30453_ (_26011_, _26010_, _25835_);
  nor _30454_ (_26012_, _26011_, _25997_);
  nor _30455_ (_26013_, _26012_, _25894_);
  nor _30456_ (_26014_, _25850_, _25526_);
  nand _30457_ (_26015_, _26014_, _25622_);
  nor _30458_ (_26016_, _26015_, _25734_);
  nor _30459_ (_26017_, _26016_, _26013_);
  not _30460_ (_26018_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _30461_ (_26019_, _25761_, _26018_);
  not _30462_ (_26020_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _30463_ (_26021_, _25771_, _26020_);
  nor _30464_ (_26023_, _26021_, _26019_);
  not _30465_ (_26024_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor _30466_ (_26025_, _25779_, _26024_);
  not _30467_ (_26026_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _30468_ (_26027_, _25783_, _26026_);
  nor _30469_ (_26028_, _26027_, _26025_);
  nand _30470_ (_26029_, _26028_, _26023_);
  not _30471_ (_26030_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _30472_ (_26031_, _25790_, _26030_);
  not _30473_ (_26032_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _30474_ (_26033_, _25774_, _26032_);
  nor _30475_ (_26034_, _26033_, _26031_);
  not _30476_ (_26035_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor _30477_ (_26036_, _25787_, _26035_);
  not _30478_ (_26037_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _30479_ (_26038_, _25766_, _26037_);
  nor _30480_ (_26039_, _26038_, _26036_);
  nand _30481_ (_26040_, _26039_, _26034_);
  nor _30482_ (_26041_, _26040_, _26029_);
  nor _30483_ (_26042_, _26041_, _25758_);
  nor _30484_ (_26043_, _25879_, _25029_);
  nor _30485_ (_26044_, _26043_, _26042_);
  nor _30486_ (_26045_, _26044_, _25852_);
  not _30487_ (_26046_, _25648_);
  nor _30488_ (_26047_, _25707_, _25700_);
  nor _30489_ (_26048_, _26047_, _25694_);
  nor _30490_ (_26049_, _26048_, _23891_);
  nor _30491_ (_26050_, _26049_, _23965_);
  nor _30492_ (_26051_, _26050_, _25635_);
  nor _30493_ (_26052_, _26051_, _26046_);
  nor _30494_ (_26053_, _26052_, _25886_);
  nor _30495_ (_26054_, _25818_, _25526_);
  nor _30496_ (_26055_, _26054_, _26053_);
  not _30497_ (_26056_, _26055_);
  nor _30498_ (_26057_, _26056_, _26045_);
  nand _30499_ (_26058_, _26057_, _26017_);
  not _30500_ (_26059_, _26058_);
  nor _30501_ (_26060_, _26059_, _23979_);
  nor _30502_ (_26061_, _26058_, _23978_);
  nor _30503_ (_26062_, _26061_, _26060_);
  nor _30504_ (_26063_, _25967_, _25819_);
  not _30505_ (_26064_, _25643_);
  nor _30506_ (_26065_, _25694_, _25645_);
  nor _30507_ (_26066_, _26065_, _25709_);
  nor _30508_ (_26067_, _26066_, _23891_);
  nor _30509_ (_26068_, _26067_, _24025_);
  nor _30510_ (_26069_, _26068_, _25635_);
  nor _30511_ (_26070_, _26069_, _26064_);
  nor _30512_ (_26071_, _26070_, _25886_);
  not _30513_ (_26072_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _30514_ (_26073_, _25761_, _26072_);
  not _30515_ (_26074_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _30516_ (_26075_, _25790_, _26074_);
  nor _30517_ (_26076_, _26075_, _26073_);
  not _30518_ (_26077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _30519_ (_26078_, _25766_, _26077_);
  not _30520_ (_26079_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _30521_ (_26080_, _25771_, _26079_);
  nor _30522_ (_26081_, _26080_, _26078_);
  nand _30523_ (_26082_, _26081_, _26076_);
  not _30524_ (_26083_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor _30525_ (_26084_, _25787_, _26083_);
  not _30526_ (_26085_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _30527_ (_26086_, _25774_, _26085_);
  nor _30528_ (_26087_, _26086_, _26084_);
  not _30529_ (_26088_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor _30530_ (_26089_, _25779_, _26088_);
  not _30531_ (_26090_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _30532_ (_26091_, _25783_, _26090_);
  nor _30533_ (_26092_, _26091_, _26089_);
  nand _30534_ (_26093_, _26092_, _26087_);
  nor _30535_ (_26094_, _26093_, _26082_);
  nor _30536_ (_26095_, _26094_, _25758_);
  not _30537_ (_26096_, _24920_);
  nor _30538_ (_26097_, _25879_, _26096_);
  nor _30539_ (_26098_, _26097_, _26095_);
  nor _30540_ (_26099_, _26098_, _25852_);
  nor _30541_ (_26100_, _24863_, _24026_);
  nor _30542_ (_26101_, _25243_, _25370_);
  not _30543_ (_26102_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _30544_ (_26103_, _24962_, _26102_);
  nor _30545_ (_26104_, _26103_, _26101_);
  not _30546_ (_26105_, _26104_);
  not _30547_ (_26106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _30548_ (_26107_, _24949_, _26106_);
  nor _30549_ (_26108_, _24957_, _25364_);
  nor _30550_ (_26109_, _26108_, _26107_);
  not _30551_ (_26110_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _30552_ (_26111_, _24953_, _26110_);
  nor _30553_ (_26112_, _24940_, _25362_);
  nor _30554_ (_26113_, _26112_, _26111_);
  nand _30555_ (_26114_, _26113_, _26109_);
  nor _30556_ (_26115_, _26114_, _26105_);
  nor _30557_ (_26117_, _26115_, _25835_);
  nor _30558_ (_26118_, _26117_, _26100_);
  nor _30559_ (_26119_, _26118_, _25894_);
  nor _30560_ (_26120_, _26119_, _26099_);
  not _30561_ (_26121_, _26120_);
  nor _30562_ (_26122_, _26121_, _26071_);
  not _30563_ (_26123_, _26122_);
  nor _30564_ (_26124_, _26123_, _26063_);
  nor _30565_ (_26125_, _26124_, _24035_);
  not _30566_ (_26126_, _26124_);
  nor _30567_ (_26127_, _26126_, _24060_);
  nor _30568_ (_26129_, _26127_, _26125_);
  nor _30569_ (_26130_, _26129_, _26062_);
  nand _30570_ (_26131_, _26130_, _25996_);
  nor _30571_ (_26132_, _26131_, _25921_);
  nor _30572_ (_26133_, _24051_, _23996_);
  not _30573_ (_26134_, _26133_);
  nor _30574_ (_26135_, _26134_, _23958_);
  nor _30575_ (_26136_, _26135_, _25631_);
  nand _30576_ (_26137_, _26136_, _26132_);
  nor _30577_ (_26138_, _26137_, _25849_);
  nor _30578_ (_26139_, _25549_, _25461_);
  nor _30579_ (_26140_, _25509_, _25423_);
  nor _30580_ (_26141_, _26140_, _26139_);
  nor _30581_ (_26142_, _26141_, _25530_);
  nor _30582_ (_26143_, _25849_, _24684_);
  nor _30583_ (_26144_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _30584_ (_26145_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _30585_ (_26146_, _26145_, _26144_);
  nor _30586_ (_26147_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _30587_ (_26148_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand _30588_ (_26149_, _26148_, _26147_);
  nor _30589_ (_26150_, _26149_, _26146_);
  nand _30590_ (_26151_, _26150_, _25508_);
  not _30591_ (_26152_, _24645_);
  nor _30592_ (_26153_, _26152_, _24578_);
  nor _30593_ (_26154_, _24645_, _24579_);
  nor _30594_ (_26155_, _26154_, _26153_);
  nand _30595_ (_26156_, _24643_, _24604_);
  not _30596_ (_26157_, _26156_);
  nor _30597_ (_26158_, _26157_, _24644_);
  nand _30598_ (_26159_, _24641_, _24607_);
  nand _30599_ (_26160_, _26159_, _24643_);
  not _30600_ (_26161_, _24639_);
  nor _30601_ (_26162_, _26161_, _24249_);
  nor _30602_ (_26163_, _24639_, _24250_);
  nor _30603_ (_26164_, _26163_, _26162_);
  not _30604_ (_26165_, _26164_);
  nand _30605_ (_26166_, _24633_, _24621_);
  not _30606_ (_26167_, _26166_);
  nor _30607_ (_26168_, _26167_, _24634_);
  not _30608_ (_26169_, _25618_);
  nor _30609_ (_26170_, _24510_, _24497_);
  nor _30610_ (_26171_, _26170_, _24512_);
  not _30611_ (_26172_, _26171_);
  nor _30612_ (_26173_, _24627_, _24624_);
  nand _30613_ (_26174_, _26173_, _26172_);
  nor _30614_ (_26175_, _26174_, _26169_);
  nand _30615_ (_26176_, _26175_, _26168_);
  nor _30616_ (_26177_, _26176_, _25846_);
  nand _30617_ (_26178_, _26177_, _26165_);
  nor _30618_ (_26179_, _26178_, _26160_);
  nand _30619_ (_26180_, _26179_, _26158_);
  nor _30620_ (_26182_, _26180_, _26155_);
  nand _30621_ (_26183_, _25846_, _25809_);
  nor _30622_ (_26184_, _26183_, _24490_);
  nor _30623_ (_26185_, _26184_, _26182_);
  nand _30624_ (_26186_, _26185_, _26151_);
  nor _30625_ (_26187_, _26186_, _26143_);
  nor _30626_ (_26188_, _25808_, _25327_);
  nor _30627_ (_26189_, _26188_, _25542_);
  nor _30628_ (_26190_, _26189_, _26187_);
  nor _30629_ (_26191_, _25393_, _25474_);
  nor _30630_ (_26192_, _26191_, _25482_);
  nor _30631_ (_26193_, _25563_, _25412_);
  nor _30632_ (_26194_, _25329_, _25235_);
  not _30633_ (_26195_, _26194_);
  nor _30634_ (_26196_, _26195_, _25563_);
  nor _30635_ (_26197_, _26196_, _26193_);
  not _30636_ (_26198_, _26197_);
  nor _30637_ (_26199_, _26198_, _26192_);
  not _30638_ (_26200_, _25574_);
  nor _30639_ (_26201_, _25548_, _25267_);
  not _30640_ (_26202_, _26201_);
  nor _30641_ (_26203_, _26202_, _25426_);
  not _30642_ (_26204_, _26203_);
  nand _30643_ (_26205_, _26204_, _26200_);
  nor _30644_ (_26206_, _26195_, _25420_);
  nor _30645_ (_26207_, _26206_, _26205_);
  not _30646_ (_26208_, _26207_);
  nor _30647_ (_26209_, _26208_, _25537_);
  nand _30648_ (_26210_, _26209_, _26199_);
  nand _30649_ (_26211_, _26210_, _26187_);
  nor _30650_ (_26212_, _25493_, _25482_);
  nor _30651_ (_26213_, _26212_, _25476_);
  not _30652_ (_26214_, _26213_);
  nor _30653_ (_26215_, _26214_, _25487_);
  nand _30654_ (_26216_, _26215_, _26211_);
  nor _30655_ (_26217_, _26216_, _26190_);
  nor _30656_ (_26218_, _25613_, _25504_);
  nor _30657_ (_26220_, _26218_, _26217_);
  nor _30658_ (_26221_, _26220_, _26142_);
  not _30659_ (_26222_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not _30660_ (_26223_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  nor _30661_ (_26224_, _26223_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _30662_ (_26225_, _26224_, _26222_);
  not _30663_ (_26226_, _26225_);
  nor _30664_ (_26227_, _26222_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _30665_ (_26228_, _26227_);
  nor _30666_ (_26229_, _26228_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  nor _30667_ (_26230_, _24035_, _23978_);
  not _30668_ (_26231_, _26230_);
  nor _30669_ (_26232_, _26231_, _25728_);
  nor _30670_ (_26233_, _26232_, _26229_);
  not _30671_ (_26234_, _26233_);
  nor _30672_ (_26235_, _26234_, _26226_);
  not _30673_ (_26236_, _26235_);
  nor _30674_ (_26237_, _25724_, _23915_);
  not _30675_ (_26238_, _26237_);
  nor _30676_ (_26239_, _26238_, _23978_);
  nor _30677_ (_26240_, _24035_, _24016_);
  not _30678_ (_26241_, _26240_);
  nor _30679_ (_26242_, _23875_, _23871_);
  not _30680_ (_26243_, _26242_);
  nor _30681_ (_26244_, _26243_, _23939_);
  not _30682_ (_26245_, _26244_);
  nor _30683_ (_26246_, _26245_, _26241_);
  nand _30684_ (_26247_, _26246_, _26239_);
  not _30685_ (_26248_, _26247_);
  nor _30686_ (_26249_, _26248_, _26236_);
  not _30687_ (_26250_, _26249_);
  nand _30688_ (_26251_, _26250_, _25508_);
  nor _30689_ (_26252_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _30690_ (_26253_, _26252_);
  nor _30691_ (_26254_, _26253_, _25729_);
  nor _30692_ (_26255_, _26238_, _23979_);
  not _30693_ (_26256_, _26255_);
  nor _30694_ (_26257_, _24060_, _24016_);
  not _30695_ (_26258_, _26257_);
  nor _30696_ (_26259_, _26258_, _26245_);
  not _30697_ (_26260_, _26259_);
  nor _30698_ (_26261_, _26260_, _26256_);
  not _30699_ (_26262_, _26261_);
  nand _30700_ (_26263_, _26262_, _26254_);
  nand _30701_ (_26264_, _26263_, _25617_);
  nand _30702_ (_26265_, _26264_, _26251_);
  nor _30703_ (_26266_, _26265_, _26221_);
  not _30704_ (_26267_, _26132_);
  not _30705_ (_26268_, _25688_);
  nor _30706_ (_26269_, _26268_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  not _30707_ (_26270_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _30708_ (_26271_, _25688_, _26270_);
  nor _30709_ (_26272_, _26271_, _26269_);
  nand _30710_ (_26273_, _26272_, _23952_);
  not _30711_ (_26274_, _26273_);
  nor _30712_ (_26275_, _26274_, _23953_);
  nor _30713_ (_26276_, _26275_, _25635_);
  nor _30714_ (_26277_, _26276_, _25687_);
  nor _30715_ (_26278_, _26277_, _25886_);
  not _30716_ (_26279_, _26278_);
  nor _30717_ (_26281_, _26015_, _25459_);
  not _30718_ (_26282_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _30719_ (_26283_, _25761_, _26282_);
  not _30720_ (_26284_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _30721_ (_26285_, _25766_, _26284_);
  nor _30722_ (_26286_, _26285_, _26283_);
  not _30723_ (_26287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _30724_ (_26288_, _25771_, _26287_);
  not _30725_ (_26289_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor _30726_ (_26290_, _25779_, _26289_);
  nor _30727_ (_26291_, _26290_, _26288_);
  nand _30728_ (_26292_, _26291_, _26286_);
  not _30729_ (_26293_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor _30730_ (_26294_, _25774_, _26293_);
  not _30731_ (_26295_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _30732_ (_26296_, _25783_, _26295_);
  nor _30733_ (_26298_, _26296_, _26294_);
  not _30734_ (_26299_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor _30735_ (_26300_, _25787_, _26299_);
  not _30736_ (_26301_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _30737_ (_26302_, _25790_, _26301_);
  nor _30738_ (_26303_, _26302_, _26300_);
  nand _30739_ (_26304_, _26303_, _26298_);
  nor _30740_ (_26305_, _26304_, _26292_);
  nor _30741_ (_26306_, _26305_, _25758_);
  nor _30742_ (_26307_, _25879_, _24820_);
  nor _30743_ (_26309_, _26307_, _26306_);
  not _30744_ (_26310_, _26309_);
  nand _30745_ (_26311_, _26310_, _25851_);
  nor _30746_ (_26312_, _24863_, _23945_);
  nor _30747_ (_26313_, _25243_, _25440_);
  not _30748_ (_26314_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _30749_ (_26315_, _24962_, _26314_);
  nor _30750_ (_26317_, _26315_, _26313_);
  not _30751_ (_26318_, _26317_);
  not _30752_ (_26319_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _30753_ (_26320_, _24949_, _26319_);
  nor _30754_ (_26322_, _24940_, _25432_);
  nor _30755_ (_26323_, _26322_, _26320_);
  nor _30756_ (_26324_, _24957_, _25434_);
  not _30757_ (_26325_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _30758_ (_26326_, _24953_, _26325_);
  nor _30759_ (_26328_, _26326_, _26324_);
  nand _30760_ (_26329_, _26328_, _26323_);
  nor _30761_ (_26330_, _26329_, _26318_);
  nor _30762_ (_26331_, _26330_, _25835_);
  nor _30763_ (_26332_, _26331_, _26312_);
  nor _30764_ (_26333_, _26332_, _25894_);
  not _30765_ (_26334_, _26333_);
  nand _30766_ (_26335_, _26334_, _26311_);
  nor _30767_ (_26337_, _26335_, _26281_);
  nand _30768_ (_26338_, _26337_, _26279_);
  nor _30769_ (_26339_, _26338_, _23958_);
  not _30770_ (_26340_, _26339_);
  not _30771_ (_26341_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _30772_ (_26342_, _25779_, _26341_);
  not _30773_ (_26343_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _30774_ (_26344_, _25774_, _26343_);
  nor _30775_ (_26345_, _26344_, _26342_);
  not _30776_ (_26346_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _30777_ (_26347_, _25783_, _26346_);
  not _30778_ (_26348_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _30779_ (_26349_, _25790_, _26348_);
  nor _30780_ (_26350_, _26349_, _26347_);
  nand _30781_ (_26351_, _26350_, _26345_);
  not _30782_ (_26352_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _30783_ (_26353_, _25766_, _26352_);
  not _30784_ (_26354_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _30785_ (_26355_, _25771_, _26354_);
  nor _30786_ (_26356_, _26355_, _26353_);
  not _30787_ (_26357_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor _30788_ (_26358_, _25787_, _26357_);
  not _30789_ (_26359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _30790_ (_26360_, _25761_, _26359_);
  nor _30791_ (_26361_, _26360_, _26358_);
  nand _30792_ (_26362_, _26361_, _26356_);
  nor _30793_ (_26363_, _26362_, _26351_);
  nor _30794_ (_26364_, _26363_, _25758_);
  nor _30795_ (_26365_, _25879_, _25703_);
  nor _30796_ (_26366_, _26365_, _26364_);
  nor _30797_ (_26367_, _26366_, _25852_);
  nor _30798_ (_26368_, _24863_, _24042_);
  nor _30799_ (_26369_, _25243_, _25277_);
  not _30800_ (_26370_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _30801_ (_26371_, _24962_, _26370_);
  nor _30802_ (_26372_, _26371_, _26369_);
  not _30803_ (_26373_, _26372_);
  not _30804_ (_26374_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _30805_ (_26375_, _24949_, _26374_);
  nor _30806_ (_26376_, _24940_, _25271_);
  nor _30807_ (_26377_, _26376_, _26375_);
  nor _30808_ (_26378_, _24957_, _25282_);
  not _30809_ (_26379_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _30810_ (_26380_, _24953_, _26379_);
  nor _30811_ (_26381_, _26380_, _26378_);
  nand _30812_ (_26382_, _26381_, _26377_);
  nor _30813_ (_26383_, _26382_, _26373_);
  nor _30814_ (_26384_, _26383_, _25835_);
  nor _30815_ (_26385_, _26384_, _26368_);
  nor _30816_ (_26386_, _26385_, _25894_);
  nor _30817_ (_26387_, _26386_, _26367_);
  not _30818_ (_26388_, _24039_);
  not _30819_ (_26389_, _25685_);
  nor _30820_ (_26390_, _25689_, _26389_);
  nor _30821_ (_26391_, _26390_, _25705_);
  nor _30822_ (_26392_, _26391_, _25692_);
  nor _30823_ (_26393_, _26392_, _23891_);
  nor _30824_ (_26394_, _26393_, _26388_);
  nor _30825_ (_26395_, _26394_, _25635_);
  nor _30826_ (_26396_, _26395_, _25704_);
  nor _30827_ (_26397_, _26396_, _25886_);
  nor _30828_ (_26398_, _26015_, _25460_);
  nor _30829_ (_26399_, _26398_, _26397_);
  nand _30830_ (_26400_, _26399_, _26387_);
  nor _30831_ (_26401_, _26400_, _24051_);
  not _30832_ (_26402_, _24051_);
  not _30833_ (_26403_, _26400_);
  nor _30834_ (_26404_, _26403_, _26402_);
  nor _30835_ (_26405_, _26404_, _26401_);
  nand _30836_ (_26406_, _26405_, _26340_);
  not _30837_ (_26407_, _26338_);
  nor _30838_ (_26408_, _26407_, _25721_);
  not _30839_ (_26409_, _26408_);
  not _30840_ (_26410_, _23996_);
  nor _30841_ (_26411_, _24863_, _23987_);
  nor _30842_ (_26412_, _25243_, _25240_);
  nor _30843_ (_26413_, _24962_, _25242_);
  nor _30844_ (_26414_, _26413_, _26412_);
  not _30845_ (_26415_, _26414_);
  not _30846_ (_26416_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor _30847_ (_26417_, _24949_, _26416_);
  nor _30848_ (_26418_, _24940_, _25253_);
  nor _30849_ (_26419_, _26418_, _26417_);
  nor _30850_ (_26420_, _24957_, _25250_);
  nor _30851_ (_26421_, _24953_, _25237_);
  nor _30852_ (_26422_, _26421_, _26420_);
  nand _30853_ (_26423_, _26422_, _26419_);
  nor _30854_ (_26424_, _26423_, _26415_);
  nor _30855_ (_26425_, _26424_, _25835_);
  nor _30856_ (_26426_, _26425_, _26411_);
  nor _30857_ (_26427_, _26426_, _25894_);
  not _30858_ (_26428_, _26427_);
  nor _30859_ (_26429_, _25818_, _25719_);
  nor _30860_ (_26430_, _26015_, _25266_);
  nor _30861_ (_26431_, _26430_, _26429_);
  nand _30862_ (_26432_, _26431_, _26428_);
  not _30863_ (_26433_, _26432_);
  not _30864_ (_26434_, _23984_);
  nor _30865_ (_26435_, _25690_, _25685_);
  nor _30866_ (_26436_, _26435_, _26390_);
  nor _30867_ (_26437_, _26436_, _23891_);
  nor _30868_ (_26438_, _26437_, _26434_);
  nor _30869_ (_26439_, _26438_, _25635_);
  nor _30870_ (_26440_, _26439_, _25684_);
  nor _30871_ (_26441_, _26440_, _25886_);
  not _30872_ (_26442_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _30873_ (_26443_, _25761_, _26442_);
  not _30874_ (_26444_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _30875_ (_26445_, _25766_, _26444_);
  nor _30876_ (_26447_, _26445_, _26443_);
  not _30877_ (_26448_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _30878_ (_26449_, _25771_, _26448_);
  not _30879_ (_26450_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _30880_ (_26451_, _25774_, _26450_);
  nor _30881_ (_26452_, _26451_, _26449_);
  nand _30882_ (_26453_, _26452_, _26447_);
  not _30883_ (_26454_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _30884_ (_26455_, _25779_, _26454_);
  not _30885_ (_26456_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _30886_ (_26457_, _25783_, _26456_);
  nor _30887_ (_26458_, _26457_, _26455_);
  not _30888_ (_26459_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _30889_ (_26460_, _25787_, _26459_);
  not _30890_ (_26461_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor _30891_ (_26463_, _25790_, _26461_);
  nor _30892_ (_26464_, _26463_, _26460_);
  nand _30893_ (_26465_, _26464_, _26458_);
  nor _30894_ (_26466_, _26465_, _26453_);
  nor _30895_ (_26467_, _26466_, _25758_);
  nor _30896_ (_26468_, _25879_, _25088_);
  nor _30897_ (_26469_, _26468_, _26467_);
  nor _30898_ (_26470_, _26469_, _25852_);
  nor _30899_ (_26471_, _26470_, _26441_);
  nand _30900_ (_26472_, _26471_, _26433_);
  not _30901_ (_26473_, _26472_);
  nor _30902_ (_26474_, _26473_, _26410_);
  nor _30903_ (_26475_, _26472_, _23996_);
  nor _30904_ (_26476_, _26475_, _26474_);
  nand _30905_ (_26477_, _26476_, _26409_);
  nor _30906_ (_26478_, _26477_, _26406_);
  nand _30907_ (_26480_, _26478_, _26242_);
  nor _30908_ (_26481_, _26480_, _26267_);
  nor _30909_ (_26482_, _23915_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand _30910_ (_26483_, _26482_, _26481_);
  nand _30911_ (_26484_, _26483_, _26266_);
  nor _30912_ (_26485_, _26484_, _26138_);
  not _30913_ (_26486_, _26485_);
  not _30914_ (_26487_, rst);
  nand _30915_ (_26488_, _25614_, _26487_);
  nor _30916_ (_28209_, _26488_, _26486_);
  not _30917_ (_26489_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r );
  nor _30918_ (_28210_, _26489_, rst);
  nor _30919_ (_26490_, _25426_, _25235_);
  nor _30920_ (_26491_, _26490_, _25427_);
  nand _30921_ (_26492_, _26491_, _25544_);
  nor _30922_ (_26493_, _26492_, _26205_);
  nor _30923_ (_26494_, _26493_, _25505_);
  nand _30924_ (_26495_, _26140_, _25499_);
  nor _30925_ (_26496_, _25530_, _25482_);
  nand _30926_ (_26498_, _26496_, _25396_);
  not _30927_ (_26499_, _26498_);
  nor _30928_ (_26500_, _26499_, _25613_);
  nand _30929_ (_26501_, _26500_, _26495_);
  nor _30930_ (_26502_, _26501_, _26494_);
  nor _30931_ (_26503_, _24863_, _23908_);
  not _30932_ (_26504_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  nor _30933_ (_26505_, _26504_, _25207_);
  nor _30934_ (_26506_, _24953_, _25825_);
  nor _30935_ (_26507_, _24957_, _25332_);
  nor _30936_ (_26508_, _26507_, _26506_);
  not _30937_ (_26509_, _26508_);
  not _30938_ (_26510_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor _30939_ (_26511_, _24949_, _26510_);
  nor _30940_ (_26512_, _24962_, _25338_);
  nor _30941_ (_26513_, _26512_, _26511_);
  nor _30942_ (_26514_, _24940_, _25343_);
  nor _30943_ (_26515_, _25243_, _25336_);
  nor _30944_ (_26517_, _26515_, _26514_);
  nand _30945_ (_26518_, _26517_, _26513_);
  nor _30946_ (_26519_, _26518_, _26509_);
  nor _30947_ (_26520_, _26519_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _30948_ (_26521_, _26520_, _26505_);
  nor _30949_ (_26522_, _26521_, _24864_);
  nor _30950_ (_26523_, _26522_, _26503_);
  not _30951_ (_26524_, _26523_);
  nor _30952_ (_26525_, _26524_, _26502_);
  not _30953_ (_26526_, _26502_);
  nor _30954_ (_26527_, _26526_, _25838_);
  nor _30955_ (_26528_, _26527_, _26525_);
  not _30956_ (_26529_, _26528_);
  nor _30957_ (_26530_, _26529_, _24090_);
  not _30958_ (_26531_, _26530_);
  nor _30959_ (_26532_, _26528_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _30960_ (_26533_, _26532_);
  nor _30961_ (_26534_, _24863_, _24012_);
  not _30962_ (_26535_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  nor _30963_ (_26536_, _26535_, _25207_);
  not _30964_ (_26537_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor _30965_ (_26538_, _24949_, _26537_);
  nor _30966_ (_26539_, _24940_, _25971_);
  nor _30967_ (_26540_, _26539_, _26538_);
  not _30968_ (_26541_, _26540_);
  nor _30969_ (_26542_, _25243_, _24945_);
  nor _30970_ (_26543_, _24957_, _24959_);
  nor _30971_ (_26544_, _26543_, _26542_);
  nor _30972_ (_26545_, _24953_, _25975_);
  nor _30973_ (_26546_, _24962_, _24951_);
  nor _30974_ (_26547_, _26546_, _26545_);
  nand _30975_ (_26548_, _26547_, _26544_);
  nor _30976_ (_26549_, _26548_, _26541_);
  nor _30977_ (_26550_, _26549_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _30978_ (_26551_, _26550_, _26536_);
  nor _30979_ (_26552_, _26551_, _24864_);
  nor _30980_ (_26553_, _26552_, _26534_);
  nand _30981_ (_26554_, _26553_, _26526_);
  nand _30982_ (_26555_, _26502_, _25985_);
  nand _30983_ (_26556_, _26555_, _26554_);
  nor _30984_ (_26557_, _26556_, _24527_);
  not _30985_ (_26558_, _26557_);
  nand _30986_ (_26559_, _26556_, _24527_);
  nand _30987_ (_26560_, _26559_, _26558_);
  not _30988_ (_26561_, _26560_);
  nor _30989_ (_26562_, _24863_, _24031_);
  not _30990_ (_26563_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  nor _30991_ (_26564_, _26563_, _25207_);
  nor _30992_ (_26565_, _25243_, _26110_);
  nor _30993_ (_26566_, _24940_, _26102_);
  nor _30994_ (_26567_, _26566_, _26565_);
  nor _30995_ (_26568_, _24953_, _26106_);
  nor _30996_ (_26569_, _24962_, _25370_);
  nor _30997_ (_26570_, _26569_, _26568_);
  nand _30998_ (_26571_, _26570_, _26567_);
  not _30999_ (_26572_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _31000_ (_26573_, _24949_, _26572_);
  nor _31001_ (_26574_, _24957_, _25362_);
  nor _31002_ (_26575_, _26574_, _26573_);
  not _31003_ (_26576_, _26575_);
  nor _31004_ (_26577_, _26576_, _26571_);
  nor _31005_ (_26578_, _26577_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _31006_ (_26579_, _26578_, _26564_);
  nor _31007_ (_26580_, _26579_, _24864_);
  nor _31008_ (_26581_, _26580_, _26562_);
  nand _31009_ (_26582_, _26581_, _26526_);
  nand _31010_ (_26583_, _26502_, _26118_);
  nand _31011_ (_26584_, _26583_, _26582_);
  nor _31012_ (_26585_, _26584_, _24153_);
  not _31013_ (_26586_, _26585_);
  nand _31014_ (_26587_, _26584_, _24153_);
  nor _31015_ (_26588_, _24863_, _23966_);
  not _31016_ (_26589_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  nor _31017_ (_26590_, _26589_, _25207_);
  not _31018_ (_26591_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _31019_ (_26592_, _24949_, _26591_);
  nor _31020_ (_26593_, _24940_, _25304_);
  nor _31021_ (_26594_, _26593_, _26592_);
  not _31022_ (_26595_, _26594_);
  nor _31023_ (_26596_, _25243_, _25299_);
  nor _31024_ (_26597_, _24957_, _25314_);
  nor _31025_ (_26598_, _26597_, _26596_);
  nor _31026_ (_26599_, _24953_, _26002_);
  nor _31027_ (_26600_, _24962_, _25301_);
  nor _31028_ (_26601_, _26600_, _26599_);
  nand _31029_ (_26602_, _26601_, _26598_);
  nor _31030_ (_26603_, _26602_, _26595_);
  nor _31031_ (_26604_, _26603_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _31032_ (_26605_, _26604_, _26590_);
  nor _31033_ (_26606_, _26605_, _24864_);
  nor _31034_ (_26607_, _26606_, _26588_);
  not _31035_ (_26608_, _26607_);
  nor _31036_ (_26609_, _26608_, _26502_);
  not _31037_ (_26610_, _26012_);
  nor _31038_ (_26611_, _26526_, _26610_);
  nor _31039_ (_26612_, _26611_, _26609_);
  not _31040_ (_26613_, _26612_);
  nor _31041_ (_26614_, _26613_, _24202_);
  not _31042_ (_26615_, _26614_);
  nor _31043_ (_26616_, _24863_, _23932_);
  not _31044_ (_26618_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  nor _31045_ (_26619_, _26618_, _25207_);
  not _31046_ (_26620_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor _31047_ (_26621_, _24949_, _26620_);
  nor _31048_ (_26622_, _24940_, _25897_);
  nor _31049_ (_26623_, _26622_, _26621_);
  not _31050_ (_26624_, _26623_);
  nor _31051_ (_26625_, _25243_, _25208_);
  nor _31052_ (_26626_, _24957_, _25903_);
  nor _31053_ (_26627_, _26626_, _26625_);
  nor _31054_ (_26628_, _24953_, _25901_);
  nor _31055_ (_26629_, _24962_, _25220_);
  nor _31056_ (_26630_, _26629_, _26628_);
  nand _31057_ (_26632_, _26630_, _26627_);
  nor _31058_ (_26633_, _26632_, _26624_);
  nor _31059_ (_26634_, _26633_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _31060_ (_26635_, _26634_, _26619_);
  nor _31061_ (_26636_, _26635_, _24864_);
  nor _31062_ (_26637_, _26636_, _26616_);
  not _31063_ (_26638_, _26637_);
  nor _31064_ (_26639_, _26638_, _26502_);
  not _31065_ (_26640_, _25912_);
  nor _31066_ (_26641_, _26526_, _26640_);
  nor _31067_ (_26642_, _26641_, _26639_);
  not _31068_ (_26643_, _26642_);
  nor _31069_ (_26644_, _26643_, _24251_);
  not _31070_ (_26645_, _26644_);
  nor _31071_ (_26646_, _26642_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _31072_ (_26647_, _26646_);
  nor _31073_ (_26648_, _24863_, _24045_);
  not _31074_ (_26649_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  nor _31075_ (_26650_, _26649_, _25207_);
  nor _31076_ (_26651_, _25243_, _26379_);
  nor _31077_ (_26652_, _24940_, _26370_);
  nor _31078_ (_26653_, _26652_, _26651_);
  nor _31079_ (_26654_, _24953_, _26374_);
  nor _31080_ (_26655_, _24962_, _25277_);
  nor _31081_ (_26656_, _26655_, _26654_);
  nand _31082_ (_26657_, _26656_, _26653_);
  not _31083_ (_26658_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor _31084_ (_26659_, _24949_, _26658_);
  nor _31085_ (_26660_, _24957_, _25271_);
  nor _31086_ (_26661_, _26660_, _26659_);
  not _31087_ (_26662_, _26661_);
  nor _31088_ (_26663_, _26662_, _26657_);
  nor _31089_ (_26664_, _26663_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _31090_ (_26665_, _26664_, _26650_);
  nor _31091_ (_26666_, _26665_, _24864_);
  nor _31092_ (_26667_, _26666_, _26648_);
  not _31093_ (_26668_, _26667_);
  nor _31094_ (_26669_, _26668_, _26502_);
  nand _31095_ (_26670_, _26502_, _26385_);
  not _31096_ (_26671_, _26670_);
  nor _31097_ (_26672_, _26671_, _26669_);
  not _31098_ (_26673_, _26672_);
  nor _31099_ (_26674_, _26673_, _24305_);
  not _31100_ (_26675_, _26674_);
  nor _31101_ (_26676_, _24863_, _23990_);
  not _31102_ (_26677_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  nor _31103_ (_26678_, _26677_, _25207_);
  not _31104_ (_26679_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor _31105_ (_26680_, _24949_, _26679_);
  nor _31106_ (_26681_, _24940_, _25242_);
  nor _31107_ (_26682_, _26681_, _26680_);
  not _31108_ (_26683_, _26682_);
  nor _31109_ (_26684_, _25243_, _25237_);
  nor _31110_ (_26685_, _24957_, _25253_);
  nor _31111_ (_26686_, _26685_, _26684_);
  nor _31112_ (_26687_, _24953_, _26416_);
  nor _31113_ (_26688_, _24962_, _25240_);
  nor _31114_ (_26689_, _26688_, _26687_);
  nand _31115_ (_26690_, _26689_, _26686_);
  nor _31116_ (_26691_, _26690_, _26683_);
  nor _31117_ (_26692_, _26691_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _31118_ (_26693_, _26692_, _26678_);
  nor _31119_ (_26694_, _26693_, _24864_);
  nor _31120_ (_26695_, _26694_, _26676_);
  not _31121_ (_26696_, _26695_);
  nor _31122_ (_26697_, _26696_, _26502_);
  nand _31123_ (_26698_, _26502_, _26426_);
  not _31124_ (_26699_, _26698_);
  nor _31125_ (_26700_, _26699_, _26697_);
  nand _31126_ (_26701_, _26700_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _31127_ (_26702_, _24863_, _24406_);
  not _31128_ (_26703_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  nor _31129_ (_26704_, _26703_, _25207_);
  not _31130_ (_26705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor _31131_ (_26706_, _24949_, _26705_);
  nor _31132_ (_26707_, _24940_, _26314_);
  nor _31133_ (_26708_, _26707_, _26706_);
  not _31134_ (_26709_, _26708_);
  nor _31135_ (_26710_, _25243_, _26325_);
  nor _31136_ (_26711_, _24957_, _25432_);
  nor _31137_ (_26712_, _26711_, _26710_);
  nor _31138_ (_26713_, _24953_, _26319_);
  nor _31139_ (_26714_, _24962_, _25440_);
  nor _31140_ (_26715_, _26714_, _26713_);
  nand _31141_ (_26716_, _26715_, _26712_);
  nor _31142_ (_26717_, _26716_, _26709_);
  nor _31143_ (_26718_, _26717_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _31144_ (_26719_, _26718_, _26704_);
  nor _31145_ (_26720_, _26719_, _24864_);
  nor _31146_ (_26721_, _26720_, _26702_);
  not _31147_ (_26722_, _26721_);
  nor _31148_ (_26723_, _26722_, _26502_);
  not _31149_ (_26724_, _26332_);
  nor _31150_ (_26725_, _26526_, _26724_);
  nor _31151_ (_26726_, _26725_, _26723_);
  nand _31152_ (_26727_, _26726_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _31153_ (_26728_, _26727_);
  not _31154_ (_26729_, _26697_);
  nand _31155_ (_26730_, _26698_, _26729_);
  nor _31156_ (_26731_, _26730_, _24364_);
  nor _31157_ (_26732_, _26700_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _31158_ (_26733_, _26732_, _26731_);
  nand _31159_ (_26734_, _26733_, _26728_);
  nand _31160_ (_26735_, _26734_, _26701_);
  nor _31161_ (_26736_, _26672_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _31162_ (_26737_, _26736_, _26674_);
  nand _31163_ (_26738_, _26737_, _26735_);
  nand _31164_ (_26739_, _26738_, _26675_);
  nand _31165_ (_26740_, _26739_, _26647_);
  nand _31166_ (_26741_, _26740_, _26645_);
  nor _31167_ (_26742_, _26612_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _31168_ (_26743_, _26742_, _26614_);
  nand _31169_ (_26744_, _26743_, _26741_);
  nand _31170_ (_26745_, _26744_, _26615_);
  nand _31171_ (_26746_, _26745_, _26587_);
  nand _31172_ (_26747_, _26746_, _26586_);
  nand _31173_ (_26748_, _26747_, _26561_);
  nand _31174_ (_26749_, _26748_, _26558_);
  nand _31175_ (_26750_, _26749_, _26533_);
  nand _31176_ (_26751_, _26750_, _26531_);
  nand _31177_ (_26752_, _26751_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _31178_ (_26753_, _26752_, _24374_);
  nand _31179_ (_26754_, _26753_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _31180_ (_26755_, _26754_, _24253_);
  nand _31181_ (_26756_, _26755_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _31182_ (_26757_, _26756_, _24151_);
  nor _31183_ (_26758_, _26757_, _26528_);
  nand _31184_ (_26759_, _26730_, _24364_);
  nand _31185_ (_26760_, _26759_, _26701_);
  nor _31186_ (_26761_, _26760_, _26727_);
  nor _31187_ (_26762_, _26761_, _26731_);
  not _31188_ (_26763_, _26737_);
  nor _31189_ (_26764_, _26763_, _26762_);
  nor _31190_ (_26765_, _26764_, _26674_);
  nor _31191_ (_26766_, _26765_, _26646_);
  nor _31192_ (_26767_, _26766_, _26644_);
  not _31193_ (_26768_, _26743_);
  nor _31194_ (_26769_, _26768_, _26767_);
  nor _31195_ (_26770_, _26769_, _26614_);
  nand _31196_ (_26771_, _26770_, _26586_);
  nand _31197_ (_26772_, _26771_, _26587_);
  nor _31198_ (_26773_, _26772_, _26560_);
  nor _31199_ (_26774_, _26773_, _26557_);
  nor _31200_ (_26775_, _26774_, _26532_);
  nor _31201_ (_26776_, _26775_, _26530_);
  nand _31202_ (_26777_, _26776_, _24398_);
  nor _31203_ (_26778_, _26777_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _31204_ (_26779_, _26778_, _24308_);
  nor _31205_ (_26780_, _26779_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _31206_ (_26781_, _26780_, _24204_);
  nor _31207_ (_26782_, _26781_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _31208_ (_26783_, _26782_, _26529_);
  nor _31209_ (_26784_, _26783_, _26758_);
  nor _31210_ (_26785_, _26528_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _31211_ (_26786_, _26529_, _24529_);
  nor _31212_ (_26787_, _26786_, _26785_);
  nand _31213_ (_26788_, _26787_, _26784_);
  nand _31214_ (_26789_, _26788_, _24095_);
  not _31215_ (_26790_, _25808_);
  nor _31216_ (_26791_, _26214_, _26790_);
  nand _31217_ (_26792_, _26791_, _26207_);
  nor _31218_ (_26793_, _26792_, _26492_);
  nor _31219_ (_26794_, _26793_, _25505_);
  nor _31220_ (_26795_, _26794_, _26499_);
  not _31221_ (_26796_, _25476_);
  nor _31222_ (_26797_, _26796_, _25505_);
  nor _31223_ (_26798_, _26797_, _26142_);
  nor _31224_ (_26799_, _26798_, _26526_);
  nor _31225_ (_26800_, _26799_, _26795_);
  not _31226_ (_26801_, _26800_);
  nor _31227_ (_26802_, _26788_, _24095_);
  nor _31228_ (_26803_, _26802_, _26801_);
  nand _31229_ (_26804_, _26803_, _26789_);
  nor _31230_ (_26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31231_ (_26806_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _31232_ (_26807_, _26805_);
  nor _31233_ (_26808_, _26807_, _24575_);
  nor _31234_ (_26809_, _26808_, _26806_);
  not _31235_ (_26810_, _26809_);
  nor _31236_ (_26811_, _24508_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _31237_ (_26812_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _31238_ (_26813_, _24353_, _26812_);
  nor _31239_ (_26814_, _26813_, _26811_);
  nor _31240_ (_26815_, _26814_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _31241_ (_26816_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31242_ (_26817_, _24247_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _31243_ (_26818_, _24558_, _26812_);
  nor _31244_ (_26819_, _26818_, _26817_);
  nor _31245_ (_26820_, _26819_, _26816_);
  nor _31246_ (_26821_, _26820_, _26815_);
  nor _31247_ (_26822_, _26821_, _26810_);
  not _31248_ (_26823_, _26822_);
  nor _31249_ (_26824_, _24396_, _26812_);
  nor _31250_ (_26825_, _26824_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31251_ (_26826_, _24296_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _31252_ (_26827_, _24199_, _26812_);
  nor _31253_ (_26828_, _26827_, _26826_);
  nor _31254_ (_26829_, _26828_, _26816_);
  nor _31255_ (_26830_, _26829_, _26825_);
  nor _31256_ (_26831_, _26807_, _24557_);
  nor _31257_ (_26832_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor _31258_ (_26833_, _26832_, _26831_);
  not _31259_ (_26834_, _26833_);
  nor _31260_ (_26835_, _26834_, _26830_);
  not _31261_ (_26836_, _26821_);
  nor _31262_ (_26837_, _26836_, _26809_);
  nor _31263_ (_26838_, _26837_, _26822_);
  nand _31264_ (_26839_, _26838_, _26835_);
  nand _31265_ (_26840_, _26839_, _26823_);
  not _31266_ (_26841_, _26830_);
  nor _31267_ (_26842_, _26833_, _26841_);
  nor _31268_ (_26843_, _26842_, _26835_);
  nand _31269_ (_26844_, _26843_, _26838_);
  nor _31270_ (_26845_, _26807_, _24196_);
  nor _31271_ (_26846_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor _31272_ (_26847_, _26846_, _26845_);
  nor _31273_ (_26848_, _24434_, _26812_);
  nor _31274_ (_26849_, _26848_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31275_ (_26850_, _24353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _31276_ (_26851_, _24247_, _26812_);
  nor _31277_ (_26852_, _26851_, _26850_);
  nor _31278_ (_26853_, _26852_, _26816_);
  nor _31279_ (_26854_, _26853_, _26849_);
  not _31280_ (_26855_, _26854_);
  nand _31281_ (_26856_, _26855_, _26847_);
  nor _31282_ (_26857_, _24439_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _31283_ (_26858_, _24296_, _26812_);
  nor _31284_ (_26859_, _26858_, _26857_);
  nand _31285_ (_26860_, _26859_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _31286_ (_26861_, _26860_);
  nor _31287_ (_26862_, _26807_, _24243_);
  nor _31288_ (_26863_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  nor _31289_ (_26864_, _26863_, _26862_);
  not _31290_ (_26865_, _26864_);
  nor _31291_ (_26866_, _26865_, _26861_);
  not _31292_ (_26867_, _26847_);
  nor _31293_ (_26868_, _26854_, _26867_);
  nor _31294_ (_26869_, _26855_, _26847_);
  nor _31295_ (_26870_, _26869_, _26868_);
  nand _31296_ (_26871_, _26870_, _26866_);
  nand _31297_ (_26872_, _26871_, _26856_);
  nand _31298_ (_26873_, _26814_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31299_ (_26874_, _26807_, _24278_);
  nor _31300_ (_26875_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor _31301_ (_26876_, _26875_, _26874_);
  nand _31302_ (_26877_, _26876_, _26873_);
  not _31303_ (_26878_, _26877_);
  nor _31304_ (_26879_, _26876_, _26873_);
  not _31305_ (_26880_, _26879_);
  nand _31306_ (_26881_, _26880_, _26877_);
  nand _31307_ (_26882_, _26824_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31308_ (_26883_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor _31309_ (_26884_, _26807_, _24350_);
  nor _31310_ (_26885_, _26884_, _26883_);
  nand _31311_ (_26886_, _26885_, _26882_);
  not _31312_ (_26887_, _26886_);
  nand _31313_ (_26888_, _26848_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31314_ (_26889_, _26807_, _24380_);
  nor _31315_ (_26890_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  nor _31316_ (_26891_, _26890_, _26889_);
  nor _31317_ (_26892_, _26891_, _26888_);
  nand _31318_ (_26893_, _24439_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _31319_ (_26894_, _26893_, _26816_);
  not _31320_ (_26895_, _26883_);
  nand _31321_ (_26896_, _26805_, _24323_);
  nand _31322_ (_26897_, _26896_, _26895_);
  nand _31323_ (_26898_, _26897_, _26894_);
  nand _31324_ (_26899_, _26898_, _26886_);
  nor _31325_ (_26900_, _26899_, _26892_);
  nor _31326_ (_26901_, _26900_, _26887_);
  nor _31327_ (_26902_, _26901_, _26881_);
  nor _31328_ (_26903_, _26902_, _26878_);
  nor _31329_ (_26904_, _26864_, _26860_);
  nor _31330_ (_26905_, _26904_, _26866_);
  nand _31331_ (_26906_, _26870_, _26905_);
  nor _31332_ (_26907_, _26906_, _26903_);
  nor _31333_ (_26908_, _26907_, _26872_);
  nor _31334_ (_26909_, _26908_, _26844_);
  nor _31335_ (_26910_, _26909_, _26840_);
  nor _31336_ (_26911_, _24558_, _24576_);
  nor _31337_ (_26912_, _26911_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _31338_ (_26913_, _26912_);
  nor _31339_ (_26914_, _26828_, _26819_);
  nor _31340_ (_26915_, _24199_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _31341_ (_26916_, _24576_, _26812_);
  nor _31342_ (_26917_, _26916_, _26915_);
  nor _31343_ (_26918_, _26917_, _26852_);
  nand _31344_ (_26919_, _26918_, _26914_);
  nand _31345_ (_26920_, _26919_, _26816_);
  nand _31346_ (_26921_, _26920_, _26913_);
  nor _31347_ (_26922_, _26859_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _31348_ (_26923_, _26917_, _26816_);
  nor _31349_ (_26924_, _26923_, _26922_);
  nor _31350_ (_26925_, _26924_, _26921_);
  not _31351_ (_26926_, _26925_);
  nor _31352_ (_26927_, _26926_, _26910_);
  nor _31353_ (_26928_, _26927_, _26810_);
  not _31354_ (_26929_, _26866_);
  nand _31355_ (_26930_, _26854_, _26867_);
  nand _31356_ (_26931_, _26930_, _26856_);
  nor _31357_ (_26932_, _26931_, _26929_);
  nor _31358_ (_26933_, _26932_, _26868_);
  nor _31359_ (_26934_, _26933_, _26844_);
  nor _31360_ (_26935_, _26934_, _26840_);
  not _31361_ (_26936_, _26903_);
  nor _31362_ (_26937_, _26906_, _26844_);
  nand _31363_ (_26938_, _26937_, _26936_);
  nand _31364_ (_26939_, _26938_, _26935_);
  nand _31365_ (_26940_, _26925_, _26939_);
  not _31366_ (_26941_, _26843_);
  nor _31367_ (_26942_, _26908_, _26941_);
  nor _31368_ (_26943_, _26942_, _26835_);
  nand _31369_ (_26944_, _26943_, _26838_);
  not _31370_ (_26945_, _26944_);
  nor _31371_ (_26946_, _26943_, _26838_);
  nor _31372_ (_26947_, _26946_, _26945_);
  nor _31373_ (_26948_, _26947_, _26940_);
  nor _31374_ (_26949_, _26948_, _26928_);
  not _31375_ (_26950_, _26924_);
  not _31376_ (_26951_, _26949_);
  nor _31377_ (_26952_, _26951_, _26950_);
  nor _31378_ (_26953_, _26949_, _26924_);
  nand _31379_ (_26954_, _26908_, _26941_);
  not _31380_ (_26955_, _26954_);
  nor _31381_ (_26956_, _26955_, _26942_);
  nor _31382_ (_26957_, _26956_, _26940_);
  nor _31383_ (_26958_, _26927_, _26833_);
  nor _31384_ (_26959_, _26958_, _26957_);
  not _31385_ (_26960_, _26959_);
  nor _31386_ (_26961_, _26960_, _26821_);
  nor _31387_ (_26962_, _26961_, _26953_);
  nor _31388_ (_26963_, _26962_, _26952_);
  nor _31389_ (_26964_, _26953_, _26952_);
  not _31390_ (_26965_, _26964_);
  nor _31391_ (_26966_, _26959_, _26836_);
  nor _31392_ (_26967_, _26966_, _26961_);
  not _31393_ (_26968_, _26967_);
  nor _31394_ (_26969_, _26968_, _26965_);
  not _31395_ (_26970_, _26969_);
  nand _31396_ (_26971_, _26905_, _26936_);
  nand _31397_ (_26972_, _26971_, _26929_);
  nor _31398_ (_26973_, _26870_, _26972_);
  nand _31399_ (_26974_, _26870_, _26972_);
  not _31400_ (_26975_, _26974_);
  nor _31401_ (_26976_, _26975_, _26973_);
  nor _31402_ (_26977_, _26976_, _26940_);
  nand _31403_ (_26978_, _26940_, _26867_);
  not _31404_ (_26979_, _26978_);
  nor _31405_ (_26980_, _26979_, _26977_);
  not _31406_ (_26981_, _26980_);
  nor _31407_ (_26982_, _26981_, _26830_);
  not _31408_ (_26983_, _26982_);
  nor _31409_ (_26984_, _26905_, _26936_);
  not _31410_ (_26985_, _26984_);
  nand _31411_ (_26986_, _26985_, _26971_);
  not _31412_ (_26987_, _26986_);
  nor _31413_ (_26988_, _26987_, _26940_);
  nand _31414_ (_26989_, _26940_, _26865_);
  not _31415_ (_26990_, _26989_);
  nor _31416_ (_26991_, _26990_, _26988_);
  nand _31417_ (_26992_, _26991_, _26855_);
  not _31418_ (_26993_, _26992_);
  nor _31419_ (_26994_, _26980_, _26841_);
  nor _31420_ (_26995_, _26982_, _26994_);
  nand _31421_ (_26996_, _26995_, _26993_);
  nand _31422_ (_26997_, _26996_, _26983_);
  not _31423_ (_26998_, _26881_);
  not _31424_ (_26999_, _26901_);
  nor _31425_ (_27000_, _26999_, _26998_);
  nor _31426_ (_27001_, _27000_, _26902_);
  nor _31427_ (_27002_, _27001_, _26940_);
  not _31428_ (_27003_, _26876_);
  nand _31429_ (_27004_, _26940_, _27003_);
  not _31430_ (_27005_, _27004_);
  nor _31431_ (_27006_, _27005_, _27002_);
  nor _31432_ (_27007_, _27006_, _26860_);
  not _31433_ (_27008_, _27007_);
  nand _31434_ (_27009_, _26940_, _26891_);
  not _31435_ (_27010_, _26888_);
  nor _31436_ (_27011_, _26891_, _27010_);
  not _31437_ (_27012_, _26891_);
  nor _31438_ (_27013_, _27012_, _26888_);
  nor _31439_ (_27014_, _27013_, _27011_);
  nand _31440_ (_27015_, _26927_, _27014_);
  nand _31441_ (_27016_, _27015_, _27009_);
  nand _31442_ (_27017_, _27016_, _26882_);
  nor _31443_ (_27018_, _26927_, _27012_);
  not _31444_ (_27019_, _27014_);
  nor _31445_ (_27020_, _26940_, _27019_);
  nor _31446_ (_27021_, _27020_, _27018_);
  nor _31447_ (_27022_, _27021_, _26894_);
  nor _31448_ (_27023_, _27016_, _26882_);
  nor _31449_ (_27024_, _27023_, _27022_);
  nor _31450_ (_27025_, _26807_, _24427_);
  nor _31451_ (_27026_, _26805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _31452_ (_27027_, _27026_, _27025_);
  nor _31453_ (_27028_, _27027_, _26888_);
  not _31454_ (_27029_, _27028_);
  nand _31455_ (_27030_, _27029_, _27024_);
  nand _31456_ (_27031_, _27030_, _27017_);
  not _31457_ (_27032_, _26892_);
  not _31458_ (_27033_, _26899_);
  nor _31459_ (_27034_, _27033_, _27032_);
  nor _31460_ (_27035_, _27034_, _26900_);
  nor _31461_ (_27036_, _27035_, _26940_);
  nor _31462_ (_27037_, _26927_, _26885_);
  nor _31463_ (_27038_, _27037_, _27036_);
  nand _31464_ (_27039_, _27038_, _26873_);
  not _31465_ (_27040_, _27039_);
  nor _31466_ (_27041_, _27038_, _26873_);
  nor _31467_ (_27042_, _27041_, _27040_);
  nand _31468_ (_27043_, _27042_, _27031_);
  not _31469_ (_27044_, _27006_);
  nor _31470_ (_27045_, _27044_, _26861_);
  nor _31471_ (_27046_, _27045_, _27040_);
  nand _31472_ (_27047_, _27046_, _27043_);
  nand _31473_ (_27048_, _27047_, _27008_);
  nor _31474_ (_27049_, _26991_, _26855_);
  nor _31475_ (_27050_, _27049_, _26993_);
  nand _31476_ (_27051_, _26995_, _27050_);
  nor _31477_ (_27052_, _27051_, _27048_);
  nor _31478_ (_27053_, _27052_, _26997_);
  nor _31479_ (_27054_, _27053_, _26970_);
  nor _31480_ (_27055_, _27054_, _26963_);
  nor _31481_ (_27056_, _27055_, _26921_);
  nor _31482_ (_27057_, _27056_, _26949_);
  not _31483_ (_27058_, _26921_);
  not _31484_ (_27059_, _26963_);
  not _31485_ (_27060_, _26997_);
  nand _31486_ (_27061_, _27021_, _26894_);
  nand _31487_ (_27062_, _27061_, _27017_);
  nor _31488_ (_27063_, _27028_, _27062_);
  nor _31489_ (_27064_, _27063_, _27022_);
  not _31490_ (_27065_, _27041_);
  nand _31491_ (_27066_, _27065_, _27039_);
  nor _31492_ (_27067_, _27066_, _27064_);
  not _31493_ (_27068_, _27046_);
  nor _31494_ (_27069_, _27068_, _27067_);
  nor _31495_ (_27070_, _27069_, _27007_);
  not _31496_ (_27071_, _27051_);
  nand _31497_ (_27072_, _27071_, _27070_);
  nand _31498_ (_27073_, _27072_, _27060_);
  nand _31499_ (_27074_, _27073_, _26969_);
  nand _31500_ (_27075_, _27074_, _27059_);
  nand _31501_ (_27076_, _27075_, _27058_);
  not _31502_ (_27077_, _26961_);
  nand _31503_ (_27078_, _27073_, _26967_);
  nand _31504_ (_27079_, _27078_, _27077_);
  nor _31505_ (_27080_, _27079_, _26965_);
  nor _31506_ (_27081_, _27053_, _26968_);
  nor _31507_ (_27082_, _27081_, _26961_);
  nor _31508_ (_27083_, _27082_, _26964_);
  nor _31509_ (_27084_, _27083_, _27080_);
  nor _31510_ (_27086_, _27084_, _27076_);
  nor _31511_ (_27087_, _27086_, _27057_);
  nor _31512_ (_27088_, _27087_, _24768_);
  nor _31513_ (_27089_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _31514_ (_27090_, _27089_);
  nand _31515_ (_27091_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not _31516_ (_27092_, _27091_);
  nand _31517_ (_27093_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  nand _31518_ (_27094_, _27089_, _24555_);
  not _31519_ (_27095_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  nor _31520_ (_27096_, _27095_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _31521_ (_27097_, _27096_);
  nor _31522_ (_27098_, _27097_, _24241_);
  not _31523_ (_27099_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nor _31524_ (_27100_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _27099_);
  not _31525_ (_27101_, _27100_);
  nor _31526_ (_27102_, _27101_, _24338_);
  nor _31527_ (_27103_, _27102_, _27098_);
  nor _31528_ (_27104_, _27100_, _27096_);
  nand _31529_ (_27105_, _24434_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nand _31530_ (_27106_, _27105_, _27104_);
  nand _31531_ (_27107_, _27106_, _27103_);
  nand _31532_ (_27108_, _27107_, _27094_);
  nor _31533_ (_27109_, _27108_, _24279_);
  nand _31534_ (_27111_, _27089_, _24149_);
  nor _31535_ (_27112_, _27097_, _24194_);
  nor _31536_ (_27113_, _27101_, _24285_);
  nor _31537_ (_27114_, _27113_, _27112_);
  nand _31538_ (_27115_, _24396_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nand _31539_ (_27116_, _27115_, _27104_);
  nand _31540_ (_27117_, _27116_, _27114_);
  nand _31541_ (_27118_, _27117_, _27111_);
  nor _31542_ (_27119_, _27118_, _24224_);
  nand _31543_ (_27120_, _27119_, _27109_);
  nor _31544_ (_27121_, _27108_, _24224_);
  nor _31545_ (_27122_, _27118_, _24179_);
  nand _31546_ (_27123_, _27122_, _27121_);
  not _31547_ (_27124_, _27111_);
  nand _31548_ (_27125_, _27096_, _24199_);
  nand _31549_ (_27126_, _27100_, _24296_);
  nand _31550_ (_27127_, _27126_, _27125_);
  not _31551_ (_27129_, _27104_);
  nor _31552_ (_27130_, _24439_, _27099_);
  nor _31553_ (_27131_, _27130_, _27129_);
  nor _31554_ (_27132_, _27131_, _27127_);
  nor _31555_ (_27133_, _27132_, _27124_);
  nand _31556_ (_27134_, _27133_, _24243_);
  not _31557_ (_27135_, _27094_);
  nand _31558_ (_27136_, _27096_, _24247_);
  nand _31559_ (_27137_, _27100_, _24353_);
  nand _31560_ (_27138_, _27137_, _27136_);
  nor _31561_ (_27139_, _24508_, _27099_);
  nor _31562_ (_27140_, _27139_, _27129_);
  nor _31563_ (_27141_, _27140_, _27138_);
  nor _31564_ (_27142_, _27141_, _27135_);
  nand _31565_ (_27143_, _27142_, _24196_);
  nand _31566_ (_27144_, _27143_, _27134_);
  nand _31567_ (_27145_, _27144_, _27123_);
  nor _31568_ (_27146_, _27145_, _27120_);
  nand _31569_ (_27147_, _27133_, _24196_);
  nand _31570_ (_27148_, _27142_, _24243_);
  nor _31571_ (_27149_, _27147_, _27148_);
  nand _31572_ (_27150_, _27149_, _24557_);
  nand _31573_ (_27151_, _27142_, _24557_);
  nand _31574_ (_27152_, _27151_, _27123_);
  nand _31575_ (_27153_, _27152_, _27150_);
  nor _31576_ (_27154_, _27153_, _27147_);
  nor _31577_ (_27155_, _27108_, _24549_);
  nor _31578_ (_27157_, _27155_, _27122_);
  nor _31579_ (_27158_, _27157_, _27154_);
  nand _31580_ (_27159_, _27158_, _27146_);
  nor _31581_ (_27160_, _27123_, _24549_);
  nor _31582_ (_27161_, _27155_, _27149_);
  nor _31583_ (_27163_, _27161_, _27160_);
  nand _31584_ (_27164_, _27163_, _27122_);
  nor _31585_ (_27166_, _27118_, _24137_);
  not _31586_ (_27167_, _27166_);
  nor _31587_ (_27168_, _27167_, _27151_);
  nor _31588_ (_27169_, _27108_, _24137_);
  nor _31589_ (_27171_, _27118_, _24549_);
  nor _31590_ (_27172_, _27171_, _27169_);
  nor _31591_ (_27173_, _27172_, _27168_);
  not _31592_ (_27174_, _27173_);
  nor _31593_ (_27175_, _27174_, _27164_);
  nor _31594_ (_27176_, _27173_, _27154_);
  nor _31595_ (_27177_, _27176_, _27175_);
  nand _31596_ (_27178_, _27177_, _27160_);
  nand _31597_ (_27179_, _27173_, _27154_);
  nand _31598_ (_27180_, _27174_, _27164_);
  nand _31599_ (_27181_, _27180_, _27179_);
  nand _31600_ (_27182_, _27181_, _27150_);
  nand _31601_ (_27183_, _27182_, _27178_);
  nor _31602_ (_27184_, _27183_, _27159_);
  nand _31603_ (_27185_, _27133_, _24380_);
  nand _31604_ (_27186_, _27142_, _24350_);
  nor _31605_ (_27187_, _27186_, _27185_);
  nand _31606_ (_27188_, _27142_, _24278_);
  nand _31607_ (_27189_, _27142_, _24380_);
  nor _31608_ (_27190_, _27118_, _24323_);
  nand _31609_ (_27191_, _27190_, _27189_);
  nor _31610_ (_27192_, _27191_, _27188_);
  nor _31611_ (_27193_, _27192_, _27187_);
  nand _31612_ (_27194_, _27133_, _24278_);
  nand _31613_ (_27195_, _27194_, _27148_);
  nand _31614_ (_27196_, _27195_, _27120_);
  nor _31615_ (_27197_, _27196_, _27193_);
  nor _31616_ (_27198_, _27134_, _27188_);
  nor _31617_ (_27199_, _27108_, _24179_);
  nor _31618_ (_27200_, _27199_, _27119_);
  nor _31619_ (_27201_, _27200_, _27149_);
  nor _31620_ (_27202_, _27201_, _27198_);
  nor _31621_ (_27203_, _27202_, _27146_);
  nand _31622_ (_27204_, _27203_, _27197_);
  nand _31623_ (_27205_, _27201_, _27198_);
  not _31624_ (_27206_, _27157_);
  nand _31625_ (_27207_, _27206_, _27164_);
  nand _31626_ (_27208_, _27207_, _27205_);
  nand _31627_ (_27209_, _27208_, _27159_);
  nor _31628_ (_27210_, _27209_, _27204_);
  nor _31629_ (_27211_, _27108_, _24381_);
  nor _31630_ (_27212_, _27118_, _24428_);
  nand _31631_ (_27213_, _27212_, _27211_);
  nor _31632_ (_27214_, _27118_, _24381_);
  nor _31633_ (_27215_, _27108_, _24323_);
  nand _31634_ (_27216_, _27215_, _27214_);
  nand _31635_ (_27217_, _27186_, _27185_);
  nand _31636_ (_27218_, _27217_, _27216_);
  nor _31637_ (_27219_, _27218_, _27213_);
  nand _31638_ (_27220_, _27133_, _24350_);
  nor _31639_ (_27221_, _27220_, _27211_);
  nor _31640_ (_27222_, _27221_, _27109_);
  nor _31641_ (_27223_, _27222_, _27192_);
  nand _31642_ (_27224_, _27223_, _27219_);
  nand _31643_ (_27225_, _27221_, _27109_);
  nand _31644_ (_27226_, _27225_, _27216_);
  nor _31645_ (_27227_, _27118_, _24279_);
  nor _31646_ (_27228_, _27227_, _27121_);
  nor _31647_ (_27229_, _27228_, _27198_);
  nand _31648_ (_27230_, _27229_, _27226_);
  nand _31649_ (_27231_, _27196_, _27193_);
  nand _31650_ (_27232_, _27231_, _27230_);
  nor _31651_ (_27233_, _27232_, _27224_);
  nand _31652_ (_27234_, _27145_, _27120_);
  nand _31653_ (_27235_, _27234_, _27205_);
  nor _31654_ (_27236_, _27235_, _27230_);
  nor _31655_ (_27237_, _27203_, _27197_);
  nor _31656_ (_27238_, _27237_, _27236_);
  nand _31657_ (_27239_, _27238_, _27233_);
  nor _31658_ (_27240_, _27207_, _27205_);
  nor _31659_ (_27241_, _27158_, _27146_);
  nor _31660_ (_27242_, _27241_, _27240_);
  nand _31661_ (_27243_, _27242_, _27236_);
  nand _31662_ (_27244_, _27209_, _27204_);
  nand _31663_ (_27245_, _27244_, _27243_);
  nor _31664_ (_27246_, _27245_, _27239_);
  nor _31665_ (_27247_, _27246_, _27210_);
  nor _31666_ (_27248_, _27181_, _27150_);
  nor _31667_ (_27249_, _27177_, _27160_);
  nor _31668_ (_27250_, _27249_, _27248_);
  nand _31669_ (_27251_, _27250_, _27240_);
  nand _31670_ (_27252_, _27183_, _27159_);
  nand _31671_ (_27253_, _27252_, _27251_);
  nor _31672_ (_27254_, _27253_, _27247_);
  nor _31673_ (_27255_, _27254_, _27184_);
  nor _31674_ (_27256_, _27167_, _27155_);
  not _31675_ (_27258_, _27256_);
  nor _31676_ (_27259_, _27248_, _27175_);
  nor _31677_ (_27261_, _27259_, _27258_);
  not _31678_ (_27262_, _27261_);
  nand _31679_ (_27263_, _27259_, _27258_);
  nand _31680_ (_27264_, _27263_, _27262_);
  nor _31681_ (_27265_, _27264_, _27255_);
  nor _31682_ (_27266_, _27261_, _27168_);
  not _31683_ (_27267_, _27266_);
  nor _31684_ (_27268_, _27267_, _27265_);
  nor _31685_ (_27269_, _27268_, _27093_);
  not _31686_ (_27270_, _27093_);
  nor _31687_ (_27271_, _27108_, _24428_);
  not _31688_ (_27272_, _27271_);
  nor _31689_ (_27273_, _27272_, _27185_);
  nor _31690_ (_27274_, _27215_, _27214_);
  nor _31691_ (_27275_, _27274_, _27187_);
  nand _31692_ (_27276_, _27275_, _27273_);
  nand _31693_ (_27277_, _27191_, _27188_);
  nand _31694_ (_27278_, _27277_, _27225_);
  nor _31695_ (_27279_, _27278_, _27276_);
  nor _31696_ (_27280_, _27229_, _27226_);
  nor _31697_ (_27281_, _27280_, _27197_);
  nand _31698_ (_27282_, _27281_, _27279_);
  nand _31699_ (_27283_, _27235_, _27230_);
  nand _31700_ (_27284_, _27283_, _27204_);
  nor _31701_ (_27285_, _27284_, _27282_);
  nor _31702_ (_27286_, _27242_, _27236_);
  nor _31703_ (_27287_, _27286_, _27210_);
  nand _31704_ (_27288_, _27287_, _27285_);
  nand _31705_ (_27289_, _27288_, _27243_);
  nor _31706_ (_27290_, _27250_, _27240_);
  nor _31707_ (_27291_, _27290_, _27184_);
  nand _31708_ (_27292_, _27291_, _27289_);
  nand _31709_ (_27293_, _27292_, _27251_);
  not _31710_ (_27294_, _27264_);
  nand _31711_ (_27295_, _27294_, _27293_);
  nand _31712_ (_27296_, _27266_, _27295_);
  nand _31713_ (_27297_, _27296_, _27270_);
  nand _31714_ (_27298_, _27268_, _27093_);
  nand _31715_ (_27299_, _27298_, _27297_);
  nand _31716_ (_27300_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  not _31717_ (_27301_, _27300_);
  nor _31718_ (_27302_, _27294_, _27293_);
  nor _31719_ (_27303_, _27302_, _27265_);
  nand _31720_ (_27304_, _27303_, _27301_);
  nor _31721_ (_27305_, _27304_, _27299_);
  nor _31722_ (_27306_, _27305_, _27269_);
  nand _31723_ (_27307_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  nand _31724_ (_27308_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor _31725_ (_27309_, _27308_, _27307_);
  not _31726_ (_27310_, _27309_);
  nor _31727_ (_27311_, _27310_, _27306_);
  nand _31728_ (_27312_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  not _31729_ (_27313_, _27312_);
  nor _31730_ (_27314_, _27291_, _27289_);
  nor _31731_ (_27315_, _27314_, _27254_);
  nand _31732_ (_27316_, _27315_, _27313_);
  not _31733_ (_27317_, _27316_);
  nand _31734_ (_27318_, _27253_, _27247_);
  nand _31735_ (_27319_, _27318_, _27292_);
  nand _31736_ (_27320_, _27319_, _27312_);
  nand _31737_ (_27321_, _27320_, _27316_);
  nand _31738_ (_27322_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  not _31739_ (_27323_, _27322_);
  nor _31740_ (_27324_, _27287_, _27285_);
  nor _31741_ (_27325_, _27324_, _27246_);
  nand _31742_ (_27326_, _27325_, _27323_);
  not _31743_ (_27327_, _27326_);
  nand _31744_ (_27328_, _27245_, _27239_);
  nand _31745_ (_27329_, _27328_, _27288_);
  nand _31746_ (_27330_, _27329_, _27322_);
  nand _31747_ (_27331_, _27330_, _27326_);
  nand _31748_ (_27332_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  not _31749_ (_27333_, _27332_);
  nor _31750_ (_27334_, _27238_, _27233_);
  nor _31751_ (_27335_, _27334_, _27285_);
  nand _31752_ (_27336_, _27335_, _27333_);
  not _31753_ (_27338_, _27336_);
  nand _31754_ (_27339_, _27284_, _27282_);
  nand _31755_ (_27340_, _27339_, _27239_);
  nand _31756_ (_27342_, _27340_, _27332_);
  nand _31757_ (_27344_, _27342_, _27336_);
  nand _31758_ (_27345_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  not _31759_ (_27346_, _27345_);
  nor _31760_ (_27347_, _27281_, _27279_);
  nor _31761_ (_27348_, _27347_, _27233_);
  nand _31762_ (_27349_, _27348_, _27346_);
  not _31763_ (_27350_, _27349_);
  nand _31764_ (_27351_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  not _31765_ (_27352_, _27351_);
  nor _31766_ (_27353_, _27223_, _27219_);
  nor _31767_ (_27354_, _27353_, _27279_);
  nand _31768_ (_27355_, _27354_, _27352_);
  not _31769_ (_27356_, _27355_);
  nand _31770_ (_27357_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  not _31771_ (_27358_, _27357_);
  nor _31772_ (_27359_, _27275_, _27273_);
  nor _31773_ (_27360_, _27359_, _27219_);
  nand _31774_ (_27361_, _27360_, _27358_);
  nand _31775_ (_27362_, _27278_, _27276_);
  nand _31776_ (_27363_, _27362_, _27224_);
  nand _31777_ (_27365_, _27363_, _27351_);
  nand _31778_ (_27366_, _27365_, _27355_);
  nor _31779_ (_27367_, _27366_, _27361_);
  nor _31780_ (_27369_, _27367_, _27356_);
  nand _31781_ (_27370_, _27232_, _27224_);
  nand _31782_ (_27371_, _27370_, _27282_);
  nand _31783_ (_27372_, _27371_, _27345_);
  nand _31784_ (_27373_, _27372_, _27349_);
  nor _31785_ (_27375_, _27373_, _27369_);
  nor _31786_ (_27376_, _27375_, _27350_);
  nor _31787_ (_27377_, _27376_, _27344_);
  nor _31788_ (_27378_, _27377_, _27338_);
  nor _31789_ (_27379_, _27378_, _27331_);
  nor _31790_ (_27380_, _27379_, _27327_);
  nor _31791_ (_27381_, _27380_, _27321_);
  nor _31792_ (_27382_, _27381_, _27317_);
  nand _31793_ (_27383_, _27264_, _27255_);
  nand _31794_ (_27384_, _27383_, _27295_);
  nand _31795_ (_27385_, _27384_, _27300_);
  nand _31796_ (_27386_, _27385_, _27304_);
  nor _31797_ (_27387_, _27386_, _27299_);
  nand _31798_ (_27388_, _27309_, _27387_);
  nor _31799_ (_27389_, _27388_, _27382_);
  nor _31800_ (_27390_, _27389_, _27311_);
  nand _31801_ (_27391_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  nand _31802_ (_27392_, _27090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _31803_ (_27393_, _27392_, _27391_);
  not _31804_ (_27394_, _27393_);
  nor _31805_ (_27395_, _27394_, _27390_);
  nand _31806_ (_27396_, _27395_, _27092_);
  not _31807_ (_27397_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _31808_ (_27398_, _27089_, _27397_);
  nand _31809_ (_27399_, _27398_, _27396_);
  nor _31810_ (_27400_, _27296_, _27270_);
  nor _31811_ (_27401_, _27400_, _27269_);
  nor _31812_ (_27402_, _27384_, _27300_);
  nand _31813_ (_27403_, _27402_, _27401_);
  nand _31814_ (_27404_, _27403_, _27297_);
  nand _31815_ (_27405_, _27309_, _27404_);
  not _31816_ (_27406_, _27382_);
  nor _31817_ (_27407_, _27303_, _27301_);
  nor _31818_ (_27408_, _27407_, _27402_);
  nand _31819_ (_27409_, _27408_, _27401_);
  nor _31820_ (_27410_, _27310_, _27409_);
  nand _31821_ (_27411_, _27410_, _27406_);
  nand _31822_ (_27412_, _27411_, _27405_);
  nand _31823_ (_27413_, _27393_, _27412_);
  nor _31824_ (_27414_, _27413_, _27091_);
  nand _31825_ (_27415_, _27414_, _27397_);
  nand _31826_ (_27416_, _27415_, _27399_);
  nand _31827_ (_27417_, _27416_, _24770_);
  nand _31828_ (_27418_, _26155_, _24590_);
  not _31829_ (_27420_, _27418_);
  not _31830_ (_27421_, _24574_);
  nor _31831_ (_27423_, _24578_, _27421_);
  nor _31832_ (_27424_, _27423_, _24580_);
  nand _31833_ (_27425_, _27424_, _24088_);
  not _31834_ (_27426_, _24657_);
  nor _31835_ (_27427_, _27426_, _24651_);
  nor _31836_ (_27429_, _27427_, _24497_);
  not _31837_ (_27430_, _27429_);
  nor _31838_ (_27431_, _27430_, _24654_);
  not _31839_ (_27432_, _27427_);
  nor _31840_ (_27433_, _27432_, _24224_);
  not _31841_ (_27434_, _27433_);
  nand _31842_ (_27436_, _27434_, _24653_);
  nor _31843_ (_27437_, _27429_, _27436_);
  nor _31844_ (_27438_, _27437_, _27431_);
  not _31845_ (_27439_, _27438_);
  nor _31846_ (_27441_, _27439_, _24575_);
  nor _31847_ (_27442_, _27438_, _24137_);
  nor _31848_ (_27443_, _27442_, _27441_);
  nor _31849_ (_27444_, _27443_, _24651_);
  nor _31850_ (_27445_, _24703_, _24498_);
  not _31851_ (_27446_, _27445_);
  not _31852_ (_27447_, _24668_);
  nor _31853_ (_27448_, _27447_, _24137_);
  nand _31854_ (_27449_, _24697_, _24427_);
  nand _31855_ (_27450_, _24775_, _24557_);
  nand _31856_ (_27451_, _27450_, _27449_);
  nor _31857_ (_27452_, _27451_, _27448_);
  nand _31858_ (_27453_, _27452_, _27446_);
  nor _31859_ (_27454_, _27453_, _24766_);
  nand _31860_ (_27455_, _27454_, _24756_);
  nor _31861_ (_27456_, _27455_, _27444_);
  nand _31862_ (_27457_, _27456_, _27425_);
  nor _31863_ (_27458_, _27457_, _27420_);
  nand _31864_ (_27459_, _27458_, _27417_);
  nor _31865_ (_27460_, _27459_, _27088_);
  nor _31866_ (_27461_, _27460_, _25614_);
  nor _31867_ (_27462_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _31868_ (_27463_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _31869_ (_27464_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _31870_ (_27465_, _27464_, _27462_);
  not _31871_ (_27466_, _27465_);
  nor _31872_ (_27467_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nor _31873_ (_27468_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _31874_ (_27469_, _27468_, _27467_);
  not _31875_ (_27470_, _27469_);
  not _31876_ (_27471_, _24581_);
  nor _31877_ (_27472_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nor _31878_ (_27473_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _31879_ (_27474_, _27473_, _27472_);
  nand _31880_ (_27476_, _27474_, _27471_);
  nor _31881_ (_27477_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor _31882_ (_27478_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _31883_ (_27479_, _27478_, _27477_);
  not _31884_ (_27480_, _27479_);
  nor _31885_ (_27481_, _27480_, _27476_);
  nor _31886_ (_27482_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor _31887_ (_27483_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _31888_ (_27484_, _27483_, _27482_);
  nand _31889_ (_27485_, _27484_, _27481_);
  nor _31890_ (_27486_, _27485_, _27470_);
  nor _31891_ (_27487_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nor _31892_ (_27488_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _31893_ (_27489_, _27488_, _27487_);
  nand _31894_ (_27491_, _27489_, _27486_);
  nor _31895_ (_27492_, _27491_, _27466_);
  nor _31896_ (_27493_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nor _31897_ (_27494_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _31898_ (_27495_, _27494_, _27493_);
  nand _31899_ (_27496_, _27495_, _27492_);
  nor _31900_ (_27497_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor _31901_ (_27498_, _27463_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _31902_ (_27499_, _27498_, _27497_);
  nor _31903_ (_27500_, _27499_, _27496_);
  not _31904_ (_27502_, _27500_);
  nand _31905_ (_27503_, _27499_, _27496_);
  nand _31906_ (_27504_, _27503_, _27502_);
  nand _31907_ (_27505_, _27504_, _24088_);
  not _31908_ (_27506_, _24770_);
  not _31909_ (_27507_, _27321_);
  not _31910_ (_27508_, _27380_);
  nor _31911_ (_27509_, _27508_, _27507_);
  nor _31912_ (_27510_, _27509_, _27381_);
  not _31913_ (_27511_, _27510_);
  nor _31914_ (_27512_, _27511_, _27506_);
  not _31915_ (_27514_, _27512_);
  nor _31916_ (_27515_, _24737_, _24137_);
  nand _31917_ (_27516_, _27515_, _24508_);
  nor _31918_ (_27517_, _27516_, _24396_);
  not _31919_ (_27519_, _27517_);
  nor _31920_ (_27520_, _27519_, _24338_);
  not _31921_ (_27521_, _27520_);
  nor _31922_ (_27522_, _27521_, _24285_);
  nand _31923_ (_27523_, _27522_, _24247_);
  nor _31924_ (_27524_, _27523_, _24194_);
  nor _31925_ (_27525_, _27524_, _24497_);
  nor _31926_ (_27526_, _24508_, _24575_);
  nand _31927_ (_27527_, _27526_, _24729_);
  nor _31928_ (_27528_, _27527_, _24439_);
  not _31929_ (_27529_, _27528_);
  nor _31930_ (_27530_, _27529_, _24353_);
  not _31931_ (_27531_, _27530_);
  nor _31932_ (_27532_, _27531_, _24296_);
  nor _31933_ (_27533_, _24247_, _24199_);
  nand _31934_ (_27534_, _27533_, _27532_);
  nand _31935_ (_27535_, _27534_, _24497_);
  not _31936_ (_27536_, _27535_);
  nor _31937_ (_27537_, _27536_, _27525_);
  nor _31938_ (_27538_, _24558_, _24497_);
  nor _31939_ (_27539_, _27538_, _25123_);
  nand _31940_ (_27540_, _27539_, _27537_);
  nor _31941_ (_27541_, _27540_, _24149_);
  nand _31942_ (_27542_, _27540_, _24149_);
  nand _31943_ (_27543_, _27542_, _24742_);
  nor _31944_ (_27544_, _27543_, _27541_);
  nor _31945_ (_27545_, _24700_, _24279_);
  nand _31946_ (_27546_, _24767_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  not _31947_ (_27547_, _27546_);
  nor _31948_ (_27548_, _27547_, _27545_);
  nor _31949_ (_27549_, _27447_, _24149_);
  not _31950_ (_27550_, _27549_);
  nand _31951_ (_27551_, _27550_, _24751_);
  nor _31952_ (_27552_, _24498_, _24137_);
  not _31953_ (_27553_, _27552_);
  not _31954_ (_27554_, _24669_);
  nand _31955_ (_27555_, _27554_, _24576_);
  nand _31956_ (_27556_, _27555_, _27553_);
  nand _31957_ (_27557_, _27556_, _27551_);
  nand _31958_ (_27558_, _27557_, _27548_);
  nor _31959_ (_27560_, _27558_, _27544_);
  nand _31960_ (_27561_, _27560_, _27514_);
  not _31961_ (_27563_, _27561_);
  nand _31962_ (_27564_, _27563_, _27505_);
  nand _31963_ (_27565_, _27564_, _26797_);
  not _31964_ (_27566_, _26495_);
  nand _31965_ (_27567_, _27566_, _25838_);
  nand _31966_ (_27568_, _27567_, _27565_);
  nor _31967_ (_27569_, _27568_, _27461_);
  nand _31968_ (_27570_, _27569_, _26804_);
  nor _31969_ (_27571_, _26794_, _26526_);
  nand _31970_ (_27572_, _27571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _31971_ (_27573_, _27572_, _26485_);
  nor _31972_ (_27574_, _27573_, _27570_);
  not _31973_ (_27575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _31974_ (_27576_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _31975_ (_27577_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _31976_ (_27578_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _31977_ (_27579_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _31978_ (_27580_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _31979_ (_27581_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _31980_ (_27582_, _24931_);
  nor _31981_ (_27583_, _27582_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _31982_ (_27584_, _27583_, _24864_);
  nor _31983_ (_27586_, _27584_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _31984_ (_27587_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _31985_ (_27589_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _31986_ (_27590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not _31987_ (_27591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _31988_ (_27592_, _27591_, _27590_);
  not _31989_ (_27594_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not _31990_ (_27595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _31991_ (_27596_, _27595_, _27594_);
  nand _31992_ (_27597_, _27596_, _27592_);
  nor _31993_ (_27598_, _27597_, _27589_);
  not _31994_ (_27599_, _27598_);
  nor _31995_ (_27600_, _27599_, _27587_);
  nand _31996_ (_27601_, _27600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _31997_ (_27602_, _27601_, _27586_);
  not _31998_ (_27603_, _27602_);
  nor _31999_ (_27604_, _27603_, _27581_);
  not _32000_ (_27605_, _27604_);
  nor _32001_ (_27606_, _27605_, _27580_);
  not _32002_ (_27607_, _27606_);
  nor _32003_ (_27608_, _27607_, _27579_);
  not _32004_ (_27609_, _27608_);
  nor _32005_ (_27610_, _27609_, _27578_);
  not _32006_ (_27611_, _27610_);
  nor _32007_ (_27612_, _27611_, _27577_);
  not _32008_ (_27613_, _27612_);
  nor _32009_ (_27614_, _27613_, _27576_);
  nor _32010_ (_27615_, _27614_, _27575_);
  not _32011_ (_27616_, _27614_);
  nor _32012_ (_27617_, _27616_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _32013_ (_27618_, _27617_, _27615_);
  nand _32014_ (_27619_, _27618_, _26486_);
  nand _32015_ (_27620_, _27619_, _26487_);
  nor _32016_ (_28211_[15], _27620_, _27574_);
  nor _32017_ (_27622_, rst, _24858_);
  nand _32018_ (_27624_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _32019_ (_27625_, _27594_, _24936_);
  not _32020_ (_27626_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _32021_ (_27628_, _27626_, _24960_);
  not _32022_ (_27629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _32023_ (_27631_, _27629_, _24938_);
  not _32024_ (_27632_, _27631_);
  nor _32025_ (_27633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _32026_ (_27634_, _27633_, _27628_);
  not _32027_ (_27635_, _27634_);
  nor _32028_ (_27636_, _27635_, _27632_);
  nor _32029_ (_27637_, _27636_, _27628_);
  nor _32030_ (_27638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _32031_ (_27639_, _27638_, _27625_);
  not _32032_ (_27640_, _27639_);
  nor _32033_ (_27641_, _27640_, _27637_);
  nor _32034_ (_27642_, _27641_, _27625_);
  not _32035_ (_27643_, _27642_);
  nor _32036_ (_27644_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not _32037_ (_27645_, _27644_);
  nor _32038_ (_27646_, _27645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not _32039_ (_27647_, _27646_);
  nor _32040_ (_27648_, _27647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _32041_ (_27649_, _27648_);
  nor _32042_ (_27650_, _27649_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _32043_ (_27651_, _27650_);
  nor _32044_ (_27652_, _27651_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _32045_ (_27653_, _27652_);
  nor _32046_ (_27654_, _27653_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _32047_ (_27656_, _27654_);
  nor _32048_ (_27657_, _27656_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _32049_ (_27659_, _27657_);
  nor _32050_ (_27660_, _27659_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand _32051_ (_27662_, _27660_, _27578_);
  nor _32052_ (_27663_, _27662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _32053_ (_27664_, _27663_);
  nor _32054_ (_27666_, _27664_, _27643_);
  not _32055_ (_27667_, _27666_);
  nor _32056_ (_27669_, _27667_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _32057_ (_27670_, _27669_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _32058_ (_27671_, _27669_);
  nor _32059_ (_27672_, _27671_, _27575_);
  nor _32060_ (_27673_, _27672_, _27670_);
  not _32061_ (_27674_, _27673_);
  nor _32062_ (_27675_, _27666_, _27576_);
  nor _32063_ (_27676_, _27675_, _27669_);
  nor _32064_ (_27677_, _27643_, _27662_);
  nor _32065_ (_27678_, _27677_, _27577_);
  nor _32066_ (_27679_, _27678_, _27666_);
  not _32067_ (_27680_, _27679_);
  nor _32068_ (_27681_, _27643_, _27659_);
  not _32069_ (_27682_, _27681_);
  nor _32070_ (_27683_, _27682_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _32071_ (_27684_, _27683_, _27578_);
  nor _32072_ (_27685_, _27684_, _27677_);
  nor _32073_ (_27686_, _27681_, _27579_);
  nor _32074_ (_27687_, _27686_, _27683_);
  not _32075_ (_27688_, _27687_);
  nor _32076_ (_27689_, _27643_, _27656_);
  nor _32077_ (_27691_, _27689_, _27580_);
  nor _32078_ (_27692_, _27691_, _27681_);
  nor _32079_ (_27694_, _27643_, _27653_);
  nor _32080_ (_27695_, _27694_, _27581_);
  nor _32081_ (_27696_, _27695_, _27689_);
  not _32082_ (_27698_, _27696_);
  not _32083_ (_27699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _32084_ (_27700_, _27643_, _27651_);
  nor _32085_ (_27701_, _27700_, _27699_);
  nor _32086_ (_27703_, _27701_, _27694_);
  nor _32087_ (_27704_, _27643_, _27649_);
  nor _32088_ (_27705_, _27704_, _27587_);
  nor _32089_ (_27707_, _27705_, _27700_);
  not _32090_ (_27708_, _27707_);
  nor _32091_ (_27709_, _27643_, _27647_);
  nor _32092_ (_27710_, _27709_, _27589_);
  nor _32093_ (_27711_, _27710_, _27704_);
  nor _32094_ (_27712_, _27643_, _27645_);
  nor _32095_ (_27713_, _27712_, _27595_);
  nor _32096_ (_27714_, _27713_, _27709_);
  not _32097_ (_27715_, _27714_);
  nor _32098_ (_27716_, _27642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not _32099_ (_27717_, _27716_);
  nand _32100_ (_27719_, _27642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand _32101_ (_27720_, _27719_, _27717_);
  not _32102_ (_27721_, _27720_);
  nor _32103_ (_27722_, _25290_, _25262_);
  not _32104_ (_27723_, _27722_);
  not _32105_ (_27724_, _25231_);
  nor _32106_ (_27725_, _27724_, _25453_);
  not _32107_ (_27726_, _27725_);
  nor _32108_ (_27727_, _27726_, _27723_);
  not _32109_ (_27728_, _27727_);
  not _32110_ (_27729_, _25351_);
  nor _32111_ (_27730_, _27729_, _24972_);
  not _32112_ (_27731_, _27730_);
  not _32113_ (_27732_, _25383_);
  not _32114_ (_27733_, _25322_);
  nor _32115_ (_27734_, _27733_, _27732_);
  nor _32116_ (_27735_, _25322_, _25383_);
  nor _32117_ (_27736_, _27735_, _27734_);
  not _32118_ (_27737_, _27736_);
  nor _32119_ (_27738_, _27737_, _27731_);
  nor _32120_ (_27739_, _25351_, _24973_);
  not _32121_ (_27740_, _27739_);
  not _32122_ (_27741_, _27734_);
  nor _32123_ (_27742_, _27741_, _27740_);
  nor _32124_ (_27743_, _27733_, _25383_);
  not _32125_ (_27744_, _27743_);
  nor _32126_ (_27745_, _27729_, _24973_);
  not _32127_ (_27746_, _27745_);
  nor _32128_ (_27747_, _27746_, _27744_);
  nor _32129_ (_27748_, _27747_, _27742_);
  not _32130_ (_27749_, _27748_);
  nor _32131_ (_27750_, _27749_, _27738_);
  nor _32132_ (_27751_, _27750_, _27728_);
  not _32133_ (_27752_, _27735_);
  nor _32134_ (_27753_, _27752_, _27740_);
  not _32135_ (_27754_, _25262_);
  not _32136_ (_27755_, _25290_);
  nor _32137_ (_27756_, _27755_, _27754_);
  not _32138_ (_27757_, _27756_);
  nand _32139_ (_27758_, _27723_, _27757_);
  not _32140_ (_27759_, _27758_);
  nor _32141_ (_27760_, _27759_, _27726_);
  nand _32142_ (_27761_, _27760_, _27753_);
  not _32143_ (_27762_, _27761_);
  not _32144_ (_27763_, _25453_);
  nor _32145_ (_27764_, _27757_, _27724_);
  not _32146_ (_27765_, _27764_);
  nor _32147_ (_27766_, _27765_, _27763_);
  not _32148_ (_27767_, _27766_);
  nor _32149_ (_27768_, _27746_, _27741_);
  nor _32150_ (_27769_, _27768_, _27753_);
  nor _32151_ (_27770_, _27769_, _27767_);
  nor _32152_ (_27771_, _27770_, _27762_);
  not _32153_ (_27772_, _27771_);
  nor _32154_ (_27773_, _27772_, _27751_);
  not _32155_ (_27774_, _27773_);
  nor _32156_ (_27775_, _27744_, _27731_);
  nor _32157_ (_27776_, _27746_, _27752_);
  nor _32158_ (_27777_, _27776_, _27775_);
  nor _32159_ (_27778_, _27777_, _27767_);
  not _32160_ (_27779_, _27775_);
  nor _32161_ (_27780_, _27765_, _25453_);
  not _32162_ (_27781_, _27780_);
  nor _32163_ (_27782_, _27781_, _27779_);
  nor _32164_ (_27783_, _27723_, _27724_);
  nand _32165_ (_27784_, _27783_, _25453_);
  not _32166_ (_27785_, _27753_);
  nor _32167_ (_27786_, _27785_, _27784_);
  nor _32168_ (_27787_, _27786_, _27782_);
  not _32169_ (_27788_, _27787_);
  nor _32170_ (_27789_, _27788_, _27778_);
  nand _32171_ (_27790_, _25231_, _25262_);
  nor _32172_ (_27791_, _27790_, _25290_);
  not _32173_ (_27792_, _27791_);
  nor _32174_ (_27793_, _27752_, _27731_);
  nor _32175_ (_27794_, _27793_, _25453_);
  nor _32176_ (_27795_, _27794_, _27792_);
  nor _32177_ (_27796_, _27740_, _27732_);
  not _32178_ (_27797_, _27796_);
  nor _32179_ (_27798_, _25322_, _27724_);
  not _32180_ (_27799_, _27798_);
  nor _32181_ (_27800_, _27799_, _27797_);
  nand _32182_ (_27801_, _27800_, _27758_);
  not _32183_ (_27802_, _27801_);
  nor _32184_ (_27803_, _27802_, _27795_);
  nand _32185_ (_27804_, _27803_, _27789_);
  nor _32186_ (_27805_, _27804_, _27774_);
  nor _32187_ (_27806_, _27792_, _25453_);
  nor _32188_ (_27807_, _25351_, _24972_);
  not _32189_ (_27808_, _27807_);
  nor _32190_ (_27809_, _27737_, _27808_);
  nand _32191_ (_27811_, _27809_, _27806_);
  nand _32192_ (_27812_, _27747_, _27766_);
  nand _32193_ (_27813_, _27812_, _27811_);
  nor _32194_ (_27814_, _27741_, _27731_);
  not _32195_ (_27815_, _27814_);
  nor _32196_ (_27816_, _27815_, _27781_);
  nor _32197_ (_27817_, _27816_, _27813_);
  not _32198_ (_27818_, _27806_);
  nand _32199_ (_27819_, _27730_, _27733_);
  nor _32200_ (_27820_, _27819_, _27732_);
  nor _32201_ (_27822_, _27746_, _25383_);
  nor _32202_ (_27823_, _27822_, _27820_);
  nor _32203_ (_27824_, _27823_, _27818_);
  nor _32204_ (_27825_, _27740_, _27744_);
  not _32205_ (_27826_, _27825_);
  nor _32206_ (_27827_, _27760_, _27766_);
  nor _32207_ (_27828_, _27827_, _27826_);
  nor _32208_ (_27829_, _27828_, _27824_);
  nand _32209_ (_27830_, _27829_, _27817_);
  not _32210_ (_27831_, _27742_);
  nor _32211_ (_27832_, _27818_, _27831_);
  not _32212_ (_27833_, _27793_);
  nor _32213_ (_27834_, _27833_, _27728_);
  nor _32214_ (_27835_, _27834_, _27832_);
  nor _32215_ (_27836_, _27831_, _27781_);
  nand _32216_ (_27837_, _27733_, _25383_);
  nor _32217_ (_27838_, _27746_, _27837_);
  nand _32218_ (_27839_, _27838_, _27766_);
  not _32219_ (_27840_, _27839_);
  nor _32220_ (_27841_, _27840_, _27836_);
  nand _32221_ (_27843_, _27841_, _27835_);
  nor _32222_ (_27844_, _27755_, _25262_);
  nor _32223_ (_27845_, _27733_, _27724_);
  nand _32224_ (_27846_, _27845_, _27844_);
  nor _32225_ (_27847_, _27846_, _27797_);
  nor _32226_ (_27848_, _27731_, _27732_);
  not _32227_ (_27849_, _27848_);
  nor _32228_ (_27850_, _27846_, _27849_);
  nor _32229_ (_27851_, _27808_, _27732_);
  not _32230_ (_27852_, _27851_);
  nor _32231_ (_27853_, _27852_, _27781_);
  nor _32232_ (_27854_, _27853_, _27850_);
  not _32233_ (_27855_, _27854_);
  nor _32234_ (_27856_, _27855_, _27847_);
  not _32235_ (_27857_, _27856_);
  nor _32236_ (_27858_, _27857_, _27843_);
  not _32237_ (_27859_, _27858_);
  nor _32238_ (_27860_, _27859_, _27830_);
  nand _32239_ (_27861_, _27860_, _27805_);
  nor _32240_ (_27862_, _27814_, _27776_);
  nor _32241_ (_27863_, _27862_, _27728_);
  nor _32242_ (_27864_, _27826_, _27784_);
  nor _32243_ (_27865_, _27815_, _27767_);
  nor _32244_ (_27866_, _27865_, _27864_);
  nor _32245_ (_27867_, _27833_, _25231_);
  not _32246_ (_27868_, _27844_);
  nor _32247_ (_27869_, _27799_, _27868_);
  nand _32248_ (_27870_, _27869_, _27730_);
  not _32249_ (_27871_, _27870_);
  nor _32250_ (_27872_, _27871_, _27867_);
  not _32251_ (_27873_, _27872_);
  nor _32252_ (_27874_, _27852_, _27767_);
  nor _32253_ (_27875_, _27874_, _27873_);
  nand _32254_ (_27876_, _27875_, _27866_);
  nor _32255_ (_27877_, _27876_, _27863_);
  not _32256_ (_27878_, _27877_);
  nor _32257_ (_27879_, _27808_, _25383_);
  not _32258_ (_27880_, _27879_);
  nor _32259_ (_27881_, _27728_, _27880_);
  nor _32260_ (_27882_, _27793_, _27742_);
  nor _32261_ (_27883_, _27882_, _27767_);
  nor _32262_ (_27884_, _27883_, _27881_);
  nor _32263_ (_27885_, _27880_, _27767_);
  nor _32264_ (_27886_, _27818_, _27826_);
  nor _32265_ (_27887_, _27808_, _27741_);
  not _32266_ (_27888_, _27887_);
  nor _32267_ (_27889_, _27888_, _27818_);
  nor _32268_ (_27890_, _27889_, _27886_);
  not _32269_ (_27891_, _27890_);
  nor _32270_ (_27892_, _27891_, _27885_);
  nand _32271_ (_27893_, _27892_, _27884_);
  nor _32272_ (_27894_, _27893_, _27878_);
  nor _32273_ (_27895_, _27749_, _27848_);
  nor _32274_ (_27896_, _27895_, _25231_);
  nor _32275_ (_27897_, _27785_, _27818_);
  nor _32276_ (_27898_, _27815_, _27818_);
  nor _32277_ (_27899_, _27898_, _27897_);
  nor _32278_ (_27900_, _27818_, _27779_);
  nor _32279_ (_27901_, _27837_, _27740_);
  not _32280_ (_27902_, _27901_);
  nor _32281_ (_27903_, _27902_, _27818_);
  nor _32282_ (_27904_, _27903_, _27900_);
  nand _32283_ (_27905_, _27904_, _27899_);
  nor _32284_ (_27907_, _27905_, _27896_);
  nand _32285_ (_27908_, _27907_, _27894_);
  nor _32286_ (_27909_, _27908_, _27861_);
  nor _32287_ (_27910_, _27634_, _27631_);
  nor _32288_ (_27911_, _27910_, _27636_);
  not _32289_ (_27912_, _27911_);
  nor _32290_ (_27914_, _27912_, _27909_);
  nor _32291_ (_27915_, _27844_, _27724_);
  nor _32292_ (_27916_, _27915_, _27815_);
  nand _32293_ (_27917_, _27884_, _27866_);
  nor _32294_ (_27918_, _27917_, _27916_);
  not _32295_ (_27919_, _27817_);
  nor _32296_ (_27920_, _27902_, _27784_);
  nor _32297_ (_27921_, _27920_, _27786_);
  nor _32298_ (_27922_, _27889_, _27900_);
  nand _32299_ (_27923_, _27922_, _27921_);
  nor _32300_ (_27924_, _27923_, _27919_);
  nand _32301_ (_27925_, _27924_, _27918_);
  nor _32302_ (_27926_, _27925_, _27909_);
  nor _32303_ (_27927_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _32304_ (_27928_, _27927_, _27631_);
  not _32305_ (_27929_, _27928_);
  nor _32306_ (_27930_, _27929_, _27926_);
  not _32307_ (_27931_, _27930_);
  not _32308_ (_27932_, _27909_);
  nor _32309_ (_27933_, _27911_, _27932_);
  nor _32310_ (_27934_, _27933_, _27914_);
  not _32311_ (_27935_, _27934_);
  nor _32312_ (_27936_, _27935_, _27931_);
  nor _32313_ (_27937_, _27936_, _27914_);
  nand _32314_ (_27938_, _27640_, _27637_);
  not _32315_ (_27939_, _27938_);
  nor _32316_ (_27940_, _27939_, _27641_);
  not _32317_ (_27941_, _27940_);
  nor _32318_ (_27942_, _27941_, _27937_);
  nand _32319_ (_27943_, _27942_, _27721_);
  nor _32320_ (_27944_, _27643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _32321_ (_27945_, _27944_, _27591_);
  nor _32322_ (_27946_, _27945_, _27712_);
  nor _32323_ (_27947_, _27946_, _27943_);
  nand _32324_ (_27948_, _27947_, _27715_);
  nor _32325_ (_27949_, _27948_, _27711_);
  nand _32326_ (_27950_, _27949_, _27708_);
  nor _32327_ (_27951_, _27950_, _27703_);
  nand _32328_ (_27952_, _27951_, _27698_);
  nor _32329_ (_27953_, _27952_, _27692_);
  nand _32330_ (_27954_, _27953_, _27688_);
  nor _32331_ (_27955_, _27954_, _27685_);
  nand _32332_ (_27956_, _27955_, _27680_);
  nor _32333_ (_27957_, _27956_, _27676_);
  nor _32334_ (_27958_, _27957_, _27674_);
  not _32335_ (_27959_, _27957_);
  nor _32336_ (_27960_, _27959_, _27673_);
  nor _32337_ (_27961_, _27960_, _27958_);
  nand _32338_ (_27962_, _27961_, _25834_);
  nor _32339_ (_27963_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _32340_ (_27964_, rst, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _32341_ (_27965_, _27964_);
  nor _32342_ (_27966_, _27965_, _27963_);
  nand _32343_ (_27967_, _27966_, _27962_);
  nand _32344_ (_28212_[15], _27967_, _27624_);
  nand _32345_ (_27968_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _25207_);
  nor _32346_ (_28213_, _27968_, rst);
  nor _32347_ (_28214_, rst, _25207_);
  nor _32348_ (_27969_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _32349_ (_27970_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nand _32350_ (_27971_, _27970_, _27969_);
  nor _32351_ (_27972_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _32352_ (_27973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nand _32353_ (_27974_, _27973_, _27972_);
  nor _32354_ (_27975_, _27974_, _27971_);
  not _32355_ (_27976_, _27975_);
  nand _32356_ (_27977_, _27976_, _26487_);
  nand _32357_ (_27978_, _24863_, _24858_);
  nand _32358_ (_27979_, _27978_, _28214_);
  nand _32359_ (_28215_, _27979_, _27977_);
  nand _32360_ (_27980_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _26487_);
  nor _32361_ (_27981_, _26504_, rst);
  nand _32362_ (_27982_, _27981_, _27975_);
  nand _32363_ (_28216_[7], _27982_, _27980_);
  nor _32364_ (_27983_, _27586_, _24864_);
  nor _32365_ (_27984_, _27909_, _24960_);
  nor _32366_ (_27986_, _27926_, _24938_);
  nor _32367_ (_27987_, _27932_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _32368_ (_27988_, _27987_, _27984_);
  nand _32369_ (_27989_, _27988_, _27986_);
  not _32370_ (_27990_, _27989_);
  nor _32371_ (_27991_, _27990_, _27984_);
  nor _32372_ (_27992_, _27991_, _24864_);
  not _32373_ (_27993_, _27992_);
  nor _32374_ (_27994_, _27993_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _32375_ (_27995_, _27992_, _24936_);
  nor _32376_ (_27996_, _27995_, _27994_);
  nor _32377_ (_27997_, _27996_, _27983_);
  not _32378_ (_27998_, _27983_);
  nand _32379_ (_27999_, _24939_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _32380_ (_28000_, _27999_, _27998_);
  nand _32381_ (_28001_, _28000_, _27925_);
  nand _32382_ (_28002_, _28001_, _24858_);
  nor _32383_ (_28003_, _28002_, _27997_);
  nor _32384_ (_28217_[2], _28003_, rst);
  nor _32385_ (_28004_, _25287_, _25450_);
  nand _32386_ (_28005_, _28004_, _25380_);
  not _32387_ (_28006_, _25347_);
  not _32388_ (_28007_, _25258_);
  nand _32389_ (_28008_, _25319_, _28007_);
  nor _32390_ (_28009_, _28008_, _28006_);
  not _32391_ (_28010_, _25226_);
  nor _32392_ (_28011_, _25268_, rst);
  nand _32393_ (_28012_, _28011_, _28010_);
  nor _32394_ (_28013_, _28012_, _24968_);
  nand _32395_ (_28014_, _28013_, _28009_);
  nor _32396_ (_28220_, _28014_, _28005_);
  nor _32397_ (_28015_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _32398_ (_28016_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _32399_ (_28017_, _28016_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _32400_ (_28019_, _28017_, _26487_);
  nor _32401_ (_28221_[7], _28019_, _28015_);
  not _32402_ (_28020_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _32403_ (_28222_, rst, _28020_);
  not _32404_ (_28021_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nand _32405_ (_28022_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  not _32406_ (_28023_, _28022_);
  nor _32407_ (_28024_, _28023_, _28021_);
  not _32408_ (_28025_, _28024_);
  nand _32409_ (_28026_, _28023_, _28021_);
  nand _32410_ (_28027_, _28026_, _28025_);
  not _32411_ (_28028_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  not _32412_ (_28029_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  nor _32413_ (_28030_, _28029_, _28021_);
  not _32414_ (_28031_, _28030_);
  nor _32415_ (_28032_, _28031_, _28028_);
  nor _32416_ (_28033_, _28030_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _32417_ (_28034_, _28033_, _28032_);
  nor _32418_ (_28035_, _28034_, _28023_);
  not _32419_ (_28036_, _28035_);
  nand _32420_ (_28037_, _28036_, _28027_);
  nor _32421_ (_28038_, _28024_, _28029_);
  nor _32422_ (_28039_, _28025_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  nor _32423_ (_28040_, _28039_, _28038_);
  nor _32424_ (_28041_, _28032_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor _32425_ (_28224_[3], _28041_, rst);
  nand _32426_ (_28042_, _28224_[3], _28040_);
  nor _32427_ (_28223_, _28042_, _28037_);
  nor _32428_ (_28043_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  nand _32429_ (_28044_, _27586_, _26510_);
  nand _32430_ (_28045_, _28044_, _26487_);
  nor _32431_ (_28225_[31], _28045_, _28043_);
  nor _32432_ (_28046_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _32433_ (_28047_, _27586_, _25343_);
  nand _32434_ (_28048_, _28047_, _26487_);
  nor _32435_ (_28226_[31], _28048_, _28046_);
  not _32436_ (_28049_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nor _32437_ (_28050_, _28049_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor _32438_ (_28227_, _28050_, rst);
  nor _32439_ (_28051_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  nand _32440_ (_28052_, _28051_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nor _32441_ (_28229_, _28052_, rst);
  not _32442_ (_28053_, _28229_);
  nand _32443_ (_28054_, _28222_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nand _32444_ (_28228_, _28054_, _28053_);
  nand _32445_ (_28055_, _25818_, _26487_);
  nor _32446_ (_28231_, _28055_, _25527_);
  nor _32447_ (_28056_, _24887_, _24068_);
  not _32448_ (_28057_, _28056_);
  nor _32449_ (_28059_, _28057_, _24882_);
  nand _32450_ (_28060_, _28059_, _25099_);
  not _32451_ (_28061_, _28059_);
  nand _32452_ (_28062_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  nand _32453_ (_27368_, _28062_, _28060_);
  nor _32454_ (_28063_, _24993_, _24059_);
  nand _32455_ (_28064_, _28063_, _24830_);
  not _32456_ (_28065_, _28063_);
  nand _32457_ (_28066_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nand _32458_ (_27475_, _28066_, _28064_);
  nor _32459_ (_28218_[6], _25985_, rst);
  nor _32460_ (_28218_[5], _26118_, rst);
  nor _32461_ (_28218_[4], _26012_, rst);
  nor _32462_ (_28218_[3], _25912_, rst);
  nor _32463_ (_28218_[2], _26385_, rst);
  nor _32464_ (_28218_[1], _26426_, rst);
  nor _32465_ (_28218_[0], _26332_, rst);
  nor _32466_ (_28219_[6], _26553_, rst);
  nor _32467_ (_28219_[5], _26581_, rst);
  nor _32468_ (_28219_[4], _26607_, rst);
  nor _32469_ (_28219_[3], _26637_, rst);
  nor _32470_ (_28219_[2], _26667_, rst);
  nor _32471_ (_28219_[1], _26695_, rst);
  nor _32472_ (_28219_[0], _26721_, rst);
  nand _32473_ (_28068_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nand _32474_ (_28069_, _25099_, _24796_);
  nand _32475_ (_01168_, _28069_, _28068_);
  nand _32476_ (_28070_, _25166_, _25039_);
  nand _32477_ (_28071_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  nand _32478_ (_01184_, _28071_, _28070_);
  nor _32479_ (_28072_, _24976_, _24995_);
  not _32480_ (_28073_, _28072_);
  nor _32481_ (_28074_, _28073_, _25051_);
  not _32482_ (_28075_, _28074_);
  nand _32483_ (_28076_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nand _32484_ (_28077_, _28074_, _25203_);
  nand _32485_ (_01387_, _28077_, _28076_);
  nor _32486_ (_28078_, _24995_, _24001_);
  not _32487_ (_28080_, _28078_);
  nor _32488_ (_28081_, _25059_, _28080_);
  nand _32489_ (_28082_, _28081_, _25099_);
  not _32490_ (_28083_, _28081_);
  nand _32491_ (_28084_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nand _32492_ (_01411_, _28084_, _28082_);
  nor _32493_ (_28085_, _24801_, _24470_);
  nand _32494_ (_28086_, _28085_, _24716_);
  nor _32495_ (_28087_, _25703_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _32496_ (_28088_, _24470_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor _32497_ (_28089_, _24328_, _23939_);
  not _32498_ (_28091_, _28089_);
  nor _32499_ (_28092_, _28091_, _28088_);
  nor _32500_ (_28093_, _28092_, _28087_);
  nand _32501_ (_28094_, _28093_, _28086_);
  not _32502_ (_28095_, _28094_);
  nor _32503_ (_28096_, _28095_, _23918_);
  nand _32504_ (_28097_, _28096_, _24985_);
  nand _32505_ (_28098_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nand _32506_ (_01439_, _28098_, _28097_);
  nor _32507_ (_28099_, _28073_, _24993_);
  nand _32508_ (_28100_, _28099_, _25203_);
  not _32509_ (_28101_, _28099_);
  nand _32510_ (_28102_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  nand _32511_ (_01627_, _28102_, _28100_);
  nor _32512_ (_28103_, _25049_, _24982_);
  not _32513_ (_28104_, _28103_);
  nor _32514_ (_28105_, _28104_, _24795_);
  nand _32515_ (_28106_, _28105_, _24927_);
  not _32516_ (_28107_, _28105_);
  nand _32517_ (_28108_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  nand _32518_ (_02571_, _28108_, _28106_);
  nor _32519_ (_28109_, _24866_, _24401_);
  not _32520_ (_28110_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _32521_ (_28111_, _24869_, _28110_);
  nor _32522_ (_28113_, _28111_, _28109_);
  nor _32523_ (_28204_[0], _28113_, rst);
  nor _32524_ (_28114_, _24866_, _24364_);
  not _32525_ (_28115_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _32526_ (_28116_, _24869_, _28115_);
  nor _32527_ (_28117_, _28116_, _28114_);
  nor _32528_ (_28204_[1], _28117_, rst);
  nor _32529_ (_28118_, _24866_, _24305_);
  not _32530_ (_28119_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _32531_ (_28120_, _24869_, _28119_);
  nor _32532_ (_28121_, _28120_, _28118_);
  nor _32533_ (_28204_[2], _28121_, rst);
  nor _32534_ (_28122_, _24866_, _24251_);
  not _32535_ (_28123_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _32536_ (_28124_, _24869_, _28123_);
  nor _32537_ (_28125_, _28124_, _28122_);
  nor _32538_ (_28204_[3], _28125_, rst);
  nor _32539_ (_28126_, _24866_, _24202_);
  not _32540_ (_28127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _32541_ (_28128_, _24869_, _28127_);
  nor _32542_ (_28129_, _28128_, _28126_);
  nor _32543_ (_28204_[4], _28129_, rst);
  nor _32544_ (_28130_, _24866_, _24153_);
  not _32545_ (_28131_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _32546_ (_28132_, _24869_, _28131_);
  nor _32547_ (_28133_, _28132_, _28130_);
  nor _32548_ (_28204_[5], _28133_, rst);
  nor _32549_ (_28134_, _24866_, _24527_);
  not _32550_ (_00001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _32551_ (_00002_, _24869_, _00001_);
  nor _32552_ (_00004_, _00002_, _28134_);
  nor _32553_ (_28204_[6], _00004_, rst);
  nor _32554_ (_00005_, _24866_, _24090_);
  not _32555_ (_00006_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _32556_ (_00007_, _24869_, _00006_);
  nor _32557_ (_00008_, _00007_, _00005_);
  nor _32558_ (_28204_[7], _00008_, rst);
  nor _32559_ (_00009_, _24866_, _24398_);
  not _32560_ (_00010_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _32561_ (_00011_, _24869_, _00010_);
  nor _32562_ (_00012_, _00011_, _00009_);
  nor _32563_ (_28204_[8], _00012_, rst);
  nor _32564_ (_00013_, _24866_, _24374_);
  not _32565_ (_00014_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _32566_ (_00015_, _24869_, _00014_);
  nor _32567_ (_00016_, _00015_, _00013_);
  nor _32568_ (_28204_[9], _00016_, rst);
  nor _32569_ (_00017_, _24866_, _24308_);
  not _32570_ (_00018_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _32571_ (_00019_, _24869_, _00018_);
  nor _32572_ (_00021_, _00019_, _00017_);
  nor _32573_ (_28204_[10], _00021_, rst);
  nor _32574_ (_00022_, _24866_, _24253_);
  not _32575_ (_00023_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _32576_ (_00024_, _24869_, _00023_);
  nor _32577_ (_00025_, _00024_, _00022_);
  nor _32578_ (_28204_[11], _00025_, rst);
  nor _32579_ (_00026_, _24866_, _24204_);
  not _32580_ (_00027_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _32581_ (_00028_, _24869_, _00027_);
  nor _32582_ (_00029_, _00028_, _00026_);
  nor _32583_ (_28204_[12], _00029_, rst);
  nor _32584_ (_00030_, _24866_, _24151_);
  not _32585_ (_00031_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _32586_ (_00032_, _24869_, _00031_);
  nor _32587_ (_00033_, _00032_, _00030_);
  nor _32588_ (_28204_[13], _00033_, rst);
  nor _32589_ (_00034_, _24866_, _24529_);
  not _32590_ (_00035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _32591_ (_00036_, _24869_, _00035_);
  nor _32592_ (_00037_, _00036_, _00034_);
  nor _32593_ (_28204_[14], _00037_, rst);
  nor _32594_ (_00038_, _24866_, _28110_);
  not _32595_ (_00039_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _32596_ (_00040_, _24869_, _00039_);
  nor _32597_ (_00041_, _00040_, _00038_);
  nor _32598_ (_28205_[0], _00041_, rst);
  nor _32599_ (_00042_, _24866_, _28115_);
  not _32600_ (_00043_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _32601_ (_00044_, _24869_, _00043_);
  nor _32602_ (_00045_, _00044_, _00042_);
  nor _32603_ (_28205_[1], _00045_, rst);
  nor _32604_ (_00046_, _24866_, _28119_);
  not _32605_ (_00047_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _32606_ (_00048_, _24869_, _00047_);
  nor _32607_ (_00049_, _00048_, _00046_);
  nor _32608_ (_28205_[2], _00049_, rst);
  nor _32609_ (_00050_, _24866_, _28123_);
  not _32610_ (_00051_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _32611_ (_00052_, _24869_, _00051_);
  nor _32612_ (_00053_, _00052_, _00050_);
  nor _32613_ (_28205_[3], _00053_, rst);
  nor _32614_ (_00054_, _24866_, _28127_);
  not _32615_ (_00055_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _32616_ (_00056_, _24869_, _00055_);
  nor _32617_ (_00057_, _00056_, _00054_);
  nor _32618_ (_28205_[4], _00057_, rst);
  nor _32619_ (_00058_, _24866_, _28131_);
  not _32620_ (_00059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _32621_ (_00060_, _24869_, _00059_);
  nor _32622_ (_00061_, _00060_, _00058_);
  nor _32623_ (_28205_[5], _00061_, rst);
  nor _32624_ (_00062_, _24866_, _00001_);
  not _32625_ (_00063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _32626_ (_00064_, _24869_, _00063_);
  nor _32627_ (_00065_, _00064_, _00062_);
  nor _32628_ (_28205_[6], _00065_, rst);
  nor _32629_ (_00066_, _24866_, _00006_);
  not _32630_ (_00067_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _32631_ (_00068_, _24869_, _00067_);
  nor _32632_ (_00069_, _00068_, _00066_);
  nor _32633_ (_28205_[7], _00069_, rst);
  nor _32634_ (_00070_, _24866_, _00010_);
  not _32635_ (_00071_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _32636_ (_00072_, _24869_, _00071_);
  nor _32637_ (_00073_, _00072_, _00070_);
  nor _32638_ (_28205_[8], _00073_, rst);
  nor _32639_ (_00074_, _24866_, _00014_);
  not _32640_ (_00075_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _32641_ (_00076_, _24869_, _00075_);
  nor _32642_ (_00077_, _00076_, _00074_);
  nor _32643_ (_28205_[9], _00077_, rst);
  nor _32644_ (_00078_, _24866_, _00018_);
  not _32645_ (_00079_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _32646_ (_00080_, _24869_, _00079_);
  nor _32647_ (_00081_, _00080_, _00078_);
  nor _32648_ (_28205_[10], _00081_, rst);
  nor _32649_ (_00082_, _24866_, _00023_);
  not _32650_ (_00083_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _32651_ (_00084_, _24869_, _00083_);
  nor _32652_ (_00085_, _00084_, _00082_);
  nor _32653_ (_28205_[11], _00085_, rst);
  nor _32654_ (_00086_, _24866_, _00027_);
  not _32655_ (_00087_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _32656_ (_00088_, _24869_, _00087_);
  nor _32657_ (_00089_, _00088_, _00086_);
  nor _32658_ (_28205_[12], _00089_, rst);
  nor _32659_ (_00090_, _24866_, _00031_);
  not _32660_ (_00091_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _32661_ (_00092_, _24869_, _00091_);
  nor _32662_ (_00093_, _00092_, _00090_);
  nor _32663_ (_28205_[13], _00093_, rst);
  nor _32664_ (_00094_, _24866_, _00035_);
  not _32665_ (_00095_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _32666_ (_00096_, _24869_, _00095_);
  nor _32667_ (_00097_, _00096_, _00094_);
  nor _32668_ (_28205_[14], _00097_, rst);
  not _32669_ (_00098_, _25844_);
  nor _32670_ (_00099_, _00098_, \oc8051_top_1.oc8051_decoder1.state [1]);
  not _32671_ (_00100_, _00099_);
  nor _32672_ (_00101_, _25806_, _00100_);
  nor _32673_ (_00102_, _25588_, _25530_);
  nor _32674_ (_00103_, _00102_, _00101_);
  nor _32675_ (_00104_, _00103_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _32676_ (_00105_, _23909_, _23870_);
  nor _32677_ (_00106_, _00105_, _00104_);
  nor _32678_ (_28190_[2], _00106_, rst);
  nand _32679_ (_00107_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  nand _32680_ (_00108_, _25099_, _24074_);
  nand _32681_ (_04256_, _00108_, _00107_);
  nand _32682_ (_00109_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nand _32683_ (_00110_, _28096_, _24074_);
  nand _32684_ (_04364_, _00110_, _00109_);
  nand _32685_ (_00111_, _25203_, _24985_);
  nand _32686_ (_00112_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  nand _32687_ (_04506_, _00112_, _00111_);
  nor _32688_ (_00113_, _24976_, _24878_);
  not _32689_ (_00114_, _00113_);
  nor _32690_ (_00115_, _00114_, _25165_);
  nand _32691_ (_00116_, _00115_, _25150_);
  not _32692_ (_00117_, _00115_);
  nand _32693_ (_00118_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  nand _32694_ (_04561_, _00118_, _00116_);
  not _32695_ (_00119_, t2_i);
  nand _32696_ (_00120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _00119_);
  nor _32697_ (_05182_, _00120_, rst);
  nor _32698_ (_05204_, _00119_, rst);
  nor _32699_ (_00121_, _25045_, _24997_);
  not _32700_ (_00122_, _00121_);
  nor _32701_ (_00123_, _00122_, _24993_);
  nand _32702_ (_00124_, _00123_, _24789_);
  not _32703_ (_00125_, _00123_);
  nand _32704_ (_00126_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  nand _32705_ (_05881_, _00126_, _00124_);
  nand _32706_ (_00127_, _00123_, _25150_);
  nand _32707_ (_00128_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nand _32708_ (_05983_, _00128_, _00127_);
  nand _32709_ (_00129_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  nand _32710_ (_00130_, _25039_, _24074_);
  nand _32711_ (_06507_, _00130_, _00129_);
  not _32712_ (_00131_, _25626_);
  nor _32713_ (_00132_, _25049_, _00131_);
  not _32714_ (_00133_, _00132_);
  nor _32715_ (_00134_, _26410_, _23958_);
  nand _32716_ (_00135_, _00134_, _26402_);
  nor _32717_ (_00136_, _25631_, _23938_);
  not _32718_ (_00137_, _00136_);
  nor _32719_ (_00138_, _00137_, _00135_);
  not _32720_ (_00139_, _00138_);
  nor _32721_ (_00140_, _00139_, _00133_);
  not _32722_ (_00141_, _00140_);
  nor _32723_ (_00142_, _00141_, _24782_);
  not _32724_ (_00143_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor _32725_ (_00144_, _26410_, _25721_);
  not _32726_ (_00145_, _00144_);
  nor _32727_ (_00146_, _00145_, _24051_);
  not _32728_ (_00147_, _00146_);
  nor _32729_ (_00148_, _00137_, _00147_);
  not _32730_ (_00149_, _00148_);
  nor _32731_ (_00150_, _00149_, _00133_);
  nand _32732_ (_00151_, _00150_, _00143_);
  not _32733_ (_00152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _32734_ (_00153_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  not _32735_ (_00154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor _32736_ (_00155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _32737_ (_00156_, _00155_, _00154_);
  nor _32738_ (_00157_, _00156_, _00153_);
  not _32739_ (_00158_, _00157_);
  nor _32740_ (_00159_, _00158_, _00152_);
  nor _32741_ (_00160_, _00150_, _00159_);
  not _32742_ (_00161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  not _32743_ (_00162_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  not _32744_ (_00163_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  nand _32745_ (_00164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _32746_ (_00165_, _00164_);
  not _32747_ (_00166_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _32748_ (_00167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _00166_);
  nor _32749_ (_00168_, _00167_, _00165_);
  nor _32750_ (_00169_, _00168_, _00163_);
  not _32751_ (_00170_, _00169_);
  not _32752_ (_00171_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  not _32753_ (_00172_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  not _32754_ (_00173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _32755_ (_00174_, _00173_, _00172_);
  nand _32756_ (_00175_, _00174_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  not _32757_ (_00176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  not _32758_ (_00177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor _32759_ (_00178_, _00177_, _00176_);
  not _32760_ (_00179_, _00178_);
  not _32761_ (_00180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  not _32762_ (_00181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _32763_ (_00182_, _00181_, _00180_);
  not _32764_ (_00183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  not _32765_ (_00184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _32766_ (_00185_, _00184_, _00183_);
  nand _32767_ (_00186_, _00185_, _00182_);
  nor _32768_ (_00187_, _00186_, _00179_);
  not _32769_ (_00188_, _00187_);
  nor _32770_ (_00189_, _00188_, _00175_);
  not _32771_ (_00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  not _32772_ (_00191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _32773_ (_00192_, _00191_, _00190_);
  nand _32774_ (_00193_, _00192_, _00189_);
  nor _32775_ (_00194_, _00193_, _00171_);
  not _32776_ (_00195_, _00194_);
  nor _32777_ (_00196_, _00195_, _00170_);
  not _32778_ (_00197_, _00196_);
  nor _32779_ (_00198_, _00197_, _00162_);
  not _32780_ (_00199_, _00198_);
  nor _32781_ (_00200_, _00199_, _00161_);
  nand _32782_ (_00201_, _00200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand _32783_ (_00202_, _00201_, _00143_);
  not _32784_ (_00203_, _00155_);
  nor _32785_ (_00204_, _00203_, _00154_);
  not _32786_ (_00205_, _00204_);
  nand _32787_ (_00206_, _00205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _32788_ (_00207_, _00206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor _32789_ (_00208_, _00207_, _00201_);
  nor _32790_ (_00209_, _00208_, _00157_);
  nand _32791_ (_00210_, _00209_, _00202_);
  nand _32792_ (_00211_, _00210_, _00160_);
  nand _32793_ (_00212_, _00211_, _00151_);
  nand _32794_ (_00213_, _00212_, _00141_);
  nand _32795_ (_00214_, _00213_, _26487_);
  nor _32796_ (_06567_, _00214_, _00142_);
  not _32797_ (_00215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  not _32798_ (_00216_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nand _32799_ (_00217_, _00216_, _00215_);
  nor _32800_ (_00218_, _23978_, _23938_);
  not _32801_ (_00219_, _00218_);
  nor _32802_ (_00220_, _00219_, _26258_);
  nor _32803_ (_00221_, _26245_, _23915_);
  nand _32804_ (_00222_, _00221_, _00220_);
  not _32805_ (_00223_, _00222_);
  nor _32806_ (_00224_, _00223_, _00217_);
  nand _32807_ (_00225_, _26135_, _24716_);
  not _32808_ (_00226_, _00225_);
  not _32809_ (_00227_, _26135_);
  nand _32810_ (_00228_, _00227_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _32811_ (_00229_, _00228_, _00223_);
  nor _32812_ (_00230_, _00229_, _00226_);
  nor _32813_ (_00231_, _00230_, _00224_);
  nor _32814_ (_00232_, _25723_, _23938_);
  not _32815_ (_00233_, _00232_);
  nor _32816_ (_00234_, _25631_, _00233_);
  not _32817_ (_00235_, _00234_);
  nor _32818_ (_00236_, _00235_, _00133_);
  nor _32819_ (_00237_, _00236_, _00231_);
  nand _32820_ (_00238_, _00236_, _25625_);
  nand _32821_ (_00239_, _00238_, _26487_);
  nor _32822_ (_06684_, _00239_, _00237_);
  nor _32823_ (_00240_, _00150_, _00140_);
  not _32824_ (_00241_, _00240_);
  not _32825_ (_00242_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _32826_ (_00243_, _00242_, _00143_);
  nand _32827_ (_00244_, _00243_, _00200_);
  not _32828_ (_00245_, _00244_);
  nor _32829_ (_00246_, _00157_, _00203_);
  nand _32830_ (_00247_, _00246_, _00245_);
  nor _32831_ (_00248_, _00247_, _00241_);
  nor _32832_ (_00249_, _00240_, _00216_);
  nor _32833_ (_00250_, _00249_, _00248_);
  nor _32834_ (_06708_, _00250_, rst);
  not _32835_ (_00251_, t2ex_i);
  nor _32836_ (_06792_, _00251_, rst);
  nand _32837_ (_00252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _26487_);
  nor _32838_ (_06839_, _00252_, t2ex_i);
  nor _32839_ (_00253_, _00170_, _00155_);
  nand _32840_ (_00254_, _00253_, _00240_);
  nor _32841_ (_00255_, _00162_, _00161_);
  nand _32842_ (_00256_, _00243_, _00255_);
  nor _32843_ (_00257_, _00256_, _00195_);
  nor _32844_ (_00258_, _00257_, _00254_);
  not _32845_ (_00259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  nand _32846_ (_00260_, _00254_, _00259_);
  nand _32847_ (_00261_, _00260_, _26487_);
  nor _32848_ (_06921_, _00261_, _00258_);
  nor _32849_ (_00262_, _23996_, _23958_);
  nand _32850_ (_00263_, _00262_, _24051_);
  nor _32851_ (_00264_, _00263_, _23938_);
  not _32852_ (_00265_, _00264_);
  nor _32853_ (_00266_, _00265_, _25631_);
  not _32854_ (_00267_, _00266_);
  nor _32855_ (_00268_, _00267_, _00133_);
  not _32856_ (_00269_, _00268_);
  nor _32857_ (_00270_, _00269_, _24782_);
  nor _32858_ (_00271_, _00205_, _00153_);
  not _32859_ (_00272_, _00271_);
  nor _32860_ (_00273_, _23996_, _25721_);
  not _32861_ (_00274_, _00273_);
  nor _32862_ (_00275_, _00274_, _26402_);
  not _32863_ (_00276_, _00275_);
  nor _32864_ (_00277_, _00137_, _00276_);
  not _32865_ (_00278_, _00277_);
  nor _32866_ (_00279_, _00278_, _00133_);
  nor _32867_ (_00280_, _00279_, _00272_);
  nor _32868_ (_00281_, _00280_, _00152_);
  not _32869_ (_00282_, _00280_);
  nor _32870_ (_00283_, _00282_, _00143_);
  nor _32871_ (_00284_, _00283_, _00281_);
  nand _32872_ (_00285_, _00269_, _00284_);
  nand _32873_ (_00286_, _00285_, _26487_);
  nor _32874_ (_06946_, _00286_, _00270_);
  not _32875_ (_00287_, _00279_);
  nor _32876_ (_00288_, _00287_, _24782_);
  not _32877_ (_00289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _32878_ (_00290_, _00271_, _00289_);
  nor _32879_ (_00291_, _00272_, _00177_);
  nor _32880_ (_00292_, _00291_, _00290_);
  nand _32881_ (_00293_, _00292_, _00287_);
  nand _32882_ (_00294_, _00293_, _00269_);
  nor _32883_ (_00295_, _00294_, _00288_);
  nor _32884_ (_00296_, _00137_, _00263_);
  nand _32885_ (_00297_, _00296_, _00132_);
  nor _32886_ (_00298_, _00297_, _00289_);
  nor _32887_ (_00299_, _00298_, _00295_);
  nor _32888_ (_06973_, _00299_, rst);
  nand _32889_ (_00300_, _28099_, _24830_);
  nand _32890_ (_00301_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  nand _32891_ (_07035_, _00301_, _00300_);
  not _32892_ (_00302_, _00150_);
  nor _32893_ (_00303_, _00302_, _24782_);
  not _32894_ (_00304_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _32895_ (_00305_, _00184_, _00176_);
  nand _32896_ (_00306_, _00305_, _00182_);
  nor _32897_ (_00307_, _00306_, _00172_);
  nand _32898_ (_00308_, _00307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _32899_ (_00309_, _00308_, _00304_);
  not _32900_ (_00310_, _00309_);
  nor _32901_ (_00311_, _00310_, _00170_);
  nor _32902_ (_00312_, _00311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor _32903_ (_00313_, _00310_, _00177_);
  not _32904_ (_00314_, _00313_);
  nor _32905_ (_00315_, _00314_, _00170_);
  nor _32906_ (_00316_, _00315_, _00312_);
  nand _32907_ (_00317_, _00205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _32908_ (_00318_, _00317_, _00244_);
  nor _32909_ (_00319_, _00318_, _00316_);
  nor _32910_ (_00320_, _00319_, _00157_);
  nor _32911_ (_00321_, _00158_, _00289_);
  nor _32912_ (_00322_, _00321_, _00320_);
  nand _32913_ (_00323_, _00322_, _00302_);
  nand _32914_ (_00324_, _00323_, _00141_);
  nor _32915_ (_00325_, _00324_, _00303_);
  nor _32916_ (_00326_, _00141_, _00177_);
  nor _32917_ (_00327_, _00326_, _00325_);
  nor _32918_ (_07103_, _00327_, rst);
  nand _32919_ (_00328_, _25000_, _24830_);
  nand _32920_ (_00329_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nand _32921_ (_08762_, _00329_, _00328_);
  nor _32922_ (_00330_, _24978_, _24073_);
  not _32923_ (_00331_, _00330_);
  nand _32924_ (_00332_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nand _32925_ (_00333_, _00330_, _28096_);
  nand _32926_ (_08986_, _00333_, _00332_);
  nand _32927_ (_00334_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  nand _32928_ (_00335_, _00330_, _25039_);
  nand _32929_ (_09316_, _00335_, _00334_);
  nand _32930_ (_00336_, _00123_, _28096_);
  nand _32931_ (_00337_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  nand _32932_ (_09479_, _00337_, _00336_);
  nand _32933_ (_00338_, _00123_, _25099_);
  nand _32934_ (_00339_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  nand _32935_ (_09544_, _00339_, _00338_);
  nand _32936_ (_00340_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  nand _32937_ (_00341_, _00330_, _25203_);
  nand _32938_ (_09650_, _00341_, _00340_);
  nand _32939_ (_00342_, _00123_, _24927_);
  nand _32940_ (_00343_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nand _32941_ (_10271_, _00343_, _00342_);
  nand _32942_ (_00344_, _00123_, _25039_);
  nand _32943_ (_00345_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nand _32944_ (_10448_, _00345_, _00344_);
  nand _32945_ (_00346_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nand _32946_ (_00347_, _00330_, _25150_);
  nand _32947_ (_10502_, _00347_, _00346_);
  nand _32948_ (_00348_, _28081_, _24830_);
  nand _32949_ (_00349_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nand _32950_ (_10558_, _00349_, _00348_);
  nand _32951_ (_00350_, _00115_, _24927_);
  nand _32952_ (_00351_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  nand _32953_ (_10612_, _00351_, _00350_);
  nand _32954_ (_00352_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  nand _32955_ (_00353_, _00330_, _24789_);
  nand _32956_ (_10719_, _00353_, _00352_);
  nand _32957_ (_00354_, _28059_, _25150_);
  nand _32958_ (_00355_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  nand _32959_ (_10987_, _00355_, _00354_);
  nor _32960_ (_00356_, _25047_, _24993_);
  nand _32961_ (_00357_, _00356_, _24927_);
  not _32962_ (_00358_, _00356_);
  nand _32963_ (_00359_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  nand _32964_ (_11178_, _00359_, _00357_);
  nor _32965_ (_28182_[4], _27733_, rst);
  nor _32966_ (_00360_, _24999_, _24073_);
  not _32967_ (_00361_, _00360_);
  nand _32968_ (_00362_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  nand _32969_ (_00363_, _00360_, _28096_);
  nand _32970_ (_11748_, _00363_, _00362_);
  nand _32971_ (_00364_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nand _32972_ (_00365_, _00360_, _25039_);
  nand _32973_ (_11816_, _00365_, _00364_);
  nand _32974_ (_00366_, _00356_, _24789_);
  nand _32975_ (_00367_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  nand _32976_ (_11868_, _00367_, _00366_);
  nand _32977_ (_00368_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  nand _32978_ (_00369_, _00360_, _25203_);
  nand _32979_ (_12042_, _00369_, _00368_);
  nand _32980_ (_00370_, _00356_, _25150_);
  nand _32981_ (_00371_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  nand _32982_ (_12057_, _00371_, _00370_);
  nor _32983_ (_00372_, _00137_, _25723_);
  not _32984_ (_00373_, _00372_);
  nor _32985_ (_00374_, _00373_, _00133_);
  not _32986_ (_00375_, _00374_);
  nor _32987_ (_00376_, _00144_, _24051_);
  nor _32988_ (_00377_, _00376_, _25722_);
  nand _32989_ (_00378_, _00377_, _00223_);
  nand _32990_ (_00379_, _00378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _32991_ (_00380_, _00379_, _00375_);
  nand _32992_ (_00381_, _00146_, _24716_);
  not _32993_ (_00382_, _00381_);
  not _32994_ (_00383_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor _32995_ (_00384_, _00144_, _26402_);
  not _32996_ (_00385_, _00384_);
  nor _32997_ (_00386_, _00385_, _00383_);
  nor _32998_ (_00387_, _00386_, _00382_);
  nor _32999_ (_00388_, _00387_, _00222_);
  nor _33000_ (_00389_, _00388_, _00380_);
  nand _33001_ (_00390_, _00236_, _25029_);
  nand _33002_ (_00391_, _00390_, _26487_);
  nor _33003_ (_12253_, _00391_, _00389_);
  nor _33004_ (_00392_, _24997_, _24878_);
  not _33005_ (_00393_, _00392_);
  nor _33006_ (_00394_, _00393_, _28057_);
  nand _33007_ (_00395_, _00394_, _25150_);
  not _33008_ (_00396_, _00394_);
  nand _33009_ (_00397_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  nand _33010_ (_12364_, _00397_, _00395_);
  nand _33011_ (_00398_, _00356_, _24830_);
  nand _33012_ (_00399_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  nand _33013_ (_12491_, _00399_, _00398_);
  nand _33014_ (_00400_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  nand _33015_ (_00401_, _00360_, _24789_);
  nand _33016_ (_12659_, _00401_, _00400_);
  nand _33017_ (_00402_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  nand _33018_ (_00403_, _00360_, _25150_);
  nand _33019_ (_12675_, _00403_, _00402_);
  nand _33020_ (_00404_, _00356_, _28096_);
  nand _33021_ (_00405_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nand _33022_ (_12718_, _00405_, _00404_);
  nand _33023_ (_00406_, _00356_, _25203_);
  nand _33024_ (_00407_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  nand _33025_ (_12867_, _00407_, _00406_);
  nor _33026_ (_00408_, _25057_, _24073_);
  not _33027_ (_00409_, _00408_);
  nand _33028_ (_00410_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nand _33029_ (_00411_, _00408_, _25203_);
  nand _33030_ (_13083_, _00411_, _00410_);
  nand _33031_ (_00412_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  nand _33032_ (_00413_, _00408_, _24927_);
  nand _33033_ (_13257_, _00413_, _00412_);
  nor _33034_ (_00414_, _25045_, _24001_);
  not _33035_ (_00415_, _00414_);
  nor _33036_ (_00416_, _00415_, _24993_);
  nand _33037_ (_00417_, _00416_, _25039_);
  not _33038_ (_00418_, _00416_);
  nand _33039_ (_00419_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  nand _33040_ (_13278_, _00419_, _00417_);
  nand _33041_ (_00420_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  nand _33042_ (_00421_, _00408_, _25039_);
  nand _33043_ (_13359_, _00421_, _00420_);
  not _33044_ (_00422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor _33045_ (_00423_, _00385_, _00422_);
  nor _33046_ (_00424_, _00423_, _00382_);
  nor _33047_ (_00425_, _23979_, _23938_);
  not _33048_ (_00426_, _00425_);
  nor _33049_ (_00427_, _24035_, _24069_);
  nand _33050_ (_00428_, _00427_, _00221_);
  nor _33051_ (_00429_, _00428_, _00426_);
  not _33052_ (_00430_, _00429_);
  nor _33053_ (_00431_, _00430_, _00424_);
  nand _33054_ (_00432_, _00429_, _00377_);
  nand _33055_ (_00433_, _00432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor _33056_ (_00434_, _00227_, _25726_);
  nor _33057_ (_00435_, _24035_, _23979_);
  not _33058_ (_00436_, _00435_);
  nor _33059_ (_00437_, _00436_, _24071_);
  nand _33060_ (_00438_, _00437_, _00434_);
  nand _33061_ (_00439_, _00438_, _00433_);
  nor _33062_ (_00440_, _00439_, _00431_);
  not _33063_ (_00441_, _00438_);
  nand _33064_ (_00442_, _00441_, _25029_);
  nand _33065_ (_00443_, _00442_, _26487_);
  nor _33066_ (_13590_, _00443_, _00440_);
  not _33067_ (_00444_, _00263_);
  nand _33068_ (_00445_, _00429_, _00444_);
  nor _33069_ (_00446_, _00445_, _24716_);
  not _33070_ (_00447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand _33071_ (_00448_, _00445_, _00447_);
  nand _33072_ (_00449_, _00448_, _00438_);
  nor _33073_ (_00450_, _00449_, _00446_);
  nor _33074_ (_00451_, _00438_, _25195_);
  nor _33075_ (_00452_, _00451_, _00450_);
  nor _33076_ (_13611_, _00452_, rst);
  nand _33077_ (_00453_, _00416_, _25150_);
  nand _33078_ (_00454_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nand _33079_ (_13632_, _00454_, _00453_);
  nor _33080_ (_00455_, _00430_, _00276_);
  not _33081_ (_00456_, _00455_);
  nor _33082_ (_00457_, _00456_, _24716_);
  nor _33083_ (_00458_, _00455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _33084_ (_00459_, _00458_, _00457_);
  nor _33085_ (_00460_, _00459_, _00441_);
  nand _33086_ (_00461_, _00441_, _25703_);
  nand _33087_ (_00462_, _00461_, _26487_);
  nor _33088_ (_13653_, _00462_, _00460_);
  nor _33089_ (_00463_, _00430_, _24842_);
  not _33090_ (_00464_, _00463_);
  nor _33091_ (_00465_, _00464_, _24716_);
  nor _33092_ (_00466_, _00463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _33093_ (_00467_, _00466_, _00465_);
  nor _33094_ (_00468_, _00467_, _00441_);
  nand _33095_ (_00469_, _00441_, _25088_);
  nand _33096_ (_00470_, _00469_, _26487_);
  nor _33097_ (_13674_, _00470_, _00468_);
  nand _33098_ (_00471_, _00429_, _25722_);
  nor _33099_ (_00472_, _00471_, _24716_);
  not _33100_ (_00473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand _33101_ (_00474_, _00471_, _00473_);
  nand _33102_ (_00475_, _00474_, _00438_);
  nor _33103_ (_00476_, _00475_, _00472_);
  nor _33104_ (_00477_, _00438_, _24820_);
  nor _33105_ (_00478_, _00477_, _00476_);
  nor _33106_ (_13695_, _00478_, rst);
  nor _33107_ (_00479_, _24978_, _24993_);
  nand _33108_ (_00480_, _00479_, _25150_);
  not _33109_ (_00481_, _00479_);
  nand _33110_ (_00482_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nand _33111_ (_13886_, _00482_, _00480_);
  nand _33112_ (_00483_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  nand _33113_ (_00484_, _00408_, _24789_);
  nand _33114_ (_13906_, _00484_, _00483_);
  nand _33115_ (_00485_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  nand _33116_ (_00486_, _00360_, _24830_);
  nand _33117_ (_13987_, _00486_, _00485_);
  nand _33118_ (_00487_, _00416_, _24830_);
  nand _33119_ (_00488_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nand _33120_ (_14118_, _00488_, _00487_);
  nand _33121_ (_00489_, _00444_, _24716_);
  not _33122_ (_00490_, _00489_);
  nand _33123_ (_00491_, _24051_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor _33124_ (_00492_, _00491_, _00262_);
  nor _33125_ (_00493_, _00492_, _00490_);
  nor _33126_ (_00494_, _00428_, _00219_);
  not _33127_ (_00495_, _00494_);
  nor _33128_ (_00496_, _00495_, _00493_);
  nor _33129_ (_00497_, _00495_, _26402_);
  not _33130_ (_00498_, _00497_);
  nand _33131_ (_00499_, _00498_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor _33132_ (_00500_, _26231_, _24071_);
  not _33133_ (_00501_, _00500_);
  nor _33134_ (_00502_, _00501_, _00373_);
  not _33135_ (_00503_, _00502_);
  nand _33136_ (_00504_, _00503_, _00499_);
  nor _33137_ (_00505_, _00504_, _00496_);
  nor _33138_ (_00506_, _00501_, _00235_);
  nand _33139_ (_00507_, _00506_, _25195_);
  nand _33140_ (_00508_, _00507_, _26487_);
  nor _33141_ (_14199_, _00508_, _00505_);
  not _33142_ (_00509_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nand _33143_ (_00510_, _00494_, _00275_);
  nand _33144_ (_00511_, _00510_, _00509_);
  nand _33145_ (_00512_, _00511_, _00503_);
  nor _33146_ (_00513_, _00510_, _24716_);
  nor _33147_ (_00514_, _00513_, _00512_);
  nor _33148_ (_00515_, _00503_, _25703_);
  nor _33149_ (_00516_, _00515_, _00514_);
  nor _33150_ (_14220_, _00516_, rst);
  not _33151_ (_00517_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nand _33152_ (_00518_, _00494_, _24840_);
  nand _33153_ (_00519_, _00518_, _00517_);
  nand _33154_ (_00520_, _00519_, _00503_);
  nor _33155_ (_00521_, _00518_, _24716_);
  nor _33156_ (_00522_, _00521_, _00520_);
  nor _33157_ (_00523_, _00503_, _25088_);
  nor _33158_ (_00524_, _00523_, _00522_);
  nor _33159_ (_14241_, _00524_, rst);
  nor _33160_ (_00525_, _00498_, _00145_);
  not _33161_ (_00526_, _00525_);
  nor _33162_ (_00527_, _00526_, _24716_);
  nor _33163_ (_00528_, _00525_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nor _33164_ (_00529_, _00528_, _00527_);
  nor _33165_ (_00530_, _00529_, _00502_);
  nand _33166_ (_00531_, _00502_, _24820_);
  nand _33167_ (_00532_, _00531_, _26487_);
  nor _33168_ (_14262_, _00532_, _00530_);
  nand _33169_ (_00533_, _00416_, _28096_);
  nand _33170_ (_00534_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  nand _33171_ (_14393_, _00534_, _00533_);
  not _33172_ (_00535_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _33173_ (_00536_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _33174_ (_00537_, _00536_);
  nor _33175_ (_00538_, _00537_, _00535_);
  not _33176_ (_00539_, _00538_);
  not _33177_ (_00540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _33178_ (_00541_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  nor _33179_ (_00542_, _00541_, _00535_);
  not _33180_ (_00543_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not _33181_ (_00544_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  nor _33182_ (_00545_, _00544_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _33183_ (_00546_, _00545_, _00543_);
  not _33184_ (_00547_, _00546_);
  nor _33185_ (_00548_, _00547_, _00542_);
  nor _33186_ (_00549_, _00548_, _00540_);
  not _33187_ (_00550_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  not _33188_ (_00551_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nor _33189_ (_00552_, _00551_, _00550_);
  not _33190_ (_00553_, _00552_);
  nor _33191_ (_00554_, _00553_, _00473_);
  not _33192_ (_00555_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  not _33193_ (_00556_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nor _33194_ (_00557_, _00517_, _00556_);
  not _33195_ (_00558_, _00557_);
  nor _33196_ (_00559_, _00558_, _00555_);
  not _33197_ (_00561_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not _33198_ (_00562_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nor _33199_ (_00563_, _00562_, _00509_);
  not _33200_ (_00564_, _00563_);
  nor _33201_ (_00565_, _00564_, _00561_);
  nor _33202_ (_00566_, _00565_, _00559_);
  not _33203_ (_00567_, _00566_);
  nor _33204_ (_00568_, _00567_, _00554_);
  not _33205_ (_00570_, _00568_);
  not _33206_ (_00571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _33207_ (_00572_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor _33208_ (_00573_, _00572_, _00571_);
  not _33209_ (_00575_, _00573_);
  nor _33210_ (_00576_, _00575_, _00422_);
  not _33211_ (_00577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _33212_ (_00578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _33213_ (_00579_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _33214_ (_00580_, _00579_, _00578_);
  not _33215_ (_00581_, _00580_);
  nor _33216_ (_00582_, _00581_, _00577_);
  nor _33217_ (_00583_, _00582_, _00576_);
  not _33218_ (_00584_, _00583_);
  nand _33219_ (_00585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor _33220_ (_00586_, _00585_, _00447_);
  nor _33221_ (_00587_, _00586_, _00584_);
  not _33222_ (_00588_, _00587_);
  nor _33223_ (_00589_, _00588_, _00570_);
  nor _33224_ (_00590_, _00589_, _00549_);
  not _33225_ (_00591_, _00590_);
  nor _33226_ (_00592_, _00591_, _00539_);
  nor _33227_ (_00593_, _00543_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _33228_ (_00594_, _00593_);
  nor _33229_ (_00595_, _00575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor _33230_ (_00596_, _00581_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  nor _33231_ (_00597_, _00596_, _00595_);
  not _33232_ (_00598_, _00597_);
  nor _33233_ (_00599_, _00585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor _33234_ (_00600_, _00599_, _00598_);
  nor _33235_ (_00601_, _00600_, _00594_);
  nor _33236_ (_00602_, _00553_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _33237_ (_00603_, _00602_);
  nor _33238_ (_00604_, _00558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  not _33239_ (_00606_, _00604_);
  nand _33240_ (_00607_, _00606_, _00603_);
  nor _33241_ (_00608_, _00564_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _33242_ (_00609_, _00608_, _00607_);
  nor _33243_ (_00610_, _00609_, _00594_);
  nor _33244_ (_00611_, _00610_, _00601_);
  nor _33245_ (_00612_, _00611_, _00539_);
  nor _33246_ (_00613_, _00612_, _00544_);
  nor _33247_ (_00614_, _00613_, _00592_);
  nor _33248_ (_14554_, _00614_, rst);
  not _33249_ (_00615_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nor _33250_ (_00616_, _24060_, _24069_);
  not _33251_ (_00617_, _00616_);
  nand _33252_ (_00618_, _00221_, _00218_);
  nor _33253_ (_00619_, _00618_, _00617_);
  nand _33254_ (_00620_, _00619_, _25722_);
  nand _33255_ (_00621_, _00620_, _00615_);
  nand _33256_ (_00622_, _00372_, _25628_);
  nand _33257_ (_00623_, _00622_, _00621_);
  nor _33258_ (_00624_, _00620_, _24716_);
  nor _33259_ (_00625_, _00624_, _00623_);
  nor _33260_ (_00626_, _00622_, _24820_);
  nor _33261_ (_00627_, _00626_, _00625_);
  nor _33262_ (_14744_, _00627_, rst);
  nor _33263_ (_00628_, _24878_, _24001_);
  not _33264_ (_00629_, _00628_);
  nor _33265_ (_00630_, _24991_, _24068_);
  not _33266_ (_00631_, _00630_);
  nor _33267_ (_00632_, _00631_, _00629_);
  nand _33268_ (_00633_, _00632_, _25099_);
  not _33269_ (_00634_, _00632_);
  nand _33270_ (_00635_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  nand _33271_ (_14775_, _00635_, _00633_);
  nor _33272_ (_00636_, _28080_, _24073_);
  not _33273_ (_00637_, _00636_);
  nand _33274_ (_00638_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  nand _33275_ (_00639_, _00636_, _24927_);
  nand _33276_ (_14926_, _00639_, _00638_);
  not _33277_ (_00640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _33278_ (_00641_, _00611_);
  nor _33279_ (_00642_, _00641_, _00590_);
  nor _33280_ (_00643_, _00642_, _00537_);
  nor _33281_ (_00644_, _00643_, _00640_);
  not _33282_ (_00645_, _00576_);
  nor _33283_ (_00646_, _00645_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _33284_ (_00647_, _00646_, _00586_);
  nand _33285_ (_00648_, _00582_, _00535_);
  nand _33286_ (_00649_, _00648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nand _33287_ (_00650_, _00649_, _00647_);
  nor _33288_ (_00651_, _00640_, _00535_);
  not _33289_ (_00652_, _00651_);
  nand _33290_ (_00653_, _00652_, _00586_);
  nand _33291_ (_00654_, _00653_, _00650_);
  nor _33292_ (_00655_, _00654_, _00565_);
  not _33293_ (_00656_, _00565_);
  nor _33294_ (_00657_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00535_);
  nor _33295_ (_00658_, _00657_, _00656_);
  nor _33296_ (_00659_, _00658_, _00655_);
  nor _33297_ (_00660_, _00659_, _00559_);
  not _33298_ (_00661_, _00554_);
  nand _33299_ (_00662_, _00651_, _00559_);
  nand _33300_ (_00663_, _00662_, _00661_);
  nor _33301_ (_00664_, _00663_, _00660_);
  nand _33302_ (_00665_, _00657_, _00554_);
  nand _33303_ (_00666_, _00665_, _00590_);
  nor _33304_ (_00667_, _00666_, _00664_);
  nor _33305_ (_00668_, _00611_, _00590_);
  not _33306_ (_00669_, _00668_);
  nor _33307_ (_00670_, _00657_, _00603_);
  not _33308_ (_00671_, _00595_);
  nor _33309_ (_00672_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _33310_ (_00674_, _00672_, _00599_);
  not _33311_ (_00675_, _00596_);
  nor _33312_ (_00676_, _00675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _33313_ (_00677_, _00676_);
  nand _33314_ (_00678_, _00677_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nand _33315_ (_00679_, _00678_, _00674_);
  nand _33316_ (_00680_, _00652_, _00599_);
  nand _33317_ (_00681_, _00680_, _00679_);
  nor _33318_ (_00682_, _00681_, _00608_);
  not _33319_ (_00683_, _00608_);
  nor _33320_ (_00684_, _00657_, _00683_);
  nor _33321_ (_00685_, _00684_, _00682_);
  nor _33322_ (_00686_, _00685_, _00604_);
  nor _33323_ (_00687_, _00652_, _00606_);
  nor _33324_ (_00688_, _00687_, _00686_);
  nor _33325_ (_00689_, _00688_, _00602_);
  nor _33326_ (_00690_, _00689_, _00670_);
  nor _33327_ (_00691_, _00690_, _00669_);
  nor _33328_ (_00692_, _00691_, _00667_);
  nor _33329_ (_00693_, _00692_, _00537_);
  nor _33330_ (_00694_, _00693_, _00644_);
  nor _33331_ (_14987_, _00694_, rst);
  nor _33332_ (_00695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00535_);
  nor _33333_ (_00696_, _00695_, _00602_);
  nor _33334_ (_00697_, _00696_, _00609_);
  not _33335_ (_00698_, _00599_);
  not _33336_ (_00699_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nor _33337_ (_00701_, _00699_, _00535_);
  not _33338_ (_00702_, _00701_);
  nor _33339_ (_00703_, _00702_, _00698_);
  nor _33340_ (_00704_, _00608_, _00604_);
  nand _33341_ (_00705_, _00677_, _00699_);
  nand _33342_ (_00706_, _00705_, _00674_);
  nand _33343_ (_00707_, _00706_, _00704_);
  nor _33344_ (_00708_, _00707_, _00703_);
  nor _33345_ (_00709_, _00708_, _00697_);
  nand _33346_ (_00710_, _00701_, _00602_);
  nand _33347_ (_00711_, _00710_, _00641_);
  nor _33348_ (_00712_, _00711_, _00709_);
  nor _33349_ (_00713_, _00641_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nor _33350_ (_00714_, _00713_, _00712_);
  nand _33351_ (_00715_, _00714_, _00591_);
  nand _33352_ (_00716_, _00701_, _00554_);
  not _33353_ (_00717_, _00695_);
  nor _33354_ (_00718_, _00717_, _00566_);
  nor _33355_ (_00719_, _00718_, _00554_);
  nand _33356_ (_00720_, _00648_, _00699_);
  nand _33357_ (_00721_, _00720_, _00647_);
  not _33358_ (_00722_, _00586_);
  nor _33359_ (_00723_, _00702_, _00722_);
  nor _33360_ (_00724_, _00723_, _00567_);
  nand _33361_ (_00725_, _00724_, _00721_);
  nand _33362_ (_00726_, _00725_, _00719_);
  nand _33363_ (_00727_, _00726_, _00716_);
  nand _33364_ (_00728_, _00727_, _00590_);
  nand _33365_ (_00729_, _00728_, _00715_);
  nor _33366_ (_00730_, _00729_, _00537_);
  nand _33367_ (_00731_, _00537_, _00699_);
  nand _33368_ (_00732_, _00731_, _26487_);
  nor _33369_ (_15098_, _00732_, _00730_);
  nand _33370_ (_00733_, _28096_, _28063_);
  nand _33371_ (_00734_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  nand _33372_ (_15309_, _00734_, _00733_);
  nor _33373_ (_00735_, _00631_, _00114_);
  nand _33374_ (_00736_, _00735_, _24789_);
  not _33375_ (_00737_, _00735_);
  nand _33376_ (_00738_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  nand _33377_ (_15340_, _00738_, _00736_);
  not _33378_ (_00739_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nand _33379_ (_00740_, _00537_, _00739_);
  nand _33380_ (_00741_, _00740_, _26487_);
  nor _33381_ (_00742_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _33382_ (_00743_, _00742_, _00586_);
  not _33383_ (_00744_, _00582_);
  nor _33384_ (_00745_, _00744_, _00535_);
  nor _33385_ (_00746_, _00745_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _33386_ (_00747_, _00645_, _00535_);
  nor _33387_ (_00749_, _00747_, _00586_);
  not _33388_ (_00750_, _00749_);
  nor _33389_ (_00751_, _00750_, _00746_);
  nor _33390_ (_00752_, _00751_, _00567_);
  nand _33391_ (_00753_, _00752_, _00743_);
  nor _33392_ (_00754_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _33393_ (_00755_, _00754_);
  nor _33394_ (_00756_, _00755_, _00566_);
  nor _33395_ (_00757_, _00756_, _00554_);
  nand _33396_ (_00758_, _00757_, _00753_);
  nand _33397_ (_00759_, _00742_, _00554_);
  nand _33398_ (_00760_, _00759_, _00758_);
  nor _33399_ (_00761_, _00760_, _00591_);
  nor _33400_ (_00762_, _00671_, _00535_);
  nor _33401_ (_00763_, _00762_, _00599_);
  not _33402_ (_00764_, _00763_);
  nor _33403_ (_00765_, _00675_, _00535_);
  nor _33404_ (_00766_, _00765_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _33405_ (_00767_, _00766_, _00764_);
  nand _33406_ (_00768_, _00742_, _00599_);
  nand _33407_ (_00769_, _00768_, _00704_);
  nor _33408_ (_00770_, _00769_, _00767_);
  nor _33409_ (_00771_, _00754_, _00602_);
  nor _33410_ (_00772_, _00771_, _00609_);
  nor _33411_ (_00773_, _00772_, _00770_);
  nand _33412_ (_00774_, _00742_, _00602_);
  nand _33413_ (_00775_, _00774_, _00641_);
  nor _33414_ (_00776_, _00775_, _00773_);
  nor _33415_ (_00777_, _00641_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _33416_ (_00778_, _00777_, _00776_);
  nor _33417_ (_00779_, _00778_, _00590_);
  nor _33418_ (_00780_, _00779_, _00761_);
  nor _33419_ (_00781_, _00780_, _00537_);
  nor _33420_ (_15361_, _00781_, _00741_);
  not _33421_ (_00782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor _33422_ (_00783_, _00643_, _00782_);
  nor _33423_ (_00784_, _00722_, _00565_);
  nor _33424_ (_00785_, _00784_, _00559_);
  nor _33425_ (_00786_, _00782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _33426_ (_00787_, _00786_, _00785_);
  nor _33427_ (_00788_, _00745_, _00782_);
  nand _33428_ (_00789_, _00749_, _00566_);
  nor _33429_ (_00790_, _00789_, _00788_);
  nor _33430_ (_00791_, _00790_, _00787_);
  nor _33431_ (_00792_, _00791_, _00554_);
  nor _33432_ (_00793_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _33433_ (_00794_, _00559_);
  nand _33434_ (_00795_, _00565_, _00794_);
  nand _33435_ (_00796_, _00795_, _00661_);
  nand _33436_ (_00797_, _00796_, _00793_);
  nand _33437_ (_00798_, _00797_, _00590_);
  nor _33438_ (_00799_, _00798_, _00792_);
  nor _33439_ (_00800_, _00765_, _00782_);
  nor _33440_ (_00801_, _00800_, _00764_);
  nor _33441_ (_00802_, _00786_, _00698_);
  nor _33442_ (_00803_, _00802_, _00801_);
  nor _33443_ (_00804_, _00803_, _00608_);
  nand _33444_ (_00805_, _00793_, _00608_);
  nand _33445_ (_00806_, _00805_, _00606_);
  nor _33446_ (_00807_, _00806_, _00804_);
  nand _33447_ (_00808_, _00786_, _00604_);
  nand _33448_ (_00809_, _00808_, _00603_);
  nor _33449_ (_00810_, _00809_, _00807_);
  nor _33450_ (_00811_, _00669_, _00602_);
  nor _33451_ (_00812_, _00793_, _00669_);
  nor _33452_ (_00813_, _00812_, _00811_);
  nor _33453_ (_00814_, _00813_, _00810_);
  nor _33454_ (_00815_, _00814_, _00799_);
  nor _33455_ (_00816_, _00815_, _00537_);
  nor _33456_ (_00817_, _00816_, _00783_);
  nor _33457_ (_15382_, _00817_, rst);
  nand _33458_ (_00818_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  nand _33459_ (_00819_, _00408_, _25099_);
  nand _33460_ (_15403_, _00819_, _00818_);
  nand _33461_ (_00820_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  nand _33462_ (_00822_, _00408_, _24830_);
  nand _33463_ (_15454_, _00822_, _00820_);
  nand _33464_ (_00823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _26487_);
  nor _33465_ (_15524_, _00823_, _00536_);
  nand _33466_ (_00824_, _00609_, _00698_);
  nor _33467_ (_00825_, _00824_, _00594_);
  nand _33468_ (_00826_, _00825_, _00598_);
  nor _33469_ (_00827_, _00826_, _00590_);
  nor _33470_ (_00828_, _00586_, _00549_);
  nor _33471_ (_00829_, _00583_, _00570_);
  nand _33472_ (_00830_, _00829_, _00828_);
  nand _33473_ (_00831_, _00830_, _00536_);
  nor _33474_ (_00832_, _00831_, _00827_);
  not _33475_ (_00833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nand _33476_ (_00834_, _00537_, _00833_);
  nand _33477_ (_00835_, _00834_, _26487_);
  nor _33478_ (_15545_, _00835_, _00832_);
  nand _33479_ (_00836_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  nand _33480_ (_00837_, _00636_, _24789_);
  nand _33481_ (_15566_, _00837_, _00836_);
  nor _33482_ (_00838_, _00590_, _00537_);
  nor _33483_ (_00839_, _00838_, _00535_);
  nor _33484_ (_00840_, _00537_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _33485_ (_00841_, _00840_, _00642_);
  nand _33486_ (_00842_, _00841_, _26487_);
  nor _33487_ (_15857_, _00842_, _00839_);
  nor _33488_ (_00843_, _28073_, _24073_);
  not _33489_ (_00844_, _00843_);
  nand _33490_ (_00845_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  nand _33491_ (_00846_, _00843_, _24927_);
  nand _33492_ (_15938_, _00846_, _00845_);
  nand _33493_ (_00847_, _24985_, _24830_);
  nand _33494_ (_00848_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  nand _33495_ (_15959_, _00848_, _00847_);
  nand _33496_ (_00849_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  nand _33497_ (_00850_, _00843_, _24789_);
  nand _33498_ (_15990_, _00850_, _00849_);
  nand _33499_ (_00851_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nand _33500_ (_00852_, _00843_, _25150_);
  nand _33501_ (_16061_, _00852_, _00851_);
  nand _33502_ (_00853_, _00735_, _24927_);
  nand _33503_ (_00854_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  nand _33504_ (_16092_, _00854_, _00853_);
  nand _33505_ (_00855_, _00735_, _25039_);
  nand _33506_ (_00856_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  nand _33507_ (_16163_, _00856_, _00855_);
  nand _33508_ (_00857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _26487_);
  nor _33509_ (_16265_, _00857_, _00536_);
  not _33510_ (_00858_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor _33511_ (_00859_, _00536_, _00858_);
  nor _33512_ (_00860_, _00859_, _00643_);
  nor _33513_ (_16306_, _00860_, rst);
  not _33514_ (_00861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor _33515_ (_00862_, _00536_, _00861_);
  nor _33516_ (_00863_, _00862_, _00643_);
  nor _33517_ (_16327_, _00863_, rst);
  nand _33518_ (_00864_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  nand _33519_ (_00865_, _00636_, _25203_);
  nand _33520_ (_16699_, _00865_, _00864_);
  nand _33521_ (_00866_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nand _33522_ (_00867_, _00636_, _28096_);
  nand _33523_ (_16780_, _00867_, _00866_);
  nand _33524_ (_00868_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nand _33525_ (_00869_, _00636_, _25099_);
  nand _33526_ (_16841_, _00869_, _00868_);
  nand _33527_ (_00870_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  nand _33528_ (_00871_, _00636_, _24830_);
  nand _33529_ (_16902_, _00871_, _00870_);
  nand _33530_ (_00872_, _00735_, _25099_);
  nand _33531_ (_00873_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  nand _33532_ (_16923_, _00873_, _00872_);
  nor _33533_ (_00874_, _25465_, _25416_);
  not _33534_ (_00875_, _25402_);
  nor _33535_ (_00876_, _00875_, _25482_);
  nor _33536_ (_00877_, _00876_, _00874_);
  nor _33537_ (_00878_, _25295_, _25266_);
  nand _33538_ (_00879_, _00878_, _25402_);
  not _33539_ (_00880_, _00879_);
  nand _33540_ (_00881_, _00880_, _25235_);
  nand _33541_ (_00882_, _00881_, _00877_);
  nor _33542_ (_00883_, _24864_, rst);
  not _33543_ (_00884_, _00883_);
  nor _33544_ (_00885_, _00884_, _00874_);
  nand _33545_ (_28184_[2], _00885_, _00882_);
  not _33546_ (_00887_, _27813_);
  nor _33547_ (_00888_, _27815_, _27765_);
  not _33548_ (_00889_, _27897_);
  nor _33549_ (_00890_, _27746_, _27732_);
  nand _33550_ (_00891_, _00890_, _27783_);
  nand _33551_ (_00892_, _00891_, _00889_);
  nor _33552_ (_00893_, _00892_, _00888_);
  nand _33553_ (_00894_, _00893_, _00887_);
  nor _33554_ (_00895_, _27852_, _27728_);
  nand _33555_ (_00896_, _00895_, _27733_);
  nand _33556_ (_00897_, _00896_, _27890_);
  nor _33557_ (_00898_, _00897_, _00894_);
  nor _33558_ (_00899_, _27819_, _27781_);
  nor _33559_ (_00900_, _27831_, _27784_);
  nor _33560_ (_00901_, _00900_, _00899_);
  nor _33561_ (_00902_, _27888_, _27728_);
  nand _33562_ (_00903_, _27730_, _27732_);
  nor _33563_ (_00904_, _27784_, _00903_);
  nor _33564_ (_00905_, _00904_, _00902_);
  nand _33565_ (_00906_, _00905_, _00901_);
  nand _33566_ (_00908_, _27806_, _27796_);
  not _33567_ (_00909_, _27916_);
  nand _33568_ (_00910_, _00909_, _00908_);
  nand _33569_ (_00911_, _27747_, _27724_);
  nand _33570_ (_00912_, _00890_, _27806_);
  nand _33571_ (_00913_, _00912_, _00911_);
  nor _33572_ (_00914_, _00913_, _00910_);
  nor _33573_ (_00915_, _27881_, _27795_);
  nand _33574_ (_00916_, _00915_, _00914_);
  nor _33575_ (_00917_, _00916_, _00906_);
  nand _33576_ (_00918_, _00917_, _00898_);
  nand _33577_ (_00919_, _00918_, _24865_);
  nor _33578_ (_00920_, _24860_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _33579_ (_00921_, _00920_);
  nor _33580_ (_00922_, _00921_, \oc8051_top_1.oc8051_decoder1.state [0]);
  nor _33581_ (_00923_, _00922_, _25501_);
  nor _33582_ (_00924_, _00923_, rst);
  nand _33583_ (_28185_[1], _00924_, _00919_);
  nor _33584_ (_00925_, _24997_, _24057_);
  not _33585_ (_00926_, _00925_);
  nor _33586_ (_00927_, _00926_, _24993_);
  nand _33587_ (_00928_, _00927_, _28096_);
  not _33588_ (_00929_, _00927_);
  nand _33589_ (_00930_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nand _33590_ (_17272_, _00930_, _00928_);
  nand _33591_ (_00931_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nand _33592_ (_00932_, _25203_, _25052_);
  nand _33593_ (_17283_, _00932_, _00931_);
  nor _33594_ (_00933_, _00122_, _24073_);
  not _33595_ (_00934_, _00933_);
  nand _33596_ (_00935_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  nand _33597_ (_00936_, _00933_, _24789_);
  nand _33598_ (_17344_, _00936_, _00935_);
  nand _33599_ (_00937_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  nand _33600_ (_00938_, _00933_, _25150_);
  nand _33601_ (_17475_, _00938_, _00937_);
  nand _33602_ (_00939_, _25152_, _24927_);
  nand _33603_ (_00940_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  nand _33604_ (_17786_, _00940_, _00939_);
  not _33605_ (_00941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not _33606_ (_00942_, _00642_);
  nor _33607_ (_00943_, _00942_, _00941_);
  nor _33608_ (_00944_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _00535_);
  not _33609_ (_00945_, _00944_);
  nand _33610_ (_00946_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _00535_);
  nand _33611_ (_00947_, _00946_, _00945_);
  nand _33612_ (_00948_, _00947_, _00590_);
  nand _33613_ (_00949_, _00948_, _00536_);
  nor _33614_ (_00950_, _00949_, _00943_);
  nand _33615_ (_00951_, _00947_, _00537_);
  nand _33616_ (_00952_, _00951_, _26487_);
  nor _33617_ (_17867_, _00952_, _00950_);
  nor _33618_ (_00953_, _25045_, _24976_);
  not _33619_ (_00954_, _00953_);
  nor _33620_ (_00955_, _00954_, _28057_);
  nand _33621_ (_00956_, _00955_, _24830_);
  not _33622_ (_00957_, _00955_);
  nand _33623_ (_00958_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  nand _33624_ (_17928_, _00958_, _00956_);
  nand _33625_ (_00959_, _25152_, _24789_);
  nand _33626_ (_00960_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  nand _33627_ (_18055_, _00960_, _00959_);
  nand _33628_ (_00961_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nand _33629_ (_00962_, _00843_, _28096_);
  nand _33630_ (_18111_, _00962_, _00961_);
  nand _33631_ (_00963_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  nand _33632_ (_00964_, _00843_, _25099_);
  nand _33633_ (_18222_, _00964_, _00963_);
  nand _33634_ (_00965_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  nand _33635_ (_00966_, _00843_, _24830_);
  nand _33636_ (_18241_, _00966_, _00965_);
  nand _33637_ (_00967_, _28063_, _25039_);
  nand _33638_ (_00968_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  nand _33639_ (_18261_, _00968_, _00967_);
  nand _33640_ (_00969_, _00927_, _24927_);
  nand _33641_ (_00970_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  nand _33642_ (_18361_, _00970_, _00969_);
  nand _33643_ (_00971_, _00927_, _25039_);
  nand _33644_ (_00972_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nand _33645_ (_18400_, _00972_, _00971_);
  nand _33646_ (_00973_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  nand _33647_ (_00974_, _00933_, _24830_);
  nand _33648_ (_18585_, _00974_, _00973_);
  nand _33649_ (_00975_, _00927_, _24789_);
  nand _33650_ (_00976_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nand _33651_ (_18635_, _00976_, _00975_);
  nand _33652_ (_00977_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  nand _33653_ (_00978_, _00933_, _28096_);
  nand _33654_ (_18653_, _00978_, _00977_);
  nor _33655_ (_00979_, _00629_, _25165_);
  nand _33656_ (_00980_, _00979_, _24830_);
  not _33657_ (_00981_, _00979_);
  nand _33658_ (_00982_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nand _33659_ (_18710_, _00982_, _00980_);
  nand _33660_ (_00983_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nand _33661_ (_00984_, _00933_, _25099_);
  nand _33662_ (_18742_, _00984_, _00983_);
  nor _33663_ (_00985_, _25059_, _24059_);
  nand _33664_ (_00986_, _00985_, _24789_);
  not _33665_ (_00987_, _00985_);
  nand _33666_ (_00988_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  nand _33667_ (_18851_, _00988_, _00986_);
  nand _33668_ (_00989_, _00985_, _25150_);
  nand _33669_ (_00990_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nand _33670_ (_18879_, _00990_, _00989_);
  nor _33671_ (_00991_, _25059_, _24882_);
  nand _33672_ (_00992_, _00991_, _25039_);
  not _33673_ (_00993_, _00991_);
  nand _33674_ (_00994_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  nand _33675_ (_18983_, _00994_, _00992_);
  nor _33676_ (_00995_, _24984_, _28080_);
  nand _33677_ (_00996_, _00995_, _24927_);
  not _33678_ (_00997_, _00995_);
  nand _33679_ (_00998_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  nand _33680_ (_19021_, _00998_, _00996_);
  nor _33681_ (_00999_, _25157_, _24887_);
  not _33682_ (_01000_, _00999_);
  nor _33683_ (_01001_, _01000_, _24978_);
  nand _33684_ (_01002_, _01001_, _28096_);
  not _33685_ (_01003_, _01001_);
  nand _33686_ (_01004_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  nand _33687_ (_19097_, _01004_, _01002_);
  nand _33688_ (_01005_, _00995_, _28096_);
  nand _33689_ (_01006_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  nand _33690_ (_19311_, _01006_, _01005_);
  nand _33691_ (_01007_, _00995_, _25039_);
  nand _33692_ (_01008_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  nand _33693_ (_19422_, _01008_, _01007_);
  nor _33694_ (_01009_, _25059_, _24795_);
  nand _33695_ (_01010_, _01009_, _25203_);
  not _33696_ (_01011_, _01009_);
  nand _33697_ (_01012_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  nand _33698_ (_19503_, _01012_, _01010_);
  nand _33699_ (_01013_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  nand _33700_ (_01014_, _00933_, _25039_);
  nand _33701_ (_19554_, _01014_, _01013_);
  nand _33702_ (_01015_, _01009_, _28096_);
  nand _33703_ (_01016_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  nand _33704_ (_19605_, _01016_, _01015_);
  nand _33705_ (_01017_, _01009_, _25099_);
  nand _33706_ (_01018_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  nand _33707_ (_19656_, _01018_, _01017_);
  nand _33708_ (_01019_, _00394_, _25099_);
  nand _33709_ (_01020_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  nand _33710_ (_19717_, _01020_, _01019_);
  nor _33711_ (_28183_[2], _25816_, rst);
  nor _33712_ (_01021_, _25572_, _25509_);
  not _33713_ (_01022_, _25587_);
  not _33714_ (_01023_, _25588_);
  nor _33715_ (_01024_, _01023_, _01022_);
  nand _33716_ (_01025_, _01024_, _25579_);
  nor _33717_ (_01026_, _01025_, _01021_);
  not _33718_ (_01027_, _25584_);
  nand _33719_ (_01028_, _01027_, _25533_);
  not _33720_ (_01029_, _25554_);
  nand _33721_ (_01030_, _25575_, _01029_);
  not _33722_ (_01031_, _01030_);
  not _33723_ (_01032_, _25605_);
  nor _33724_ (_01033_, _00875_, _25329_);
  nor _33725_ (_01034_, _01033_, _25474_);
  nor _33726_ (_01035_, _01034_, _25551_);
  nor _33727_ (_01036_, _01035_, _01032_);
  nand _33728_ (_01037_, _01036_, _25568_);
  nor _33729_ (_01038_, _01037_, _25556_);
  nand _33730_ (_01039_, _01038_, _01031_);
  nor _33731_ (_01040_, _01039_, _01028_);
  nand _33732_ (_01041_, _01040_, _01026_);
  nor _33733_ (_01042_, _25412_, _25401_);
  not _33734_ (_01043_, _25424_);
  nand _33735_ (_01044_, _25599_, _01043_);
  nor _33736_ (_01045_, _01044_, _01042_);
  nor _33737_ (_01046_, _26195_, _25401_);
  nor _33738_ (_01047_, _01046_, _25546_);
  nor _33739_ (_01048_, _25327_, _25235_);
  not _33740_ (_01049_, _01048_);
  nor _33741_ (_01050_, _01049_, _25420_);
  nor _33742_ (_01051_, _01050_, _25421_);
  not _33743_ (_01052_, _01051_);
  nor _33744_ (_01053_, _01049_, _25416_);
  nand _33745_ (_01054_, _26139_, _25327_);
  not _33746_ (_01055_, _01054_);
  nor _33747_ (_01056_, _01055_, _01053_);
  not _33748_ (_01057_, _01056_);
  nor _33749_ (_01058_, _01057_, _01052_);
  nand _33750_ (_01059_, _01058_, _01047_);
  nor _33751_ (_01060_, _01049_, _25423_);
  not _33752_ (_01061_, _25423_);
  nor _33753_ (_01062_, _01061_, _25418_);
  nor _33754_ (_01063_, _01062_, _26195_);
  nor _33755_ (_01064_, _01063_, _01060_);
  not _33756_ (_01065_, _25603_);
  nor _33757_ (_01066_, _01065_, _25494_);
  nand _33758_ (_01067_, _01066_, _01064_);
  nor _33759_ (_01068_, _01067_, _01059_);
  nand _33760_ (_01069_, _01068_, _01045_);
  nor _33761_ (_01070_, _01069_, _01041_);
  nor _33762_ (_01071_, _01070_, _24864_);
  nand _33763_ (_01072_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _33764_ (_01073_, _01055_, _01021_);
  nor _33765_ (_01074_, _01073_, _25505_);
  nor _33766_ (_01075_, _01074_, _00101_);
  not _33767_ (_01076_, _01075_);
  nor _33768_ (_01077_, _25541_, _25505_);
  nor _33769_ (_01078_, _01077_, _01076_);
  nand _33770_ (_01079_, _01078_, _01072_);
  nor _33771_ (_01080_, _01079_, _01071_);
  nor _33772_ (_28195_, _01080_, rst);
  nand _33773_ (_01081_, _00985_, _25099_);
  nand _33774_ (_01082_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nand _33775_ (_19921_, _01082_, _01081_);
  nand _33776_ (_01083_, _00985_, _24830_);
  nand _33777_ (_01084_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  nand _33778_ (_19973_, _01084_, _01083_);
  nor _33779_ (_01085_, _25047_, _24073_);
  not _33780_ (_01086_, _01085_);
  nand _33781_ (_01087_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  nand _33782_ (_01088_, _01085_, _25203_);
  nand _33783_ (_19987_, _01088_, _01087_);
  nor _33784_ (_28182_[5], _27732_, rst);
  nand _33785_ (_01089_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  nand _33786_ (_01090_, _01085_, _28096_);
  nand _33787_ (_20109_, _01090_, _01089_);
  nand _33788_ (_01091_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nand _33789_ (_01093_, _01085_, _25099_);
  nand _33790_ (_20174_, _01093_, _01091_);
  nand _33791_ (_01094_, _00985_, _25039_);
  nand _33792_ (_01095_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  nand _33793_ (_20263_, _01095_, _01094_);
  nand _33794_ (_01096_, _00985_, _25203_);
  nand _33795_ (_01097_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nand _33796_ (_20330_, _01097_, _01096_);
  nand _33797_ (_01098_, _00985_, _28096_);
  nand _33798_ (_01099_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nand _33799_ (_20409_, _01099_, _01098_);
  nand _33800_ (_01100_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  nand _33801_ (_01101_, _01085_, _24927_);
  nand _33802_ (_20458_, _01101_, _01100_);
  nand _33803_ (_01102_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  nand _33804_ (_01103_, _01085_, _25150_);
  nand _33805_ (_20605_, _01103_, _01102_);
  nor _33806_ (_01104_, _25057_, _24984_);
  nand _33807_ (_01105_, _01104_, _28096_);
  not _33808_ (_01106_, _01104_);
  nand _33809_ (_01107_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nand _33810_ (_20873_, _01107_, _01105_);
  nor _33811_ (_01108_, _01000_, _00114_);
  nand _33812_ (_01109_, _01108_, _25039_);
  not _33813_ (_01110_, _01108_);
  nand _33814_ (_01111_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nand _33815_ (_20898_, _01111_, _01109_);
  nand _33816_ (_01112_, _00995_, _24789_);
  nand _33817_ (_01113_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  nand _33818_ (_21000_, _01113_, _01112_);
  nand _33819_ (_01114_, _01104_, _24830_);
  nand _33820_ (_01115_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nand _33821_ (_21036_, _01115_, _01114_);
  nor _33822_ (_01116_, _01000_, _24999_);
  nand _33823_ (_01117_, _01116_, _24789_);
  not _33824_ (_01118_, _01116_);
  nand _33825_ (_01119_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  nand _33826_ (_21091_, _01119_, _01117_);
  nor _33827_ (_01120_, _28073_, _24984_);
  nand _33828_ (_01121_, _01120_, _28096_);
  not _33829_ (_01123_, _01120_);
  nand _33830_ (_01124_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nand _33831_ (_21130_, _01124_, _01121_);
  nand _33832_ (_01125_, _01104_, _25039_);
  nand _33833_ (_01126_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nand _33834_ (_21268_, _01126_, _01125_);
  nand _33835_ (_01127_, _01104_, _25150_);
  nand _33836_ (_01128_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nand _33837_ (_21283_, _01128_, _01127_);
  nor _33838_ (_01129_, _00415_, _24073_);
  not _33839_ (_01130_, _01129_);
  nand _33840_ (_01131_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  nand _33841_ (_01132_, _01129_, _25039_);
  nand _33842_ (_21304_, _01132_, _01131_);
  nand _33843_ (_01133_, _01104_, _25203_);
  nand _33844_ (_01134_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nand _33845_ (_21572_, _01134_, _01133_);
  nand _33846_ (_01135_, _00995_, _25150_);
  nand _33847_ (_01136_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  nand _33848_ (_21623_, _01136_, _01135_);
  nand _33849_ (_01137_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nand _33850_ (_01138_, _01129_, _25150_);
  nand _33851_ (_21654_, _01138_, _01137_);
  nor _33852_ (_01140_, _00926_, _25059_);
  nand _33853_ (_01141_, _01140_, _24789_);
  not _33854_ (_01142_, _01140_);
  nand _33855_ (_01143_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  nand _33856_ (_21845_, _01143_, _01141_);
  nand _33857_ (_01144_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  nand _33858_ (_01145_, _01129_, _24927_);
  nand _33859_ (_22016_, _01145_, _01144_);
  nand _33860_ (_01146_, _01108_, _28096_);
  nand _33861_ (_01147_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  nand _33862_ (_22242_, _01147_, _01146_);
  nand _33863_ (_01149_, _01108_, _25099_);
  nand _33864_ (_01150_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nand _33865_ (_22307_, _01150_, _01149_);
  nand _33866_ (_01151_, _01108_, _24830_);
  nand _33867_ (_01152_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  nand _33868_ (_22334_, _01152_, _01151_);
  nor _33869_ (_01153_, _00629_, _28057_);
  nand _33870_ (_01154_, _01153_, _25150_);
  not _33871_ (_01155_, _01153_);
  nand _33872_ (_01156_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nand _33873_ (_22413_, _01156_, _01154_);
  nand _33874_ (_01157_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  nand _33875_ (_01158_, _01085_, _24830_);
  nand _33876_ (_22462_, _01158_, _01157_);
  nand _33877_ (_01159_, _01140_, _25099_);
  nand _33878_ (_01160_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  nand _33879_ (_22593_, _01160_, _01159_);
  nand _33880_ (_01161_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  nand _33881_ (_01162_, _01129_, _24789_);
  nand _33882_ (_22674_, _01162_, _01161_);
  nand _33883_ (_01163_, _01140_, _24830_);
  nand _33884_ (_01164_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nand _33885_ (_22695_, _01164_, _01163_);
  nand _33886_ (_01165_, _01009_, _24789_);
  nand _33887_ (_01166_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nand _33888_ (_22786_, _01166_, _01165_);
  nand _33889_ (_01167_, _01140_, _25203_);
  nand _33890_ (_01169_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  nand _33891_ (_23037_, _01169_, _01167_);
  nand _33892_ (_01170_, _01140_, _24927_);
  nand _33893_ (_01171_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  nand _33894_ (_23058_, _01171_, _01170_);
  nand _33895_ (_01172_, _01140_, _25039_);
  nand _33896_ (_01173_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  nand _33897_ (_23199_, _01173_, _01172_);
  nor _33898_ (_01174_, _00954_, _24073_);
  not _33899_ (_01175_, _01174_);
  nand _33900_ (_01176_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  nand _33901_ (_01177_, _01174_, _24789_);
  nand _33902_ (_23350_, _01177_, _01176_);
  nor _33903_ (_01178_, _00926_, _25159_);
  nand _33904_ (_01179_, _01178_, _24830_);
  not _33905_ (_01180_, _01178_);
  nand _33906_ (_01181_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand _33907_ (_23552_, _01181_, _01179_);
  nor _33908_ (_01182_, _28057_, _24999_);
  nand _33909_ (_01183_, _01182_, _25099_);
  not _33910_ (_01185_, _01182_);
  nand _33911_ (_01186_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  nand _33912_ (_23654_, _01186_, _01183_);
  nand _33913_ (_01187_, _01009_, _25150_);
  nand _33914_ (_01188_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  nand _33915_ (_23680_, _01188_, _01187_);
  nand _33916_ (_01190_, _25160_, _24830_);
  nand _33917_ (_01191_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand _33918_ (_23681_, _01191_, _01190_);
  nand _33919_ (_01192_, _01009_, _24927_);
  nand _33920_ (_01193_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  nand _33921_ (_23682_, _01193_, _01192_);
  nand _33922_ (_01194_, _28081_, _25039_);
  nand _33923_ (_01195_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  nand _33924_ (_23683_, _01195_, _01194_);
  nand _33925_ (_01196_, _28105_, _24789_);
  nand _33926_ (_01197_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nand _33927_ (_23684_, _01197_, _01196_);
  nand _33928_ (_01198_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  nand _33929_ (_01199_, _01129_, _25099_);
  nand _33930_ (_23685_, _01199_, _01198_);
  not _33931_ (_01200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nand _33932_ (_01201_, _00223_, _24840_);
  nand _33933_ (_01202_, _01201_, _01200_);
  nand _33934_ (_01203_, _01202_, _00375_);
  nor _33935_ (_01204_, _01201_, _24716_);
  nor _33936_ (_01205_, _01204_, _01203_);
  nor _33937_ (_01206_, _00375_, _25088_);
  nor _33938_ (_01207_, _01206_, _01205_);
  nor _33939_ (_23686_, _01207_, rst);
  nor _33940_ (_01208_, _25059_, _24999_);
  nand _33941_ (_01209_, _01208_, _25203_);
  not _33942_ (_01210_, _01208_);
  nand _33943_ (_01211_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nand _33944_ (_23687_, _01211_, _01209_);
  nand _33945_ (_01212_, _28081_, _25203_);
  nand _33946_ (_01213_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nand _33947_ (_23688_, _01213_, _01212_);
  nand _33948_ (_01214_, _01208_, _28096_);
  nand _33949_ (_01215_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  nand _33950_ (_23689_, _01215_, _01214_);
  nor _33951_ (_01216_, _00415_, _25051_);
  not _33952_ (_01217_, _01216_);
  nand _33953_ (_01218_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  nand _33954_ (_01219_, _01216_, _25099_);
  nand _33955_ (_23690_, _01219_, _01218_);
  nor _33956_ (_28182_[1], _25262_, rst);
  nor _33957_ (_28182_[3], _25231_, rst);
  nor _33958_ (_28182_[0], _27763_, rst);
  nor _33959_ (_28182_[2], _27755_, rst);
  nand _33960_ (_01221_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  nand _33961_ (_01222_, _01174_, _28096_);
  nand _33962_ (_23691_, _01222_, _01221_);
  nand _33963_ (_01224_, _01208_, _24789_);
  nand _33964_ (_01226_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  nand _33965_ (_23692_, _01226_, _01224_);
  nand _33966_ (_01228_, _01208_, _25150_);
  nand _33967_ (_01229_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  nand _33968_ (_23693_, _01229_, _01228_);
  nand _33969_ (_01230_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nand _33970_ (_01231_, _01174_, _25099_);
  nand _33971_ (_23694_, _01231_, _01230_);
  nand _33972_ (_01232_, _01208_, _24927_);
  nand _33973_ (_01233_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  nand _33974_ (_23695_, _01233_, _01232_);
  nand _33975_ (_01234_, _25061_, _24927_);
  nand _33976_ (_01236_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  nand _33977_ (_23696_, _01236_, _01234_);
  nand _33978_ (_01237_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  nand _33979_ (_01238_, _01174_, _24927_);
  nand _33980_ (_23697_, _01238_, _01237_);
  not _33981_ (_01239_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _33982_ (_01240_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _33983_ (_01241_, _01240_);
  nor _33984_ (_01242_, _01241_, _00166_);
  not _33985_ (_01243_, _01242_);
  nor _33986_ (_01245_, _01243_, _01239_);
  nand _33987_ (_01246_, _01241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  nor _33988_ (_01247_, _01246_, _01239_);
  not _33989_ (_01248_, _01247_);
  nor _33990_ (_01249_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _33991_ (_01250_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nand _33992_ (_01251_, _01250_, _01249_);
  nor _33993_ (_01252_, _01251_, _01248_);
  nor _33994_ (_01253_, _01252_, _01245_);
  not _33995_ (_01254_, _01253_);
  nand _33996_ (_01255_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand _33997_ (_01256_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nand _33998_ (_01257_, _01256_, _01255_);
  nor _33999_ (_01258_, _24833_, _24071_);
  nor _34000_ (_01259_, _00137_, _24842_);
  nand _34001_ (_01260_, _01259_, _01258_);
  not _34002_ (_01261_, _01260_);
  nor _34003_ (_01262_, _01261_, rst);
  nand _34004_ (_01263_, _01262_, _01257_);
  nand _34005_ (_01264_, _01240_, _24920_);
  nand _34006_ (_01265_, _01241_, _25028_);
  nand _34007_ (_01266_, _01265_, _01264_);
  nor _34008_ (_01267_, _01260_, rst);
  nand _34009_ (_01269_, _01267_, _01266_);
  nand _34010_ (_23698_, _01269_, _01263_);
  not _34011_ (_01271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  not _34012_ (_01272_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nand _34013_ (_01274_, _01272_, _01271_);
  not _34014_ (_01275_, _00221_);
  nor _34015_ (_01276_, _01275_, _00617_);
  not _34016_ (_01277_, _01276_);
  nor _34017_ (_01278_, _01277_, _00426_);
  nor _34018_ (_01279_, _01278_, _01274_);
  nand _34019_ (_01280_, _24840_, _24716_);
  not _34020_ (_01281_, _01280_);
  nand _34021_ (_01282_, _24842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _34022_ (_01283_, _01282_, _01278_);
  nor _34023_ (_01284_, _01283_, _01281_);
  nor _34024_ (_01285_, _01284_, _01279_);
  not _34025_ (_01286_, _01258_);
  nor _34026_ (_01287_, _01286_, _00235_);
  nor _34027_ (_01288_, _01287_, _01285_);
  nor _34028_ (_01290_, _01286_, _00373_);
  nand _34029_ (_01291_, _01290_, _25088_);
  nand _34030_ (_01292_, _01291_, _26487_);
  nor _34031_ (_23699_, _01292_, _01288_);
  not _34032_ (_01293_, _01290_);
  not _34033_ (_01294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand _34034_ (_01295_, _01278_, _00444_);
  nand _34035_ (_01296_, _01295_, _01294_);
  nand _34036_ (_01297_, _01296_, _01293_);
  nor _34037_ (_01298_, _01295_, _24716_);
  nor _34038_ (_01299_, _01298_, _01297_);
  nor _34039_ (_01300_, _01293_, _25195_);
  nor _34040_ (_01301_, _01300_, _01299_);
  nor _34041_ (_23700_, _01301_, rst);
  nor _34042_ (_01302_, _01260_, _01241_);
  not _34043_ (_01303_, _01302_);
  nor _34044_ (_01304_, _01303_, _25029_);
  nand _34045_ (_01305_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nand _34046_ (_01306_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand _34047_ (_01307_, _01306_, _01305_);
  nand _34048_ (_01308_, _01307_, _01260_);
  nor _34049_ (_01309_, _01260_, _01240_);
  nand _34050_ (_01310_, _01309_, _25194_);
  nand _34051_ (_01312_, _01310_, _01308_);
  nor _34052_ (_01313_, _01312_, _01304_);
  nor _34053_ (_23701_, _01313_, rst);
  not _34054_ (_01314_, _01309_);
  nor _34055_ (_01315_, _01314_, _25703_);
  nand _34056_ (_01316_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand _34057_ (_01317_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nand _34058_ (_01318_, _01317_, _01316_);
  nand _34059_ (_01319_, _01318_, _01260_);
  nand _34060_ (_01320_, _01302_, _25194_);
  nand _34061_ (_01321_, _01320_, _01319_);
  nor _34062_ (_01322_, _01321_, _01315_);
  nor _34063_ (_23702_, _01322_, rst);
  nor _34064_ (_01323_, _01303_, _25703_);
  nand _34065_ (_01324_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nand _34066_ (_01325_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nand _34067_ (_01326_, _01325_, _01324_);
  nand _34068_ (_01327_, _01326_, _01260_);
  nand _34069_ (_01328_, _01309_, _25089_);
  nand _34070_ (_01329_, _01328_, _01327_);
  nor _34071_ (_01330_, _01329_, _01323_);
  nor _34072_ (_23703_, _01330_, rst);
  nor _34073_ (_01331_, _01303_, _25088_);
  nand _34074_ (_01332_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nand _34075_ (_01333_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nand _34076_ (_01334_, _01333_, _01332_);
  nand _34077_ (_01335_, _01334_, _01260_);
  nand _34078_ (_01336_, _01309_, _24821_);
  nand _34079_ (_01337_, _01336_, _01335_);
  nor _34080_ (_01338_, _01337_, _01331_);
  nor _34081_ (_23704_, _01338_, rst);
  nor _34082_ (_01339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not _34083_ (_01340_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _34084_ (_01341_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  not _34085_ (_01342_, _01341_);
  nor _34086_ (_01343_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _34087_ (_01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nand _34088_ (_01345_, _01344_, _01343_);
  nor _34089_ (_01346_, _01345_, _01342_);
  not _34090_ (_01347_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _34091_ (_01348_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nand _34092_ (_01349_, _01348_, _01347_);
  nor _34093_ (_01350_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nand _34094_ (_01351_, _01350_, _01346_);
  nand _34095_ (_01352_, _01351_, _01340_);
  nand _34096_ (_01354_, _01352_, _01245_);
  nor _34097_ (_01355_, _01354_, _01339_);
  nor _34098_ (_01357_, _01252_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not _34099_ (_01358_, _01245_);
  nand _34100_ (_01360_, _01252_, _01340_);
  nand _34101_ (_01361_, _01360_, _01358_);
  nor _34102_ (_01362_, _01361_, _01357_);
  nor _34103_ (_01363_, _01362_, _01355_);
  nor _34104_ (_01364_, _01363_, _01261_);
  nand _34105_ (_01366_, _01240_, _24821_);
  nor _34106_ (_01367_, _01366_, _01260_);
  nor _34107_ (_01368_, _01367_, _01364_);
  nor _34108_ (_23705_, _01368_, rst);
  nand _34109_ (_01369_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  nand _34110_ (_01370_, _01174_, _25039_);
  nand _34111_ (_23706_, _01370_, _01369_);
  nor _34112_ (_01371_, _28073_, _28057_);
  nand _34113_ (_01372_, _01371_, _25203_);
  not _34114_ (_01373_, _01371_);
  nand _34115_ (_01374_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  nand _34116_ (_23707_, _01374_, _01372_);
  nand _34117_ (_01375_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  nand _34118_ (_01376_, _01174_, _25203_);
  nand _34119_ (_23708_, _01376_, _01375_);
  not _34120_ (_01377_, _01262_);
  not _34121_ (_01378_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  not _34122_ (_01379_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nand _34123_ (_01380_, _01247_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _34124_ (_01381_, _01380_, _01379_);
  not _34125_ (_01382_, _01381_);
  nor _34126_ (_01383_, _01382_, _01378_);
  not _34127_ (_01384_, _01383_);
  nand _34128_ (_01385_, _01382_, _01378_);
  nand _34129_ (_01386_, _01385_, _01384_);
  nor _34130_ (_23709_, _01386_, _01377_);
  nor _34131_ (_01388_, _00926_, _24073_);
  not _34132_ (_01389_, _01388_);
  nand _34133_ (_01391_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  nand _34134_ (_01392_, _01388_, _24927_);
  nand _34135_ (_23710_, _01392_, _01391_);
  nand _34136_ (_01393_, _01380_, _01379_);
  nand _34137_ (_01394_, _01393_, _01382_);
  nor _34138_ (_23711_, _01394_, _01377_);
  not _34139_ (_01395_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nand _34140_ (_01396_, _01248_, _01395_);
  nand _34141_ (_01397_, _01396_, _01380_);
  nor _34142_ (_23712_, _01397_, _01377_);
  nor _34143_ (_01398_, _28073_, _25059_);
  nand _34144_ (_01399_, _01398_, _25203_);
  not _34145_ (_01400_, _01398_);
  nand _34146_ (_01401_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  nand _34147_ (_23713_, _01401_, _01399_);
  nor _34148_ (_01402_, _00629_, _24889_);
  nand _34149_ (_01403_, _01402_, _25203_);
  not _34150_ (_01404_, _01402_);
  nand _34151_ (_01405_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nand _34152_ (_23714_, _01405_, _01403_);
  nand _34153_ (_01406_, _01208_, _24830_);
  nand _34154_ (_01407_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nand _34155_ (_23715_, _01407_, _01406_);
  nand _34156_ (_01408_, _25061_, _24789_);
  nand _34157_ (_01409_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  nand _34158_ (_23716_, _01409_, _01408_);
  nor _34159_ (_01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  nand _34160_ (_01413_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not _34161_ (_01414_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _34162_ (_01415_, _01414_, rst);
  nand _34163_ (_01416_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  nand _34164_ (_23717_, _01416_, _01413_);
  nand _34165_ (_01418_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nand _34166_ (_01419_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  nand _34167_ (_23718_, _01419_, _01418_);
  nand _34168_ (_01420_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  nand _34169_ (_01421_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand _34170_ (_23719_, _01421_, _01420_);
  nand _34171_ (_01422_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  nand _34172_ (_01423_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  nand _34173_ (_23720_, _01423_, _01422_);
  nand _34174_ (_01424_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  nand _34175_ (_01425_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  nand _34176_ (_23721_, _01425_, _01424_);
  not _34177_ (_01426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not _34178_ (_01427_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  nor _34179_ (_01428_, _01427_, _01426_);
  not _34180_ (_01429_, _01428_);
  nor _34181_ (_01430_, _01429_, _01240_);
  not _34182_ (_01431_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _34183_ (_01432_, _01431_, _01427_);
  not _34184_ (_01433_, _01432_);
  nor _34185_ (_01434_, _01433_, _01240_);
  not _34186_ (_01435_, _01434_);
  nor _34187_ (_01436_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01426_);
  nor _34188_ (_01437_, _01241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _34189_ (_01438_, _01437_, _01436_);
  nand _34190_ (_01440_, _01438_, _01435_);
  nor _34191_ (_01441_, _01440_, _01430_);
  not _34192_ (_01443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _34193_ (_01444_, _01443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not _34194_ (_01445_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _34195_ (_01447_, _01445_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nand _34196_ (_01448_, _01447_, _01444_);
  not _34197_ (_01450_, _01448_);
  nor _34198_ (_01452_, _01450_, _01435_);
  nor _34199_ (_01453_, _01452_, _01441_);
  not _34200_ (_01454_, _01453_);
  nor _34201_ (_01456_, _01243_, _01431_);
  nor _34202_ (_01457_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  nand _34203_ (_01459_, _01457_, _01454_);
  not _34204_ (_01460_, _01415_);
  nor _34205_ (_01461_, _01448_, _01435_);
  nor _34206_ (_01462_, _01461_, _01456_);
  nor _34207_ (_01463_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  nor _34208_ (_01464_, _01463_, _01460_);
  nand _34209_ (_01465_, _01464_, _01459_);
  nand _34210_ (_23722_, _01465_, _01424_);
  not _34211_ (_01467_, _01462_);
  nand _34212_ (_01468_, _01467_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  not _34213_ (_01470_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor _34214_ (_01471_, _01456_, _01470_);
  nand _34215_ (_01473_, _01471_, _01454_);
  nand _34216_ (_01474_, _01473_, _01468_);
  nand _34217_ (_01475_, _01474_, _01415_);
  nand _34218_ (_23723_, _01475_, _01413_);
  not _34219_ (_01476_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _34220_ (_01477_, _01240_, _01414_);
  nand _34221_ (_01479_, _01477_, _01432_);
  nand _34222_ (_01480_, _01430_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nand _34223_ (_01481_, _01480_, _01479_);
  nor _34224_ (_01482_, _01481_, _01476_);
  nor _34225_ (_01483_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01476_);
  nor _34226_ (_01484_, _01483_, _01447_);
  nor _34227_ (_01485_, _01484_, _01479_);
  nor _34228_ (_01486_, _01485_, _01482_);
  nor _34229_ (_23724_, _01486_, rst);
  nand _34230_ (_01488_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  nand _34231_ (_01489_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _34232_ (_23725_, _01489_, _01488_);
  nand _34233_ (_01490_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  nor _34234_ (_01491_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  nand _34235_ (_01492_, _01491_, _01454_);
  nor _34236_ (_01493_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  nor _34237_ (_01494_, _01493_, _01460_);
  nand _34238_ (_01496_, _01494_, _01492_);
  nand _34239_ (_23726_, _01496_, _01490_);
  nor _34240_ (_01497_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  nand _34241_ (_01498_, _01497_, _01454_);
  nor _34242_ (_01499_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  nor _34243_ (_01500_, _01499_, _01460_);
  nand _34244_ (_01501_, _01500_, _01498_);
  nand _34245_ (_23727_, _01501_, _01488_);
  not _34246_ (_01502_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  not _34247_ (_01503_, _01456_);
  nand _34248_ (_01504_, _01503_, _01502_);
  nor _34249_ (_01506_, _01504_, _01453_);
  not _34250_ (_01507_, _01410_);
  nor _34251_ (_01508_, _01507_, _01502_);
  nor _34252_ (_01509_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  nor _34253_ (_01511_, _01509_, _01460_);
  nor _34254_ (_01512_, _01511_, _01508_);
  nor _34255_ (_23728_, _01512_, _01506_);
  not _34256_ (_01513_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  nand _34257_ (_01514_, _01503_, _01513_);
  nor _34258_ (_01515_, _01514_, _01453_);
  nor _34259_ (_01516_, _01507_, _01513_);
  nor _34260_ (_01517_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  nor _34261_ (_01518_, _01517_, _01460_);
  nor _34262_ (_01519_, _01518_, _01516_);
  nor _34263_ (_23729_, _01519_, _01515_);
  nor _34264_ (_01520_, _00393_, _24073_);
  not _34265_ (_01521_, _01520_);
  nand _34266_ (_01522_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  nand _34267_ (_01523_, _01520_, _24927_);
  nand _34268_ (_23730_, _01523_, _01522_);
  not _34269_ (_01524_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _34270_ (_01525_, _01503_, _01524_);
  nor _34271_ (_01526_, _01525_, _01453_);
  nor _34272_ (_01527_, _01507_, _01524_);
  nor _34273_ (_01528_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  nor _34274_ (_01529_, _01528_, _01460_);
  nor _34275_ (_01530_, _01529_, _01527_);
  nor _34276_ (_23731_, _01530_, _01526_);
  nand _34277_ (_01531_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nand _34278_ (_01532_, _01520_, _25039_);
  nand _34279_ (_23732_, _01532_, _01531_);
  nor _34280_ (_01533_, _25059_, _24978_);
  nand _34281_ (_01534_, _01533_, _28096_);
  not _34282_ (_01535_, _01533_);
  nand _34283_ (_01536_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nand _34284_ (_23733_, _01536_, _01534_);
  nand _34285_ (_01537_, _01533_, _25099_);
  nand _34286_ (_01538_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  nand _34287_ (_23734_, _01538_, _01537_);
  nor _34288_ (_01539_, _24071_, _25724_);
  not _34289_ (_01540_, _01539_);
  nor _34290_ (_01541_, _01540_, _00436_);
  not _34291_ (_01542_, _01541_);
  nor _34292_ (_01543_, _01542_, _24842_);
  nand _34293_ (_01544_, _01543_, _24717_);
  nor _34294_ (_01545_, _01543_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor _34295_ (_01546_, _01545_, _26245_);
  nand _34296_ (_01547_, _01546_, _01544_);
  nor _34297_ (_01548_, _25723_, _25724_);
  not _34298_ (_01549_, _01548_);
  nor _34299_ (_01550_, _00436_, _01549_);
  nand _34300_ (_01551_, _01550_, _24070_);
  not _34301_ (_01552_, _01551_);
  nand _34302_ (_01553_, _01552_, _25088_);
  nor _34303_ (_01554_, _01552_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor _34304_ (_01555_, _01554_, _25631_);
  nand _34305_ (_01556_, _01555_, _01553_);
  nand _34306_ (_01557_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nand _34307_ (_01558_, _01557_, _01556_);
  nor _34308_ (_01559_, _01558_, rst);
  nand _34309_ (_23735_, _01559_, _01547_);
  nor _34310_ (_01560_, _01542_, _25723_);
  nand _34311_ (_01561_, _01560_, _24717_);
  nor _34312_ (_01562_, _01552_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _34313_ (_01563_, _01562_, _26245_);
  nand _34314_ (_01564_, _01563_, _01561_);
  nand _34315_ (_01565_, _01552_, _24820_);
  nand _34316_ (_01566_, _01565_, _25630_);
  nor _34317_ (_01567_, _01566_, _01562_);
  nand _34318_ (_01568_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nand _34319_ (_01569_, _01568_, _26487_);
  nor _34320_ (_01570_, _01569_, _01567_);
  nand _34321_ (_23736_, _01570_, _01564_);
  nand _34322_ (_01571_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nand _34323_ (_01572_, _01388_, _25150_);
  nand _34324_ (_23737_, _01572_, _01571_);
  nor _34325_ (_01573_, _00278_, _25627_);
  nor _34326_ (_01574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not _34327_ (_01575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not _34328_ (_01577_, t0_i);
  nand _34329_ (_01578_, _01577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  nand _34330_ (_01580_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _34331_ (_01582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _34332_ (_01584_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _34333_ (_01585_, _01584_, _01582_);
  nand _34334_ (_01587_, _01585_, _01580_);
  not _34335_ (_01588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  not _34336_ (_01589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _34337_ (_01590_, _01589_, _01588_);
  not _34338_ (_01591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand _34339_ (_01592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _34340_ (_01593_, _01592_, _01591_);
  nand _34341_ (_01594_, _01593_, _01590_);
  nor _34342_ (_01595_, _01594_, _01587_);
  not _34343_ (_01597_, _01595_);
  nor _34344_ (_01598_, _01597_, _01575_);
  nor _34345_ (_01599_, _01595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _34346_ (_01601_, _01599_, _01598_);
  nand _34347_ (_01602_, _01601_, _01574_);
  not _34348_ (_01603_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _34349_ (_01604_, _01603_, _00166_);
  not _34350_ (_01605_, _01604_);
  nor _34351_ (_01606_, _01605_, _01575_);
  nand _34352_ (_01607_, _01605_, _01575_);
  not _34353_ (_01608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not _34354_ (_01609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _34355_ (_01611_, _01609_, _01608_);
  nand _34356_ (_01612_, _01611_, _01607_);
  nor _34357_ (_01613_, _01612_, _01606_);
  nor _34358_ (_01614_, _01609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor _34359_ (_01615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _01608_);
  nor _34360_ (_01616_, _01615_, _01614_);
  not _34361_ (_01617_, _01616_);
  not _34362_ (_01618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _34363_ (_01619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _34364_ (_01620_, _01594_, _01619_);
  nand _34365_ (_01621_, _01620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _34366_ (_01622_, _01621_, _01618_);
  nor _34367_ (_01624_, _01587_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand _34368_ (_01625_, _01624_, _01622_);
  nand _34369_ (_01626_, _01625_, _01575_);
  nand _34370_ (_01628_, _01626_, _01617_);
  not _34371_ (_01630_, _01622_);
  nor _34372_ (_01631_, _01630_, _01587_);
  not _34373_ (_01632_, _01631_);
  nor _34374_ (_01633_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _34375_ (_01634_, _01633_);
  nor _34376_ (_01635_, _01634_, _01575_);
  nor _34377_ (_01636_, _01635_, _01628_);
  nor _34378_ (_01637_, _01636_, _01613_);
  nand _34379_ (_01638_, _01637_, _01602_);
  nor _34380_ (_01639_, _24051_, _23938_);
  nand _34381_ (_01640_, _01639_, _00144_);
  nor _34382_ (_01641_, _01640_, _25627_);
  nand _34383_ (_01642_, _01641_, _25630_);
  nand _34384_ (_01643_, _01642_, _01638_);
  not _34385_ (_01644_, _01642_);
  nand _34386_ (_01645_, _01644_, _24821_);
  nand _34387_ (_01646_, _01645_, _01643_);
  nor _34388_ (_01647_, _01646_, _01573_);
  nand _34389_ (_01648_, _01573_, _01575_);
  nand _34390_ (_01649_, _01648_, _26487_);
  nor _34391_ (_23738_, _01649_, _01647_);
  nor _34392_ (_01650_, _01542_, _00147_);
  nand _34393_ (_01651_, _01650_, _24717_);
  nor _34394_ (_01652_, _01650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor _34395_ (_01653_, _01652_, _26245_);
  nand _34396_ (_01654_, _01653_, _01651_);
  nand _34397_ (_01655_, _01551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand _34398_ (_01657_, _01552_, _25028_);
  nand _34399_ (_01658_, _01657_, _01655_);
  nand _34400_ (_01659_, _01658_, _25630_);
  nand _34401_ (_01660_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand _34402_ (_01661_, _01660_, _01659_);
  nor _34403_ (_01662_, _01661_, rst);
  nand _34404_ (_23739_, _01662_, _01654_);
  nand _34405_ (_01663_, _01398_, _28096_);
  nand _34406_ (_01664_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  nand _34407_ (_23740_, _01664_, _01663_);
  nor _34408_ (_01665_, _26134_, _25721_);
  not _34409_ (_01666_, _01665_);
  nor _34410_ (_01667_, _01542_, _01666_);
  nand _34411_ (_01668_, _01667_, _24717_);
  nor _34412_ (_01669_, _01667_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _34413_ (_01670_, _01669_, _26245_);
  nand _34414_ (_01671_, _01670_, _01668_);
  nand _34415_ (_01672_, _01552_, _25140_);
  nor _34416_ (_01673_, _01552_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _34417_ (_01674_, _01673_, _25631_);
  nand _34418_ (_01675_, _01674_, _01672_);
  nand _34419_ (_01676_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nand _34420_ (_01677_, _01676_, _01675_);
  nor _34421_ (_01678_, _01677_, rst);
  nand _34422_ (_23741_, _01678_, _01671_);
  nor _34423_ (_01680_, _01542_, _00135_);
  nand _34424_ (_01681_, _01680_, _24717_);
  nor _34425_ (_01682_, _01680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor _34426_ (_01683_, _01682_, _26245_);
  nand _34427_ (_01684_, _01683_, _01681_);
  nand _34428_ (_01685_, _01552_, _26096_);
  nor _34429_ (_01686_, _01552_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor _34430_ (_01687_, _01686_, _25631_);
  nand _34431_ (_01688_, _01687_, _01685_);
  nand _34432_ (_01689_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand _34433_ (_01690_, _01689_, _01688_);
  nor _34434_ (_01691_, _01690_, rst);
  nand _34435_ (_23742_, _01691_, _01684_);
  nor _34436_ (_01692_, _01542_, _00263_);
  nand _34437_ (_01693_, _01692_, _24717_);
  nor _34438_ (_01694_, _01692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor _34439_ (_01695_, _01694_, _26245_);
  nand _34440_ (_01696_, _01695_, _01693_);
  nand _34441_ (_01697_, _01551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nand _34442_ (_01699_, _01552_, _25194_);
  nand _34443_ (_01700_, _01699_, _01697_);
  nand _34444_ (_01701_, _01700_, _25630_);
  nand _34445_ (_01702_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nand _34446_ (_01704_, _01702_, _01701_);
  nor _34447_ (_01705_, _01704_, rst);
  nand _34448_ (_23743_, _01705_, _01696_);
  nand _34449_ (_01706_, _01533_, _24927_);
  nand _34450_ (_01707_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  nand _34451_ (_23744_, _01707_, _01706_);
  nand _34452_ (_01709_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  nand _34453_ (_01710_, _01520_, _24789_);
  nand _34454_ (_23745_, _01710_, _01709_);
  nand _34455_ (_01711_, _01533_, _25039_);
  nand _34456_ (_01712_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nand _34457_ (_23746_, _01712_, _01711_);
  nor _34458_ (_01713_, _01540_, _26231_);
  not _34459_ (_01714_, _01713_);
  nor _34460_ (_01715_, _01714_, _00263_);
  nand _34461_ (_01716_, _01715_, _24717_);
  nor _34462_ (_01717_, _01715_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor _34463_ (_01718_, _01717_, _26245_);
  nand _34464_ (_01719_, _01718_, _01716_);
  nor _34465_ (_01720_, _00501_, _01549_);
  nand _34466_ (_01722_, _01720_, _25195_);
  nor _34467_ (_01723_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor _34468_ (_01724_, _01723_, _25631_);
  nand _34469_ (_01725_, _01724_, _01722_);
  nand _34470_ (_01726_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nand _34471_ (_01728_, _01726_, _01725_);
  nor _34472_ (_01729_, _01728_, rst);
  nand _34473_ (_23747_, _01729_, _01719_);
  nor _34474_ (_01730_, _01714_, _00276_);
  nand _34475_ (_01731_, _01730_, _24717_);
  nor _34476_ (_01732_, _01730_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor _34477_ (_01733_, _01732_, _26245_);
  nand _34478_ (_01734_, _01733_, _01731_);
  nand _34479_ (_01735_, _01720_, _25703_);
  nor _34480_ (_01737_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor _34481_ (_01738_, _01737_, _25631_);
  nand _34482_ (_01739_, _01738_, _01735_);
  nand _34483_ (_01740_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nand _34484_ (_01741_, _01740_, _01739_);
  nor _34485_ (_01742_, _01741_, rst);
  nand _34486_ (_23748_, _01742_, _01734_);
  nor _34487_ (_01743_, _01714_, _24842_);
  nand _34488_ (_01745_, _01743_, _24717_);
  nor _34489_ (_01746_, _01743_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor _34490_ (_01747_, _01746_, _26245_);
  nand _34491_ (_01748_, _01747_, _01745_);
  nand _34492_ (_01749_, _01720_, _25088_);
  nor _34493_ (_01750_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor _34494_ (_01751_, _01750_, _25631_);
  nand _34495_ (_01752_, _01751_, _01749_);
  nand _34496_ (_01753_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nand _34497_ (_01754_, _01753_, _01752_);
  nor _34498_ (_01756_, _01754_, rst);
  nand _34499_ (_23749_, _01756_, _01748_);
  nand _34500_ (_01757_, _01720_, _24717_);
  nor _34501_ (_01758_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _34502_ (_01759_, _01758_, _26245_);
  nand _34503_ (_01760_, _01759_, _01757_);
  nand _34504_ (_01761_, _01720_, _24820_);
  nand _34505_ (_01762_, _01761_, _25630_);
  nor _34506_ (_01763_, _01762_, _01758_);
  nand _34507_ (_01764_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nand _34508_ (_01765_, _01764_, _26487_);
  nor _34509_ (_01766_, _01765_, _01763_);
  nand _34510_ (_23750_, _01766_, _01760_);
  nand _34511_ (_01767_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nand _34512_ (_01768_, _01216_, _28096_);
  nand _34513_ (_23751_, _01768_, _01767_);
  nand _34514_ (_01769_, _00991_, _25150_);
  nand _34515_ (_01770_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  nand _34516_ (_23752_, _01770_, _01769_);
  nor _34517_ (_01771_, _01714_, _00135_);
  nand _34518_ (_01772_, _01771_, _24717_);
  nor _34519_ (_01773_, _01771_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor _34520_ (_01774_, _01773_, _26245_);
  nand _34521_ (_01775_, _01774_, _01772_);
  nand _34522_ (_01776_, _01720_, _26096_);
  nor _34523_ (_01777_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor _34524_ (_01778_, _01777_, _25631_);
  nand _34525_ (_01779_, _01778_, _01776_);
  nand _34526_ (_01780_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand _34527_ (_01781_, _01780_, _01779_);
  nor _34528_ (_01782_, _01781_, rst);
  nand _34529_ (_23754_, _01782_, _01775_);
  nand _34530_ (_01783_, _01533_, _24789_);
  nand _34531_ (_01785_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  nand _34532_ (_23755_, _01785_, _01783_);
  nand _34533_ (_01786_, _01402_, _25099_);
  nand _34534_ (_01787_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  nand _34535_ (_23756_, _01787_, _01786_);
  nor _34536_ (_01788_, _01714_, _01666_);
  nand _34537_ (_01789_, _01788_, _24717_);
  nor _34538_ (_01790_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor _34539_ (_01791_, _01790_, _26245_);
  nand _34540_ (_01792_, _01791_, _01789_);
  nand _34541_ (_01793_, _01720_, _25140_);
  nor _34542_ (_01794_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor _34543_ (_01795_, _01794_, _25631_);
  nand _34544_ (_01796_, _01795_, _01793_);
  nand _34545_ (_01797_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nand _34546_ (_01799_, _01797_, _01796_);
  nor _34547_ (_01800_, _01799_, rst);
  nand _34548_ (_23757_, _01800_, _01792_);
  nor _34549_ (_28207_[0], _25459_, rst);
  nor _34550_ (_28207_[1], _25266_, rst);
  nor _34551_ (_28207_[2], _25460_, rst);
  nor _34552_ (_28207_[3], _25743_, rst);
  nor _34553_ (_01801_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _34554_ (_01803_, _27586_, _25440_);
  nand _34555_ (_01804_, _01803_, _26487_);
  nor _34556_ (_28225_[0], _01804_, _01801_);
  nor _34557_ (_01806_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _34558_ (_01808_, _27586_, _25240_);
  nand _34559_ (_01809_, _01808_, _26487_);
  nor _34560_ (_28225_[1], _01809_, _01806_);
  nor _34561_ (_01810_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _34562_ (_01811_, _27586_, _25277_);
  nand _34563_ (_01812_, _01811_, _26487_);
  nor _34564_ (_28225_[2], _01812_, _01810_);
  nor _34565_ (_01813_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand _34566_ (_01814_, _27586_, _25220_);
  nand _34567_ (_01815_, _01814_, _26487_);
  nor _34568_ (_28225_[3], _01815_, _01813_);
  nor _34569_ (_01816_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand _34570_ (_01818_, _27586_, _25301_);
  nand _34571_ (_01819_, _01818_, _26487_);
  nor _34572_ (_28225_[4], _01819_, _01816_);
  nor _34573_ (_01820_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _34574_ (_01822_, _27586_, _25370_);
  nand _34575_ (_01823_, _01822_, _26487_);
  nor _34576_ (_28225_[5], _01823_, _01820_);
  nor _34577_ (_01824_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _34578_ (_01825_, _27586_, _24951_);
  nand _34579_ (_01826_, _01825_, _26487_);
  nor _34580_ (_28225_[6], _01826_, _01824_);
  nor _34581_ (_01827_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _34582_ (_01828_, _27586_, _25338_);
  nand _34583_ (_01829_, _01828_, _26487_);
  nor _34584_ (_28225_[7], _01829_, _01827_);
  nor _34585_ (_01830_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand _34586_ (_01831_, _27586_, _26325_);
  nand _34587_ (_01832_, _01831_, _26487_);
  nor _34588_ (_28225_[8], _01832_, _01830_);
  nor _34589_ (_01833_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand _34590_ (_01834_, _27586_, _25237_);
  nand _34591_ (_01835_, _01834_, _26487_);
  nor _34592_ (_28225_[9], _01835_, _01833_);
  nor _34593_ (_01836_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand _34594_ (_01837_, _27586_, _26379_);
  nand _34595_ (_01838_, _01837_, _26487_);
  nor _34596_ (_28225_[10], _01838_, _01836_);
  nor _34597_ (_01839_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _34598_ (_01840_, _27586_, _25208_);
  nand _34599_ (_01841_, _01840_, _26487_);
  nor _34600_ (_28225_[11], _01841_, _01839_);
  nor _34601_ (_01842_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand _34602_ (_01843_, _27586_, _25299_);
  nand _34603_ (_01844_, _01843_, _26487_);
  nor _34604_ (_28225_[12], _01844_, _01842_);
  nor _34605_ (_01845_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand _34606_ (_01846_, _27586_, _26110_);
  nand _34607_ (_01848_, _01846_, _26487_);
  nor _34608_ (_28225_[13], _01848_, _01845_);
  nor _34609_ (_01849_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand _34610_ (_01850_, _27586_, _24945_);
  nand _34611_ (_01851_, _01850_, _26487_);
  nor _34612_ (_28225_[14], _01851_, _01849_);
  nor _34613_ (_01852_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _34614_ (_01853_, _27586_, _25336_);
  nand _34615_ (_01854_, _01853_, _26487_);
  nor _34616_ (_28225_[15], _01854_, _01852_);
  nor _34617_ (_01855_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  nand _34618_ (_01856_, _27586_, _26319_);
  nand _34619_ (_01857_, _01856_, _26487_);
  nor _34620_ (_28225_[16], _01857_, _01855_);
  nor _34621_ (_01858_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  nand _34622_ (_01859_, _27586_, _26416_);
  nand _34623_ (_01860_, _01859_, _26487_);
  nor _34624_ (_28225_[17], _01860_, _01858_);
  nor _34625_ (_01861_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  nand _34626_ (_01862_, _27586_, _26374_);
  nand _34627_ (_01863_, _01862_, _26487_);
  nor _34628_ (_28225_[18], _01863_, _01861_);
  nor _34629_ (_01864_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  nand _34630_ (_01865_, _27586_, _25901_);
  nand _34631_ (_01866_, _01865_, _26487_);
  nor _34632_ (_28225_[19], _01866_, _01864_);
  nor _34633_ (_01867_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  nand _34634_ (_01868_, _27586_, _26002_);
  nand _34635_ (_01869_, _01868_, _26487_);
  nor _34636_ (_28225_[20], _01869_, _01867_);
  nor _34637_ (_01870_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  nand _34638_ (_01871_, _27586_, _26106_);
  nand _34639_ (_01873_, _01871_, _26487_);
  nor _34640_ (_28225_[21], _01873_, _01870_);
  nor _34641_ (_01874_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  nand _34642_ (_01875_, _27586_, _25975_);
  nand _34643_ (_01877_, _01875_, _26487_);
  nor _34644_ (_28225_[22], _01877_, _01874_);
  nor _34645_ (_01878_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  nand _34646_ (_01879_, _27586_, _25825_);
  nand _34647_ (_01880_, _01879_, _26487_);
  nor _34648_ (_28225_[23], _01880_, _01878_);
  nor _34649_ (_01881_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  nand _34650_ (_01882_, _27586_, _26705_);
  nand _34651_ (_01883_, _01882_, _26487_);
  nor _34652_ (_28225_[24], _01883_, _01881_);
  nor _34653_ (_01884_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  nand _34654_ (_01885_, _27586_, _26679_);
  nand _34655_ (_01887_, _01885_, _26487_);
  nor _34656_ (_28225_[25], _01887_, _01884_);
  nor _34657_ (_01888_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  nand _34658_ (_01889_, _27586_, _26658_);
  nand _34659_ (_01890_, _01889_, _26487_);
  nor _34660_ (_28225_[26], _01890_, _01888_);
  nor _34661_ (_01892_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  nand _34662_ (_01893_, _27586_, _26620_);
  nand _34663_ (_01894_, _01893_, _26487_);
  nor _34664_ (_28225_[27], _01894_, _01892_);
  nor _34665_ (_01895_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand _34666_ (_01896_, _27586_, _26591_);
  nand _34667_ (_01898_, _01896_, _26487_);
  nor _34668_ (_28225_[28], _01898_, _01895_);
  nor _34669_ (_01899_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  nand _34670_ (_01900_, _27586_, _26572_);
  nand _34671_ (_01901_, _01900_, _26487_);
  nor _34672_ (_28225_[29], _01901_, _01899_);
  nor _34673_ (_01902_, _27586_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  nand _34674_ (_01903_, _27586_, _26537_);
  nand _34675_ (_01904_, _01903_, _26487_);
  nor _34676_ (_28225_[30], _01904_, _01902_);
  nor _34677_ (_28208_[0], _26309_, rst);
  nor _34678_ (_28208_[1], _26469_, rst);
  nor _34679_ (_28208_[2], _26366_, rst);
  nor _34680_ (_28208_[3], _25881_, rst);
  nor _34681_ (_28208_[4], _26044_, rst);
  nor _34682_ (_28208_[5], _26098_, rst);
  nor _34683_ (_28208_[6], _25965_, rst);
  nor _34684_ (_01905_, _25159_, _24882_);
  nand _34685_ (_01906_, _01905_, _25203_);
  not _34686_ (_01907_, _01905_);
  nand _34687_ (_01908_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nand _34688_ (_23758_, _01908_, _01906_);
  nand _34689_ (_01909_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  nand _34690_ (_01910_, _01520_, _25099_);
  nand _34691_ (_23759_, _01910_, _01909_);
  nand _34692_ (_01911_, _01905_, _28096_);
  nand _34693_ (_01912_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nand _34694_ (_23760_, _01912_, _01911_);
  nand _34695_ (_01913_, _26255_, _00616_);
  nor _34696_ (_01914_, _01913_, _24842_);
  nand _34697_ (_01915_, _01914_, _24717_);
  nor _34698_ (_01916_, _01914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor _34699_ (_01917_, _01916_, _26245_);
  nand _34700_ (_01918_, _01917_, _01915_);
  nor _34701_ (_01919_, _01286_, _01549_);
  nand _34702_ (_01920_, _01919_, _25088_);
  nor _34703_ (_01921_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor _34704_ (_01922_, _01921_, _25631_);
  nand _34705_ (_01923_, _01922_, _01920_);
  nand _34706_ (_01924_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nand _34707_ (_01925_, _01924_, _01923_);
  nor _34708_ (_01926_, _01925_, rst);
  nand _34709_ (_23761_, _01926_, _01918_);
  nor _34710_ (_01927_, _01913_, _25723_);
  nand _34711_ (_01928_, _01927_, _24717_);
  nor _34712_ (_01929_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _34713_ (_01930_, _01929_, _26245_);
  nand _34714_ (_01931_, _01930_, _01928_);
  nand _34715_ (_01932_, _01919_, _24820_);
  nand _34716_ (_01933_, _01932_, _25630_);
  nor _34717_ (_01934_, _01933_, _01929_);
  nand _34718_ (_01935_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nand _34719_ (_01936_, _01935_, _26487_);
  nor _34720_ (_01937_, _01936_, _01934_);
  nand _34721_ (_23762_, _01937_, _01931_);
  nand _34722_ (_01938_, _01905_, _25099_);
  nand _34723_ (_01939_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand _34724_ (_23763_, _01939_, _01938_);
  nand _34725_ (_01940_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  nand _34726_ (_01941_, _01520_, _24830_);
  nand _34727_ (_23764_, _01941_, _01940_);
  nand _34728_ (_01942_, _27076_, _27027_);
  nor _34729_ (_01943_, _27027_, _27010_);
  not _34730_ (_01944_, _27027_);
  nor _34731_ (_01945_, _01944_, _26888_);
  nor _34732_ (_01946_, _01945_, _01943_);
  nand _34733_ (_01947_, _27056_, _01946_);
  nand _34734_ (_01948_, _01947_, _01942_);
  nand _34735_ (_01949_, _01948_, _24767_);
  nor _34736_ (_01950_, _27386_, _27382_);
  nor _34737_ (_01951_, _27408_, _27406_);
  nor _34738_ (_01952_, _01951_, _01950_);
  not _34739_ (_01953_, _01952_);
  nor _34740_ (_01954_, _01953_, _27506_);
  nor _34741_ (_01955_, _24590_, _24088_);
  nor _34742_ (_01956_, _01955_, _26172_);
  nor _34743_ (_01957_, _24700_, _24498_);
  nand _34744_ (_01958_, _24773_, _24380_);
  nand _34745_ (_01959_, _24686_, _24575_);
  not _34746_ (_01960_, _01959_);
  nor _34747_ (_01961_, _24668_, _24650_);
  nor _34748_ (_01962_, _01961_, _24428_);
  nor _34749_ (_01963_, _01962_, _01960_);
  nand _34750_ (_01964_, _01963_, _01958_);
  nor _34751_ (_01965_, _01964_, _24816_);
  nand _34752_ (_01966_, _01965_, _24811_);
  nor _34753_ (_01967_, _01966_, _24808_);
  not _34754_ (_01968_, _01967_);
  nor _34755_ (_01969_, _01968_, _01957_);
  not _34756_ (_01970_, _01969_);
  nor _34757_ (_01971_, _01970_, _01956_);
  not _34758_ (_01972_, _01971_);
  nor _34759_ (_01973_, _01972_, _01954_);
  nand _34760_ (_01974_, _01973_, _01949_);
  not _34761_ (_01975_, _26794_);
  nand _34762_ (_01976_, _26798_, _01975_);
  nor _34763_ (_01977_, _01976_, _26526_);
  nor _34764_ (_01978_, _01977_, _26797_);
  not _34765_ (_01979_, _01978_);
  nand _34766_ (_01980_, _01979_, _01974_);
  nor _34767_ (_01981_, _25614_, _27629_);
  nand _34768_ (_01982_, _26722_, _27566_);
  nand _34769_ (_01983_, _26799_, _01975_);
  not _34770_ (_01984_, _01983_);
  nand _34771_ (_01985_, _01984_, _26724_);
  nand _34772_ (_01986_, _01985_, _01982_);
  nor _34773_ (_01987_, _01986_, _01981_);
  nand _34774_ (_01988_, _01987_, _01980_);
  nor _34775_ (_01989_, _26726_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _34776_ (_01990_, _01989_, _26728_);
  nand _34777_ (_01991_, _01990_, _26800_);
  nand _34778_ (_01992_, _01991_, _26485_);
  nor _34779_ (_01993_, _01992_, _01988_);
  nand _34780_ (_01994_, _26486_, _27629_);
  nand _34781_ (_01995_, _01994_, _26487_);
  nor _34782_ (_28211_[0], _01995_, _01993_);
  nor _34783_ (_01996_, _01950_, _27402_);
  nor _34784_ (_01997_, _01996_, _27299_);
  not _34785_ (_01998_, _01996_);
  nor _34786_ (_01999_, _01998_, _27401_);
  nor _34787_ (_02000_, _01999_, _01997_);
  nand _34788_ (_02001_, _02000_, _24770_);
  not _34789_ (_02002_, _02001_);
  nor _34790_ (_02003_, _27029_, _27024_);
  nor _34791_ (_02004_, _02003_, _27063_);
  nor _34792_ (_02005_, _02004_, _27076_);
  nor _34793_ (_02006_, _27056_, _27016_);
  nor _34794_ (_02007_, _02006_, _02005_);
  nand _34795_ (_02008_, _02007_, _24767_);
  nor _34796_ (_02009_, _24441_, _24435_);
  nor _34797_ (_02010_, _02009_, _24443_);
  nor _34798_ (_02011_, _02010_, _24512_);
  nor _34799_ (_02012_, _24514_, _24089_);
  not _34800_ (_02013_, _02012_);
  nor _34801_ (_02014_, _02013_, _02011_);
  nand _34802_ (_02015_, _24629_, _24627_);
  nand _34803_ (_02016_, _02015_, _24631_);
  nand _34804_ (_02017_, _02016_, _24590_);
  not _34805_ (_02018_, _02017_);
  nor _34806_ (_02019_, _02018_, _02014_);
  not _34807_ (_02020_, _02019_);
  not _34808_ (_02021_, _25074_);
  nor _34809_ (_02022_, _24657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  not _34810_ (_02023_, _02022_);
  nor _34811_ (_02024_, _02023_, _24381_);
  nor _34812_ (_02025_, _02022_, _24380_);
  nor _34813_ (_02026_, _02025_, _02024_);
  nor _34814_ (_02027_, _02026_, _24651_);
  nor _34815_ (_02028_, _27447_, _24381_);
  not _34816_ (_02029_, _24775_);
  nor _34817_ (_02030_, _02029_, _24428_);
  nand _34818_ (_02031_, _24773_, _24350_);
  not _34819_ (_02032_, _02031_);
  nor _34820_ (_02033_, _02032_, _02030_);
  not _34821_ (_02034_, _02033_);
  nor _34822_ (_02035_, _02034_, _02028_);
  nand _34823_ (_02036_, _02035_, _25086_);
  nor _34824_ (_02037_, _02036_, _02027_);
  nand _34825_ (_02038_, _02037_, _02021_);
  nor _34826_ (_02039_, _02038_, _02020_);
  nand _34827_ (_02040_, _02039_, _02008_);
  nor _34828_ (_02041_, _02040_, _02002_);
  nor _34829_ (_02042_, _02041_, _01978_);
  nand _34830_ (_02043_, _25613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _34831_ (_02044_, _26733_, _26728_);
  nand _34832_ (_02045_, _26800_, _26734_);
  nor _34833_ (_02046_, _02045_, _02044_);
  nand _34834_ (_02047_, _26696_, _27566_);
  not _34835_ (_02048_, _26426_);
  nand _34836_ (_02049_, _01984_, _02048_);
  nand _34837_ (_02050_, _02049_, _02047_);
  nor _34838_ (_02051_, _02050_, _02046_);
  nand _34839_ (_02052_, _02051_, _02043_);
  nor _34840_ (_02053_, _02052_, _02042_);
  nor _34841_ (_02054_, _02053_, _26486_);
  nor _34842_ (_02055_, _26485_, _27626_);
  nor _34843_ (_02056_, _02055_, _02054_);
  nor _34844_ (_28211_[1], _02056_, rst);
  nor _34845_ (_02057_, _27042_, _27031_);
  nor _34846_ (_02058_, _02057_, _27067_);
  nor _34847_ (_02059_, _02058_, _27076_);
  nor _34848_ (_02060_, _27056_, _27038_);
  nor _34849_ (_02061_, _02060_, _02059_);
  nand _34850_ (_02062_, _02061_, _24767_);
  nor _34851_ (_02063_, _01997_, _27269_);
  nor _34852_ (_02064_, _02063_, _27307_);
  not _34853_ (_02065_, _02064_);
  nand _34854_ (_02066_, _02063_, _27307_);
  nand _34855_ (_02067_, _02066_, _02065_);
  nor _34856_ (_02068_, _02067_, _27506_);
  not _34857_ (_02069_, _24518_);
  nor _34858_ (_02070_, _24517_, _24514_);
  not _34859_ (_02071_, _02070_);
  nand _34860_ (_02072_, _02071_, _24088_);
  nor _34861_ (_02073_, _02072_, _02069_);
  nand _34862_ (_02074_, _24631_, _24624_);
  nand _34863_ (_02075_, _02074_, _24633_);
  nand _34864_ (_02076_, _02075_, _24590_);
  nor _34865_ (_02077_, _02025_, _24323_);
  not _34866_ (_02078_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  not _34867_ (_02079_, _24656_);
  nor _34868_ (_02080_, _02079_, _02078_);
  nor _34869_ (_02081_, _02080_, _02077_);
  nor _34870_ (_02082_, _02081_, _24651_);
  nor _34871_ (_02083_, _27447_, _24323_);
  nand _34872_ (_02084_, _24775_, _24380_);
  nand _34873_ (_02085_, _24773_, _24278_);
  nand _34874_ (_02086_, _02085_, _02084_);
  nor _34875_ (_02087_, _02086_, _02083_);
  not _34876_ (_02088_, _02087_);
  nor _34877_ (_02089_, _02088_, _25677_);
  not _34878_ (_02090_, _02089_);
  nor _34879_ (_02091_, _02090_, _02082_);
  nand _34880_ (_02092_, _02091_, _02076_);
  nor _34881_ (_02093_, _02092_, _02073_);
  nand _34882_ (_02094_, _02093_, _25669_);
  nor _34883_ (_02095_, _02094_, _02068_);
  nand _34884_ (_02096_, _02095_, _02062_);
  nand _34885_ (_02097_, _02096_, _01979_);
  nor _34886_ (_02098_, _01983_, _26385_);
  nand _34887_ (_02099_, _25613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nand _34888_ (_02100_, _26668_, _27566_);
  nand _34889_ (_02101_, _02100_, _02099_);
  nor _34890_ (_02102_, _02101_, _02098_);
  nand _34891_ (_02103_, _02102_, _02097_);
  nor _34892_ (_02104_, _26737_, _26735_);
  nor _34893_ (_02105_, _02104_, _26764_);
  nand _34894_ (_02106_, _02105_, _26800_);
  nand _34895_ (_02107_, _02106_, _26485_);
  nor _34896_ (_02108_, _02107_, _02103_);
  nor _34897_ (_02109_, _27586_, _27594_);
  not _34898_ (_02110_, _27586_);
  nor _34899_ (_02111_, _02110_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _34900_ (_02112_, _02111_, _02109_);
  not _34901_ (_02113_, _02112_);
  nand _34902_ (_02114_, _02113_, _26486_);
  nand _34903_ (_02115_, _02114_, _26487_);
  nor _34904_ (_28211_[2], _02115_, _02108_);
  nor _34905_ (_02116_, _27056_, _27044_);
  not _34906_ (_02117_, _27045_);
  nand _34907_ (_02118_, _02117_, _27008_);
  not _34908_ (_02119_, _02118_);
  nor _34909_ (_02120_, _27067_, _27040_);
  nand _34910_ (_02122_, _02120_, _02119_);
  not _34911_ (_02123_, _02122_);
  nor _34912_ (_02124_, _02120_, _02119_);
  nor _34913_ (_02125_, _02124_, _02123_);
  nor _34914_ (_02127_, _02125_, _27076_);
  nor _34915_ (_02128_, _02127_, _02116_);
  nor _34916_ (_02129_, _02128_, _24768_);
  not _34917_ (_02130_, _27308_);
  nor _34918_ (_02131_, _02130_, _02064_);
  nor _34919_ (_02132_, _02131_, _27412_);
  nand _34920_ (_02133_, _02132_, _24770_);
  nor _34921_ (_02134_, _26168_, _24591_);
  not _34922_ (_02135_, _24450_);
  nor _34923_ (_02136_, _02069_, _02135_);
  nor _34924_ (_02137_, _24519_, _24089_);
  not _34925_ (_02138_, _02137_);
  nor _34926_ (_02139_, _02138_, _02136_);
  nor _34927_ (_02141_, _24656_, _02078_);
  nor _34928_ (_02142_, _02141_, _24278_);
  nor _34929_ (_02143_, _02142_, _24651_);
  nand _34930_ (_02145_, _02143_, _27426_);
  nor _34931_ (_02146_, _27447_, _24279_);
  nand _34932_ (_02147_, _24773_, _24243_);
  nand _34933_ (_02149_, _24775_, _24350_);
  nand _34934_ (_02150_, _02149_, _02147_);
  nor _34935_ (_02151_, _02150_, _02146_);
  nand _34936_ (_02152_, _02151_, _25179_);
  nor _34937_ (_02153_, _02152_, _25192_);
  nand _34938_ (_02154_, _02153_, _02145_);
  nor _34939_ (_02155_, _02154_, _02139_);
  not _34940_ (_02156_, _02155_);
  nor _34941_ (_02158_, _02156_, _02134_);
  nand _34942_ (_02159_, _02158_, _02133_);
  nor _34943_ (_02160_, _02159_, _02129_);
  nor _34944_ (_02161_, _02160_, _01978_);
  nand _34945_ (_02162_, _26647_, _26645_);
  not _34946_ (_02163_, _02162_);
  nand _34947_ (_02164_, _02163_, _26765_);
  nand _34948_ (_02165_, _02162_, _26739_);
  nand _34949_ (_02166_, _02165_, _02164_);
  nand _34950_ (_02167_, _02166_, _26800_);
  nor _34951_ (_02168_, _25614_, _27590_);
  nand _34952_ (_02169_, _26638_, _27566_);
  nand _34953_ (_02170_, _01984_, _26640_);
  nand _34954_ (_02172_, _02170_, _02169_);
  nor _34955_ (_02173_, _02172_, _02168_);
  nand _34956_ (_02174_, _02173_, _02167_);
  nor _34957_ (_02176_, _02174_, _02161_);
  nor _34958_ (_02177_, _02176_, _26486_);
  not _34959_ (_02178_, _02109_);
  nor _34960_ (_02179_, _02178_, _27590_);
  nor _34961_ (_02181_, _02109_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _34962_ (_02182_, _02181_, _02179_);
  not _34963_ (_02183_, _02182_);
  nor _34964_ (_02184_, _02183_, _26485_);
  nor _34965_ (_02185_, _02184_, _02177_);
  nor _34966_ (_28211_[3], _02185_, rst);
  nand _34967_ (_02186_, _27050_, _27070_);
  not _34968_ (_02187_, _27050_);
  nand _34969_ (_02188_, _02187_, _27048_);
  nand _34970_ (_02189_, _02188_, _02186_);
  nand _34971_ (_02190_, _02189_, _27056_);
  not _34972_ (_02191_, _26991_);
  nand _34973_ (_02192_, _27076_, _02191_);
  nand _34974_ (_02194_, _02192_, _02190_);
  nor _34975_ (_02195_, _02194_, _24768_);
  nor _34976_ (_02196_, _27391_, _27390_);
  not _34977_ (_02197_, _27391_);
  nor _34978_ (_02199_, _02197_, _27412_);
  nor _34979_ (_02200_, _02199_, _02196_);
  nand _34980_ (_02201_, _02200_, _24770_);
  nor _34981_ (_02202_, _26165_, _24591_);
  not _34982_ (_02203_, _24523_);
  nor _34983_ (_02204_, _02203_, _24249_);
  nor _34984_ (_02205_, _24524_, _24089_);
  not _34985_ (_02206_, _02205_);
  nor _34986_ (_02207_, _02206_, _02204_);
  nor _34987_ (_02208_, _27427_, _24243_);
  not _34988_ (_02210_, _02208_);
  nand _34989_ (_02211_, _02210_, _24650_);
  nor _34990_ (_02212_, _02211_, _27433_);
  nand _34991_ (_02213_, _24773_, _24196_);
  nor _34992_ (_02214_, _27447_, _24224_);
  nand _34993_ (_02215_, _24775_, _24278_);
  not _34994_ (_02216_, _02215_);
  nor _34995_ (_02217_, _02216_, _02214_);
  nand _34996_ (_02218_, _02217_, _02213_);
  nor _34997_ (_02219_, _02218_, _25025_);
  not _34998_ (_02220_, _02219_);
  nor _34999_ (_02221_, _02220_, _02212_);
  nand _35000_ (_02222_, _02221_, _25017_);
  nor _35001_ (_02224_, _02222_, _02207_);
  not _35002_ (_02225_, _02224_);
  nor _35003_ (_02226_, _02225_, _02202_);
  nand _35004_ (_02228_, _02226_, _02201_);
  nor _35005_ (_02229_, _02228_, _02195_);
  nor _35006_ (_02230_, _02229_, _01978_);
  nand _35007_ (_02231_, _26768_, _26767_);
  nor _35008_ (_02232_, _26801_, _26769_);
  nand _35009_ (_02233_, _02232_, _02231_);
  nor _35010_ (_02234_, _25614_, _27591_);
  nand _35011_ (_02235_, _26608_, _27566_);
  nand _35012_ (_02236_, _01984_, _26610_);
  nand _35013_ (_02238_, _02236_, _02235_);
  nor _35014_ (_02239_, _02238_, _02234_);
  nand _35015_ (_02240_, _02239_, _02233_);
  nor _35016_ (_02241_, _02240_, _02230_);
  nor _35017_ (_02242_, _02241_, _26486_);
  not _35018_ (_02243_, _27592_);
  nor _35019_ (_02244_, _02243_, _02178_);
  not _35020_ (_02245_, _02244_);
  not _35021_ (_02246_, _02179_);
  nand _35022_ (_02248_, _02246_, _27591_);
  nand _35023_ (_02249_, _02248_, _02245_);
  nor _35024_ (_02251_, _02249_, _26485_);
  nor _35025_ (_02252_, _02251_, _02242_);
  nor _35026_ (_28211_[4], _02252_, rst);
  nor _35027_ (_02254_, _27056_, _26981_);
  not _35028_ (_02255_, _26995_);
  nand _35029_ (_02257_, _02186_, _26992_);
  nor _35030_ (_02258_, _02257_, _02255_);
  nor _35031_ (_02259_, _02187_, _27048_);
  nor _35032_ (_02261_, _02259_, _26993_);
  nor _35033_ (_02262_, _02261_, _26995_);
  nor _35034_ (_02263_, _02262_, _02258_);
  nor _35035_ (_02264_, _02263_, _27076_);
  nor _35036_ (_02265_, _02264_, _02254_);
  nor _35037_ (_02266_, _02265_, _24768_);
  not _35038_ (_02267_, _27392_);
  nor _35039_ (_02268_, _02267_, _02196_);
  nor _35040_ (_02269_, _02268_, _27395_);
  nand _35041_ (_02270_, _02269_, _24770_);
  nor _35042_ (_02271_, _24242_, _24201_);
  nor _35043_ (_02272_, _02271_, _24564_);
  nor _35044_ (_02273_, _02272_, _24524_);
  not _35045_ (_02274_, _24525_);
  nor _35046_ (_02276_, _02274_, _24089_);
  not _35047_ (_02277_, _02276_);
  nor _35048_ (_02278_, _02277_, _02273_);
  nand _35049_ (_02279_, _26160_, _24590_);
  not _35050_ (_02280_, _02279_);
  not _35051_ (_02281_, _27431_);
  nor _35052_ (_02282_, _27433_, _24196_);
  nor _35053_ (_02283_, _27434_, _24179_);
  nor _35054_ (_02285_, _02283_, _02282_);
  not _35055_ (_02286_, _02285_);
  nor _35056_ (_02287_, _02286_, _02281_);
  nor _35057_ (_02288_, _02285_, _27431_);
  nor _35058_ (_02289_, _02288_, _02287_);
  nor _35059_ (_02290_, _02289_, _24651_);
  nor _35060_ (_02291_, _27447_, _24179_);
  nand _35061_ (_02292_, _24775_, _24243_);
  nand _35062_ (_02293_, _24773_, _24557_);
  nand _35063_ (_02294_, _02293_, _02292_);
  nor _35064_ (_02295_, _02294_, _02291_);
  not _35065_ (_02296_, _02295_);
  nor _35066_ (_02297_, _02296_, _24917_);
  not _35067_ (_02299_, _02297_);
  nor _35068_ (_02300_, _02299_, _02290_);
  nand _35069_ (_02301_, _02300_, _24908_);
  nor _35070_ (_02302_, _02301_, _02280_);
  not _35071_ (_02303_, _02302_);
  nor _35072_ (_02304_, _02303_, _02278_);
  nand _35073_ (_02305_, _02304_, _02270_);
  nor _35074_ (_02307_, _02305_, _02266_);
  nor _35075_ (_02308_, _02307_, _01978_);
  nand _35076_ (_02309_, _26587_, _26586_);
  not _35077_ (_02311_, _02309_);
  nor _35078_ (_02312_, _02311_, _26770_);
  nor _35079_ (_02313_, _02309_, _26745_);
  nor _35080_ (_02314_, _02313_, _02312_);
  nor _35081_ (_02316_, _02314_, _26801_);
  nand _35082_ (_02317_, _25613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _35083_ (_02318_, _26581_, _26495_);
  nor _35084_ (_02319_, _01983_, _26118_);
  nor _35085_ (_02320_, _02319_, _02318_);
  nand _35086_ (_02321_, _02320_, _02317_);
  nor _35087_ (_02322_, _02321_, _02316_);
  nand _35088_ (_02323_, _02322_, _26485_);
  nor _35089_ (_02324_, _02323_, _02308_);
  nand _35090_ (_02325_, _02244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nand _35091_ (_02326_, _02245_, _27595_);
  nand _35092_ (_02327_, _02326_, _02325_);
  nand _35093_ (_02328_, _02327_, _26486_);
  nand _35094_ (_02329_, _02328_, _26487_);
  nor _35095_ (_28211_[5], _02329_, _02324_);
  nor _35096_ (_02330_, _26158_, _24591_);
  not _35097_ (_02331_, _02330_);
  nand _35098_ (_02332_, _27053_, _26968_);
  nand _35099_ (_02333_, _02332_, _27078_);
  nand _35100_ (_02334_, _02333_, _27056_);
  nand _35101_ (_02335_, _27076_, _26960_);
  nand _35102_ (_02336_, _02335_, _02334_);
  nor _35103_ (_02337_, _02336_, _24768_);
  nand _35104_ (_02338_, _27413_, _27091_);
  nor _35105_ (_02339_, _27414_, _27506_);
  nand _35106_ (_02341_, _02339_, _02338_);
  not _35107_ (_02342_, _24569_);
  nor _35108_ (_02343_, _02342_, _02274_);
  nor _35109_ (_02344_, _24570_, _24089_);
  not _35110_ (_02346_, _02344_);
  nor _35111_ (_02347_, _02346_, _02343_);
  nand _35112_ (_02348_, _02282_, _02281_);
  not _35113_ (_02350_, _02348_);
  nor _35114_ (_02351_, _02350_, _24557_);
  nor _35115_ (_02352_, _02348_, _24549_);
  nor _35116_ (_02353_, _02352_, _24651_);
  not _35117_ (_02354_, _02353_);
  nor _35118_ (_02355_, _02354_, _02351_);
  nand _35119_ (_02356_, _24775_, _24196_);
  nand _35120_ (_02357_, _24773_, _24575_);
  not _35121_ (_02358_, _02357_);
  nor _35122_ (_02360_, _27447_, _24549_);
  nor _35123_ (_02361_, _02360_, _02358_);
  nand _35124_ (_02362_, _02361_, _02356_);
  nor _35125_ (_02364_, _02362_, _25136_);
  nand _35126_ (_02365_, _02364_, _25128_);
  nor _35127_ (_02366_, _02365_, _02355_);
  not _35128_ (_02367_, _02366_);
  nor _35129_ (_02369_, _02367_, _02347_);
  nand _35130_ (_02370_, _02369_, _02341_);
  nor _35131_ (_02372_, _02370_, _02337_);
  nand _35132_ (_02373_, _02372_, _02331_);
  nand _35133_ (_02374_, _02373_, _01979_);
  nor _35134_ (_02375_, _26747_, _26561_);
  nand _35135_ (_02376_, _26800_, _26748_);
  nor _35136_ (_02377_, _02376_, _02375_);
  nand _35137_ (_02378_, _25613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _35138_ (_02379_, _26553_, _26495_);
  nor _35139_ (_02380_, _01983_, _25985_);
  nor _35140_ (_02381_, _02380_, _02379_);
  nand _35141_ (_02382_, _02381_, _02378_);
  nor _35142_ (_02383_, _02382_, _02377_);
  nand _35143_ (_02384_, _02383_, _02374_);
  nor _35144_ (_02385_, _02384_, _26486_);
  nor _35145_ (_02386_, _27599_, _27586_);
  not _35146_ (_02387_, _02386_);
  nand _35147_ (_02388_, _02325_, _27589_);
  nand _35148_ (_02389_, _02388_, _02387_);
  nand _35149_ (_02390_, _02389_, _26486_);
  nand _35150_ (_02392_, _02390_, _26487_);
  nor _35151_ (_28211_[6], _02392_, _02385_);
  nand _35152_ (_02393_, _26531_, _26533_);
  nor _35153_ (_02394_, _02393_, _26774_);
  nand _35154_ (_02396_, _02393_, _26774_);
  nand _35155_ (_02397_, _02396_, _26800_);
  nor _35156_ (_02398_, _02397_, _02394_);
  nand _35157_ (_02399_, _27076_, _26951_);
  nand _35158_ (_02401_, _27082_, _26964_);
  nand _35159_ (_02402_, _27079_, _26965_);
  nand _35160_ (_02403_, _02402_, _02401_);
  nand _35161_ (_02404_, _02403_, _27056_);
  nand _35162_ (_02406_, _02404_, _02399_);
  nand _35163_ (_02407_, _02406_, _24767_);
  not _35164_ (_02408_, _27398_);
  nor _35165_ (_02409_, _02408_, _27414_);
  nor _35166_ (_02410_, _27396_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _35167_ (_02411_, _02410_, _02409_);
  nor _35168_ (_02412_, _02411_, _27506_);
  not _35169_ (_02413_, _27458_);
  nor _35170_ (_02414_, _02413_, _02412_);
  nand _35171_ (_02415_, _02414_, _02407_);
  nand _35172_ (_02416_, _01979_, _02415_);
  nor _35173_ (_02417_, _01983_, _25837_);
  nand _35174_ (_02419_, _26524_, _27566_);
  nand _35175_ (_02420_, _25613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nand _35176_ (_02421_, _02420_, _02419_);
  nor _35177_ (_02422_, _02421_, _02417_);
  nand _35178_ (_02424_, _02422_, _02416_);
  nor _35179_ (_02425_, _02424_, _02398_);
  nor _35180_ (_02426_, _02425_, _26486_);
  nand _35181_ (_02428_, _02386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nand _35182_ (_02429_, _02387_, _27587_);
  nand _35183_ (_02431_, _02429_, _02428_);
  nor _35184_ (_02432_, _02431_, _26485_);
  nor _35185_ (_02433_, _02432_, _02426_);
  nor _35186_ (_28211_[7], _02433_, rst);
  nand _35187_ (_02434_, _26751_, _24398_);
  nand _35188_ (_02435_, _26776_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand _35189_ (_02436_, _02435_, _02434_);
  nand _35190_ (_02437_, _02436_, _26528_);
  nor _35191_ (_02438_, _02436_, _26528_);
  nor _35192_ (_02439_, _02438_, _26801_);
  nand _35193_ (_02441_, _02439_, _02437_);
  nor _35194_ (_02442_, _27056_, _01944_);
  not _35195_ (_02443_, _01946_);
  nor _35196_ (_02444_, _27076_, _02443_);
  nor _35197_ (_02445_, _02444_, _02442_);
  nor _35198_ (_02446_, _02445_, _24768_);
  not _35199_ (_02447_, _01973_);
  nor _35200_ (_02448_, _02447_, _02446_);
  nor _35201_ (_02450_, _02448_, _25614_);
  nand _35202_ (_02451_, _01984_, _25383_);
  not _35203_ (_02452_, _26797_);
  nor _35204_ (_02453_, _27474_, _27471_);
  not _35205_ (_02454_, _02453_);
  nand _35206_ (_02455_, _02454_, _27476_);
  nor _35207_ (_02456_, _02455_, _24089_);
  nand _35208_ (_02457_, _27056_, _24767_);
  nor _35209_ (_02458_, _24752_, _27552_);
  nand _35210_ (_02459_, _02458_, _24740_);
  not _35211_ (_02460_, _02459_);
  nor _35212_ (_02461_, _02460_, _24508_);
  nor _35213_ (_02462_, _02459_, _24434_);
  nor _35214_ (_02463_, _02462_, _24743_);
  not _35215_ (_02464_, _02463_);
  nor _35216_ (_02465_, _02464_, _02461_);
  nor _35217_ (_02467_, _27447_, _24434_);
  nor _35218_ (_02468_, _27272_, _27506_);
  not _35219_ (_02469_, _02468_);
  nor _35220_ (_02470_, _24700_, _24224_);
  nor _35221_ (_02471_, _24751_, _24428_);
  nor _35222_ (_02472_, _02471_, _02470_);
  nand _35223_ (_02473_, _02472_, _02469_);
  nor _35224_ (_02474_, _02473_, _02467_);
  not _35225_ (_02475_, _02474_);
  nor _35226_ (_02476_, _02475_, _02465_);
  nand _35227_ (_02477_, _02476_, _02457_);
  nor _35228_ (_02478_, _02477_, _02456_);
  nor _35229_ (_02479_, _02478_, _02452_);
  nand _35230_ (_02480_, _27566_, _26724_);
  nand _35231_ (_02481_, _01977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand _35232_ (_02482_, _02481_, _02480_);
  nor _35233_ (_02484_, _02482_, _02479_);
  nand _35234_ (_02485_, _02484_, _02451_);
  nor _35235_ (_02486_, _02485_, _02450_);
  nand _35236_ (_02487_, _02486_, _02441_);
  nor _35237_ (_02488_, _02487_, _26486_);
  nand _35238_ (_02490_, _02428_, _27699_);
  nand _35239_ (_02491_, _02490_, _27603_);
  nand _35240_ (_02492_, _02491_, _26486_);
  nand _35241_ (_02493_, _02492_, _26487_);
  nor _35242_ (_28211_[8], _02493_, _02488_);
  nand _35243_ (_02494_, _27603_, _27581_);
  nand _35244_ (_02495_, _02494_, _27605_);
  nor _35245_ (_02497_, _02495_, _26485_);
  not _35246_ (_02498_, _26777_);
  nor _35247_ (_02499_, _02498_, _26529_);
  not _35248_ (_02500_, _26752_);
  nor _35249_ (_02501_, _02500_, _26528_);
  nor _35250_ (_02502_, _02501_, _02499_);
  nor _35251_ (_02503_, _02502_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _35252_ (_02504_, _02502_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _35253_ (_02505_, _02504_, _26800_);
  nor _35254_ (_02506_, _02505_, _02503_);
  not _35255_ (_02507_, _02039_);
  nor _35256_ (_02508_, _02507_, _02002_);
  nand _35257_ (_02509_, _02508_, _02008_);
  nand _35258_ (_02510_, _02509_, _25613_);
  not _35259_ (_02511_, _27476_);
  nor _35260_ (_02512_, _27479_, _02511_);
  nor _35261_ (_02513_, _27481_, _24089_);
  not _35262_ (_02514_, _02513_);
  nor _35263_ (_02515_, _02514_, _02512_);
  nor _35264_ (_02516_, _27516_, _24497_);
  nor _35265_ (_02517_, _27527_, _24498_);
  nor _35266_ (_02518_, _02517_, _02516_);
  nor _35267_ (_02519_, _02518_, _24439_);
  nand _35268_ (_02520_, _02518_, _24439_);
  not _35269_ (_02521_, _02520_);
  nor _35270_ (_02522_, _02521_, _02519_);
  nor _35271_ (_02523_, _02522_, _24743_);
  nor _35272_ (_02524_, _26940_, _24768_);
  not _35273_ (_02525_, _02524_);
  nor _35274_ (_02526_, _27447_, _24396_);
  nor _35275_ (_02527_, _27212_, _27211_);
  nor _35276_ (_02528_, _02527_, _27273_);
  not _35277_ (_02529_, _02528_);
  nor _35278_ (_02530_, _02529_, _27506_);
  not _35279_ (_02531_, _02530_);
  nor _35280_ (_02532_, _24700_, _24179_);
  nor _35281_ (_02533_, _24751_, _24381_);
  nor _35282_ (_02534_, _02533_, _02532_);
  nand _35283_ (_02535_, _02534_, _02531_);
  nor _35284_ (_02536_, _02535_, _02526_);
  nand _35285_ (_02537_, _02536_, _02525_);
  nor _35286_ (_02538_, _02537_, _02523_);
  not _35287_ (_02539_, _02538_);
  nor _35288_ (_02540_, _02539_, _02515_);
  nor _35289_ (_02541_, _02540_, _02452_);
  nor _35290_ (_02542_, _26495_, _26426_);
  nor _35291_ (_02543_, _01983_, _24973_);
  nor _35292_ (_02544_, _02543_, _02542_);
  nand _35293_ (_02545_, _01977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nand _35294_ (_02546_, _02545_, _02544_);
  nor _35295_ (_02547_, _02546_, _02541_);
  nand _35296_ (_02548_, _02547_, _02510_);
  nor _35297_ (_02549_, _02548_, _02506_);
  nor _35298_ (_02550_, _02549_, _26486_);
  nor _35299_ (_02551_, _02550_, _02497_);
  nor _35300_ (_28211_[9], _02551_, rst);
  not _35301_ (_02552_, _26778_);
  nor _35302_ (_02553_, _02552_, _26529_);
  not _35303_ (_02554_, _26753_);
  nor _35304_ (_02555_, _02554_, _26528_);
  nor _35305_ (_02556_, _02555_, _02553_);
  nand _35306_ (_02557_, _02556_, _24308_);
  not _35307_ (_02558_, _02556_);
  nand _35308_ (_02559_, _02558_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand _35309_ (_02560_, _02559_, _02557_);
  nor _35310_ (_02561_, _02560_, _26801_);
  not _35311_ (_02562_, _02094_);
  nand _35312_ (_02563_, _02562_, _02062_);
  nor _35313_ (_02564_, _02563_, _02068_);
  nor _35314_ (_02565_, _02564_, _25614_);
  nor _35315_ (_02566_, _27484_, _27481_);
  not _35316_ (_02567_, _02566_);
  nand _35317_ (_02568_, _02567_, _27485_);
  nor _35318_ (_02569_, _02568_, _24089_);
  nor _35319_ (_02570_, _27528_, _24498_);
  nor _35320_ (_02572_, _27517_, _24497_);
  nor _35321_ (_02573_, _02572_, _02570_);
  nor _35322_ (_02574_, _02573_, _24353_);
  nand _35323_ (_02575_, _02573_, _24353_);
  nand _35324_ (_02576_, _02575_, _24742_);
  nor _35325_ (_02577_, _02576_, _02574_);
  not _35326_ (_02578_, _27361_);
  nor _35327_ (_02579_, _27360_, _27358_);
  nor _35328_ (_02580_, _02579_, _02578_);
  not _35329_ (_02581_, _02580_);
  nor _35330_ (_02582_, _02581_, _27506_);
  nor _35331_ (_02583_, _24700_, _24549_);
  nor _35332_ (_02584_, _24751_, _24323_);
  nor _35333_ (_02585_, _27447_, _24338_);
  not _35334_ (_02586_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _35335_ (_02587_, _24768_, _02586_);
  nor _35336_ (_02588_, _02587_, _02585_);
  not _35337_ (_02589_, _02588_);
  nor _35338_ (_02590_, _02589_, _02584_);
  not _35339_ (_02591_, _02590_);
  nor _35340_ (_02592_, _02591_, _02583_);
  not _35341_ (_02593_, _02592_);
  nor _35342_ (_02594_, _02593_, _02582_);
  not _35343_ (_02595_, _02594_);
  nor _35344_ (_02596_, _02595_, _02577_);
  not _35345_ (_02597_, _02596_);
  nor _35346_ (_02598_, _02597_, _02569_);
  not _35347_ (_02599_, _02598_);
  nand _35348_ (_02600_, _02599_, _26797_);
  nor _35349_ (_02601_, _01983_, _27729_);
  not _35350_ (_02602_, _26385_);
  nand _35351_ (_02603_, _27566_, _02602_);
  nand _35352_ (_02604_, _01977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nand _35353_ (_02605_, _02604_, _02603_);
  nor _35354_ (_02606_, _02605_, _02601_);
  nand _35355_ (_02607_, _02606_, _02600_);
  nor _35356_ (_02608_, _02607_, _02565_);
  nand _35357_ (_02609_, _02608_, _26485_);
  nor _35358_ (_02610_, _02609_, _02561_);
  nand _35359_ (_02611_, _27605_, _27580_);
  nand _35360_ (_02612_, _02611_, _27607_);
  nand _35361_ (_02613_, _02612_, _26486_);
  nand _35362_ (_02614_, _02613_, _26487_);
  nor _35363_ (_28211_[10], _02614_, _02610_);
  not _35364_ (_02615_, _27571_);
  nor _35365_ (_02616_, _02615_, _27579_);
  not _35366_ (_02617_, _02134_);
  nand _35367_ (_02618_, _02155_, _02133_);
  nor _35368_ (_02619_, _02618_, _02129_);
  nand _35369_ (_02620_, _02619_, _02617_);
  nand _35370_ (_02621_, _02620_, _25613_);
  not _35371_ (_02622_, _27485_);
  nor _35372_ (_02623_, _02622_, _27469_);
  nor _35373_ (_02624_, _27486_, _24089_);
  not _35374_ (_02625_, _02624_);
  nor _35375_ (_02626_, _02625_, _02623_);
  nor _35376_ (_02627_, _27521_, _24497_);
  nor _35377_ (_02628_, _27531_, _24498_);
  nor _35378_ (_02629_, _02628_, _02627_);
  nor _35379_ (_02630_, _02629_, _24285_);
  nand _35380_ (_02631_, _02629_, _24285_);
  nand _35381_ (_02632_, _02631_, _24742_);
  nor _35382_ (_02633_, _02632_, _02630_);
  not _35383_ (_02635_, _27366_);
  nor _35384_ (_02636_, _02635_, _02578_);
  nor _35385_ (_02637_, _02636_, _27367_);
  not _35386_ (_02638_, _02637_);
  nor _35387_ (_02639_, _02638_, _27506_);
  not _35388_ (_02640_, _02639_);
  not _35389_ (_02641_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _35390_ (_02642_, _24768_, _02641_);
  not _35391_ (_02643_, _24701_);
  nor _35392_ (_02644_, _24751_, _24279_);
  nor _35393_ (_02645_, _27447_, _24285_);
  nor _35394_ (_02646_, _02645_, _02644_);
  nand _35395_ (_02647_, _02646_, _02643_);
  nor _35396_ (_02648_, _02647_, _02642_);
  nand _35397_ (_02649_, _02648_, _02640_);
  nor _35398_ (_02650_, _02649_, _02633_);
  not _35399_ (_02651_, _02650_);
  nor _35400_ (_02652_, _02651_, _02626_);
  nor _35401_ (_02653_, _02652_, _02452_);
  nor _35402_ (_02654_, _26495_, _25912_);
  nor _35403_ (_02655_, _02654_, _02653_);
  nand _35404_ (_02656_, _02655_, _02621_);
  nor _35405_ (_02657_, _02656_, _02616_);
  nand _35406_ (_02658_, _02657_, _26485_);
  nor _35407_ (_02659_, _26754_, _26528_);
  nor _35408_ (_02660_, _26779_, _26529_);
  nor _35409_ (_02661_, _02660_, _02659_);
  nand _35410_ (_02662_, _02661_, _24253_);
  not _35411_ (_02663_, _02661_);
  nand _35412_ (_02664_, _02663_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _35413_ (_02665_, _02664_, _02662_);
  nor _35414_ (_02666_, _02665_, _26801_);
  nor _35415_ (_02667_, _02666_, _02658_);
  nand _35416_ (_02668_, _27607_, _27579_);
  nand _35417_ (_02669_, _02668_, _27609_);
  nand _35418_ (_02670_, _02669_, _26486_);
  nand _35419_ (_02671_, _02670_, _26487_);
  nor _35420_ (_28211_[11], _02671_, _02667_);
  not _35421_ (_02672_, _26755_);
  nor _35422_ (_02673_, _02672_, _26528_);
  not _35423_ (_02674_, _26780_);
  nor _35424_ (_02675_, _02674_, _26529_);
  nor _35425_ (_02676_, _02675_, _02673_);
  nand _35426_ (_02677_, _02676_, _24204_);
  not _35427_ (_02678_, _02676_);
  nand _35428_ (_02679_, _02678_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _35429_ (_02680_, _02679_, _02677_);
  nor _35430_ (_02681_, _02680_, _26801_);
  not _35431_ (_02682_, _02202_);
  nand _35432_ (_02683_, _02224_, _02201_);
  nor _35433_ (_02684_, _02683_, _02195_);
  nand _35434_ (_02685_, _02684_, _02682_);
  nand _35435_ (_02686_, _02685_, _25613_);
  nor _35436_ (_02687_, _27489_, _27486_);
  not _35437_ (_02688_, _02687_);
  nand _35438_ (_02689_, _02688_, _27491_);
  nor _35439_ (_02690_, _02689_, _24089_);
  nor _35440_ (_02691_, _24497_, _24285_);
  nand _35441_ (_02692_, _02691_, _27520_);
  not _35442_ (_02693_, _02692_);
  not _35443_ (_02694_, _27532_);
  nor _35444_ (_02695_, _02694_, _24498_);
  nor _35445_ (_02696_, _02695_, _02693_);
  not _35446_ (_02697_, _02696_);
  nor _35447_ (_02698_, _02697_, _24247_);
  nor _35448_ (_02699_, _02696_, _24241_);
  nor _35449_ (_02700_, _02699_, _24743_);
  not _35450_ (_02701_, _02700_);
  nor _35451_ (_02702_, _02701_, _02698_);
  not _35452_ (_02703_, _27369_);
  not _35453_ (_02704_, _27373_);
  nor _35454_ (_02705_, _02704_, _02703_);
  nor _35455_ (_02706_, _02705_, _27375_);
  not _35456_ (_02707_, _02706_);
  nor _35457_ (_02708_, _02707_, _27506_);
  not _35458_ (_02709_, _02708_);
  not _35459_ (_02710_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _35460_ (_02711_, _24768_, _02710_);
  nor _35461_ (_02712_, _24498_, _24243_);
  nor _35462_ (_02713_, _24497_, _24247_);
  nor _35463_ (_02714_, _02713_, _24751_);
  not _35464_ (_02715_, _02714_);
  nor _35465_ (_02716_, _02715_, _02712_);
  not _35466_ (_02717_, _02716_);
  nor _35467_ (_02718_, _24700_, _24428_);
  nor _35468_ (_02719_, _27447_, _24241_);
  nor _35469_ (_02720_, _02719_, _02718_);
  nand _35470_ (_02721_, _02720_, _02717_);
  nor _35471_ (_02722_, _02721_, _02711_);
  nand _35472_ (_02723_, _02722_, _02709_);
  nor _35473_ (_02724_, _02723_, _02702_);
  not _35474_ (_02725_, _02724_);
  nor _35475_ (_02726_, _02725_, _02690_);
  not _35476_ (_02727_, _02726_);
  nand _35477_ (_02728_, _02727_, _26797_);
  nor _35478_ (_02729_, _26495_, _26012_);
  nor _35479_ (_02730_, _02615_, _27578_);
  nor _35480_ (_02731_, _02730_, _02729_);
  nand _35481_ (_02732_, _02731_, _02728_);
  nor _35482_ (_02733_, _02732_, _26486_);
  nand _35483_ (_02734_, _02733_, _02686_);
  nor _35484_ (_02735_, _02734_, _02681_);
  nor _35485_ (_02736_, _27601_, _27581_);
  nand _35486_ (_02737_, _02736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _35487_ (_02738_, _02737_, _27579_);
  nand _35488_ (_02739_, _02738_, _02110_);
  nand _35489_ (_02740_, _02739_, _27578_);
  nand _35490_ (_02741_, _02740_, _27611_);
  nand _35491_ (_02742_, _02741_, _26486_);
  nand _35492_ (_02743_, _02742_, _26487_);
  nor _35493_ (_28211_[12], _02743_, _02735_);
  nor _35494_ (_02745_, _26756_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _35495_ (_02746_, _26756_);
  nor _35496_ (_02747_, _02746_, _24151_);
  nor _35497_ (_02748_, _02747_, _02745_);
  nor _35498_ (_02749_, _02748_, _26528_);
  not _35499_ (_02750_, _26781_);
  nor _35500_ (_02752_, _02750_, _24151_);
  nor _35501_ (_02753_, _02752_, _26782_);
  nor _35502_ (_02754_, _02753_, _26529_);
  nor _35503_ (_02755_, _02754_, _02749_);
  nor _35504_ (_02756_, _02755_, _26801_);
  not _35505_ (_02757_, _02278_);
  nand _35506_ (_02758_, _02302_, _02270_);
  nor _35507_ (_02760_, _02758_, _02266_);
  nand _35508_ (_02761_, _02760_, _02757_);
  nand _35509_ (_02762_, _02761_, _25613_);
  not _35510_ (_02764_, _27491_);
  nor _35511_ (_02765_, _02764_, _27465_);
  nor _35512_ (_02766_, _27492_, _24089_);
  not _35513_ (_02767_, _02766_);
  nor _35514_ (_02768_, _02767_, _02765_);
  nor _35515_ (_02769_, _02694_, _24247_);
  nor _35516_ (_02770_, _02769_, _02693_);
  nor _35517_ (_02771_, _02770_, _02713_);
  nor _35518_ (_02772_, _02771_, _24199_);
  nand _35519_ (_02773_, _02771_, _24199_);
  nand _35520_ (_02775_, _02773_, _24742_);
  nor _35521_ (_02776_, _02775_, _02772_);
  not _35522_ (_02777_, _27344_);
  not _35523_ (_02778_, _27376_);
  nor _35524_ (_02779_, _02778_, _02777_);
  nor _35525_ (_02781_, _02779_, _27377_);
  not _35526_ (_02782_, _02781_);
  nor _35527_ (_02783_, _02782_, _27506_);
  not _35528_ (_02784_, _02783_);
  nor _35529_ (_02785_, _24497_, _24194_);
  nor _35530_ (_02786_, _24498_, _24179_);
  nor _35531_ (_02787_, _02786_, _02785_);
  nor _35532_ (_02788_, _02787_, _24751_);
  nor _35533_ (_02789_, _24700_, _24381_);
  nor _35534_ (_02790_, _27447_, _24194_);
  not _35535_ (_02791_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _35536_ (_02792_, _24768_, _02791_);
  nor _35537_ (_02793_, _02792_, _02790_);
  not _35538_ (_02794_, _02793_);
  nor _35539_ (_02795_, _02794_, _02789_);
  not _35540_ (_02796_, _02795_);
  nor _35541_ (_02797_, _02796_, _02788_);
  nand _35542_ (_02798_, _02797_, _02784_);
  nor _35543_ (_02799_, _02798_, _02776_);
  not _35544_ (_02800_, _02799_);
  nor _35545_ (_02802_, _02800_, _02768_);
  not _35546_ (_02803_, _02802_);
  nand _35547_ (_02804_, _02803_, _26797_);
  nor _35548_ (_02806_, _26495_, _26118_);
  nor _35549_ (_02807_, _02615_, _27577_);
  nor _35550_ (_02808_, _02807_, _02806_);
  nand _35551_ (_02809_, _02808_, _02804_);
  nor _35552_ (_02810_, _02809_, _26486_);
  nand _35553_ (_02811_, _02810_, _02762_);
  nor _35554_ (_02813_, _02811_, _02756_);
  nor _35555_ (_02814_, _02739_, _27578_);
  nand _35556_ (_02815_, _02814_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _35557_ (_02816_, _27611_, _27577_);
  nand _35558_ (_02817_, _02816_, _02815_);
  nand _35559_ (_02818_, _02817_, _26486_);
  nand _35560_ (_02819_, _02818_, _26487_);
  nor _35561_ (_28211_[13], _02819_, _02813_);
  nor _35562_ (_02820_, _26784_, _24529_);
  not _35563_ (_02821_, _26784_);
  nor _35564_ (_02822_, _02821_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _35565_ (_02823_, _02822_, _02820_);
  nor _35566_ (_02824_, _02823_, _26801_);
  nand _35567_ (_02825_, _02373_, _25613_);
  not _35568_ (_02826_, _27496_);
  nor _35569_ (_02828_, _27495_, _27492_);
  nor _35570_ (_02829_, _02828_, _02826_);
  nand _35571_ (_02830_, _02829_, _24088_);
  not _35572_ (_02831_, _27537_);
  nor _35573_ (_02832_, _02831_, _24558_);
  nor _35574_ (_02833_, _27537_, _24555_);
  nor _35575_ (_02835_, _02833_, _02832_);
  nor _35576_ (_02836_, _02835_, _24743_);
  not _35577_ (_02837_, _27331_);
  not _35578_ (_02838_, _27378_);
  nor _35579_ (_02839_, _02838_, _02837_);
  nor _35580_ (_02840_, _02839_, _27379_);
  not _35581_ (_02841_, _02840_);
  nor _35582_ (_02842_, _02841_, _27506_);
  not _35583_ (_02843_, _02842_);
  nor _35584_ (_02844_, _24557_, _24498_);
  nor _35585_ (_02845_, _27538_, _24751_);
  not _35586_ (_02846_, _02845_);
  nor _35587_ (_02847_, _02846_, _02844_);
  nor _35588_ (_02849_, _24700_, _24323_);
  nor _35589_ (_02850_, _27447_, _24555_);
  nand _35590_ (_02851_, _24767_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  not _35591_ (_02852_, _02851_);
  nor _35592_ (_02853_, _02852_, _02850_);
  not _35593_ (_02854_, _02853_);
  nor _35594_ (_02856_, _02854_, _02849_);
  not _35595_ (_02857_, _02856_);
  nor _35596_ (_02858_, _02857_, _02847_);
  nand _35597_ (_02859_, _02858_, _02843_);
  nor _35598_ (_02860_, _02859_, _02836_);
  nand _35599_ (_02861_, _02860_, _02830_);
  nand _35600_ (_02862_, _02861_, _26797_);
  nor _35601_ (_02863_, _26495_, _25985_);
  nor _35602_ (_02864_, _02615_, _27576_);
  nor _35603_ (_02865_, _02864_, _02863_);
  nand _35604_ (_02866_, _02865_, _02862_);
  nor _35605_ (_02867_, _02866_, _26486_);
  nand _35606_ (_02868_, _02867_, _02825_);
  nor _35607_ (_02870_, _02868_, _02824_);
  nand _35608_ (_02871_, _02815_, _27576_);
  nand _35609_ (_02872_, _02871_, _27616_);
  nand _35610_ (_02873_, _02872_, _26486_);
  nand _35611_ (_02875_, _02873_, _26487_);
  nor _35612_ (_28211_[14], _02875_, _02870_);
  nor _35613_ (_02876_, _01913_, _00147_);
  nand _35614_ (_02878_, _02876_, _24717_);
  nor _35615_ (_02879_, _02876_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor _35616_ (_02880_, _02879_, _26245_);
  nand _35617_ (_02881_, _02880_, _02878_);
  nand _35618_ (_02882_, _01919_, _25029_);
  nor _35619_ (_02883_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor _35620_ (_02884_, _02883_, _25631_);
  nand _35621_ (_02886_, _02884_, _02882_);
  nand _35622_ (_02887_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand _35623_ (_02888_, _02887_, _02886_);
  nor _35624_ (_02889_, _02888_, rst);
  nand _35625_ (_23765_, _02889_, _02881_);
  nand _35626_ (_02891_, _27929_, _27926_);
  nand _35627_ (_02892_, _02891_, _27931_);
  nand _35628_ (_02893_, _02892_, _25834_);
  nor _35629_ (_02894_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _35630_ (_02895_, _02894_, _27965_);
  nand _35631_ (_02896_, _02895_, _02893_);
  nand _35632_ (_02897_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nand _35633_ (_28212_[0], _02897_, _02896_);
  not _35634_ (_02899_, _27936_);
  nand _35635_ (_02900_, _27935_, _27931_);
  nand _35636_ (_02901_, _02900_, _02899_);
  nand _35637_ (_02902_, _02901_, _25834_);
  nor _35638_ (_02904_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _35639_ (_02905_, _02904_, _27965_);
  nand _35640_ (_02906_, _02905_, _02902_);
  nand _35641_ (_02907_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nand _35642_ (_28212_[1], _02907_, _02906_);
  nand _35643_ (_02908_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not _35644_ (_02909_, _27942_);
  nand _35645_ (_02910_, _27941_, _27937_);
  nand _35646_ (_02911_, _02910_, _02909_);
  nand _35647_ (_02912_, _02911_, _25834_);
  nor _35648_ (_02913_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _35649_ (_02914_, _02913_, _27965_);
  nand _35650_ (_02915_, _02914_, _02912_);
  nand _35651_ (_28212_[2], _02915_, _02908_);
  nand _35652_ (_02916_, _02909_, _27720_);
  nand _35653_ (_02917_, _02916_, _27943_);
  nand _35654_ (_02918_, _02917_, _25834_);
  nor _35655_ (_02919_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _35656_ (_02920_, _02919_, _27965_);
  nand _35657_ (_02921_, _02920_, _02918_);
  nand _35658_ (_02922_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand _35659_ (_28212_[3], _02922_, _02921_);
  not _35660_ (_02923_, _27947_);
  nand _35661_ (_02924_, _27946_, _27943_);
  nand _35662_ (_02926_, _02924_, _02923_);
  nand _35663_ (_02927_, _02926_, _25834_);
  nor _35664_ (_02928_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _35665_ (_02929_, _02928_, _27965_);
  nand _35666_ (_02930_, _02929_, _02927_);
  nand _35667_ (_02931_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nand _35668_ (_28212_[4], _02931_, _02930_);
  nand _35669_ (_02932_, _02923_, _27714_);
  nand _35670_ (_02933_, _02932_, _27948_);
  nand _35671_ (_02934_, _02933_, _25834_);
  nor _35672_ (_02935_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _35673_ (_02936_, _02935_, _27965_);
  nand _35674_ (_02937_, _02936_, _02934_);
  nand _35675_ (_02938_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nand _35676_ (_28212_[5], _02938_, _02937_);
  not _35677_ (_02939_, _27949_);
  nand _35678_ (_02940_, _27948_, _27711_);
  nand _35679_ (_02941_, _02940_, _02939_);
  nand _35680_ (_02942_, _02941_, _25834_);
  nor _35681_ (_02943_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _35682_ (_02945_, _02943_, _27965_);
  nand _35683_ (_02946_, _02945_, _02942_);
  nand _35684_ (_02947_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nand _35685_ (_28212_[6], _02947_, _02946_);
  nand _35686_ (_02948_, _02939_, _27707_);
  nand _35687_ (_02949_, _02948_, _27950_);
  nand _35688_ (_02950_, _02949_, _25834_);
  nor _35689_ (_02951_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _35690_ (_02952_, _02951_, _27965_);
  nand _35691_ (_02953_, _02952_, _02950_);
  nand _35692_ (_02954_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nand _35693_ (_28212_[7], _02954_, _02953_);
  not _35694_ (_02955_, _27951_);
  nand _35695_ (_02956_, _27950_, _27703_);
  nand _35696_ (_02957_, _02956_, _02955_);
  nand _35697_ (_02959_, _02957_, _25834_);
  nor _35698_ (_02960_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _35699_ (_02961_, _02960_, _27965_);
  nand _35700_ (_02962_, _02961_, _02959_);
  nand _35701_ (_02963_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand _35702_ (_28212_[8], _02963_, _02962_);
  nand _35703_ (_02964_, _02955_, _27696_);
  nand _35704_ (_02965_, _02964_, _27952_);
  nand _35705_ (_02966_, _02965_, _25834_);
  nor _35706_ (_02967_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _35707_ (_02968_, _02967_, _27965_);
  nand _35708_ (_02969_, _02968_, _02966_);
  nand _35709_ (_02971_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nand _35710_ (_28212_[9], _02971_, _02969_);
  not _35711_ (_02972_, _27953_);
  nand _35712_ (_02973_, _27952_, _27692_);
  nand _35713_ (_02974_, _02973_, _02972_);
  nand _35714_ (_02975_, _02974_, _25834_);
  nor _35715_ (_02976_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _35716_ (_02977_, _02976_, _27965_);
  nand _35717_ (_02979_, _02977_, _02975_);
  nand _35718_ (_02980_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nand _35719_ (_28212_[10], _02980_, _02979_);
  nand _35720_ (_02981_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand _35721_ (_02982_, _02972_, _27687_);
  nand _35722_ (_02984_, _02982_, _27954_);
  nand _35723_ (_02985_, _02984_, _25834_);
  nor _35724_ (_02986_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _35725_ (_02987_, _02986_, _27965_);
  nand _35726_ (_02988_, _02987_, _02985_);
  nand _35727_ (_28212_[11], _02988_, _02981_);
  not _35728_ (_02990_, _27955_);
  nand _35729_ (_02991_, _27954_, _27685_);
  nand _35730_ (_02992_, _02991_, _02990_);
  nand _35731_ (_02993_, _02992_, _25834_);
  nor _35732_ (_02994_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _35733_ (_02995_, _02994_, _27965_);
  nand _35734_ (_02996_, _02995_, _02993_);
  nand _35735_ (_02997_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand _35736_ (_28212_[12], _02997_, _02996_);
  nand _35737_ (_02999_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _35738_ (_03000_, _02990_, _27679_);
  nand _35739_ (_03001_, _03000_, _27956_);
  nand _35740_ (_03003_, _03001_, _25834_);
  nor _35741_ (_03004_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _35742_ (_03005_, _03004_, _27965_);
  nand _35743_ (_03006_, _03005_, _03003_);
  nand _35744_ (_28212_[13], _03006_, _02999_);
  nand _35745_ (_03008_, _27956_, _27676_);
  nand _35746_ (_03009_, _03008_, _27959_);
  nand _35747_ (_03011_, _03009_, _25834_);
  nor _35748_ (_03012_, _25834_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _35749_ (_03013_, _03012_, _27965_);
  nand _35750_ (_03014_, _03013_, _03011_);
  nand _35751_ (_03015_, _27622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _35752_ (_28212_[14], _03015_, _03014_);
  nor _35753_ (_03016_, _01913_, _01666_);
  nand _35754_ (_03017_, _03016_, _24717_);
  nor _35755_ (_03018_, _03016_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _35756_ (_03019_, _03018_, _26245_);
  nand _35757_ (_03020_, _03019_, _03017_);
  nand _35758_ (_03021_, _01919_, _25140_);
  nor _35759_ (_03022_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _35760_ (_03023_, _03022_, _25631_);
  nand _35761_ (_03024_, _03023_, _03021_);
  nand _35762_ (_03025_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nand _35763_ (_03026_, _03025_, _03024_);
  nor _35764_ (_03028_, _03026_, rst);
  nand _35765_ (_23766_, _03028_, _03020_);
  nor _35766_ (_03029_, _27976_, _26703_);
  nor _35767_ (_03031_, _03029_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor _35768_ (_28216_[0], _03031_, rst);
  nor _35769_ (_03032_, _27976_, _26677_);
  nor _35770_ (_03033_, _03032_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor _35771_ (_28216_[1], _03033_, rst);
  nor _35772_ (_03034_, _27976_, _26649_);
  nor _35773_ (_03035_, _03034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor _35774_ (_28216_[2], _03035_, rst);
  nor _35775_ (_03036_, _27976_, _26618_);
  nor _35776_ (_03037_, _03036_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _35777_ (_28216_[3], _03037_, rst);
  nor _35778_ (_03038_, _27976_, _26589_);
  nor _35779_ (_03039_, _03038_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _35780_ (_28216_[4], _03039_, rst);
  nor _35781_ (_03040_, _27976_, _26563_);
  nor _35782_ (_03041_, _03040_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor _35783_ (_28216_[5], _03041_, rst);
  nor _35784_ (_03043_, _27976_, _26535_);
  nor _35785_ (_03044_, _03043_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor _35786_ (_28216_[6], _03044_, rst);
  nor _35787_ (_03045_, _01913_, _00135_);
  nand _35788_ (_03047_, _03045_, _24717_);
  nor _35789_ (_03048_, _03045_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor _35790_ (_03049_, _03048_, _26245_);
  nand _35791_ (_03050_, _03049_, _03047_);
  nand _35792_ (_03051_, _01919_, _26096_);
  nor _35793_ (_03052_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor _35794_ (_03053_, _03052_, _25631_);
  nand _35795_ (_03054_, _03053_, _03051_);
  nand _35796_ (_03055_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand _35797_ (_03056_, _03055_, _03054_);
  nor _35798_ (_03057_, _03056_, rst);
  nand _35799_ (_23767_, _03057_, _03050_);
  not _35800_ (_03058_, _27926_);
  nand _35801_ (_03059_, _03058_, _24863_);
  nor _35802_ (_03060_, _03059_, _24938_);
  nand _35803_ (_03061_, _03059_, _24938_);
  nand _35804_ (_03062_, _03061_, _27964_);
  nor _35805_ (_28217_[0], _03062_, _03060_);
  nor _35806_ (_03063_, _27988_, _27986_);
  nor _35807_ (_03064_, _03063_, _27990_);
  nor _35808_ (_03065_, _03064_, _24864_);
  nand _35809_ (_03066_, _24864_, _24960_);
  nand _35810_ (_03067_, _03066_, _27964_);
  nor _35811_ (_28217_[1], _03067_, _03065_);
  nor _35812_ (_03068_, _01913_, _00263_);
  nand _35813_ (_03069_, _03068_, _24717_);
  nor _35814_ (_03070_, _03068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor _35815_ (_03072_, _03070_, _26245_);
  nand _35816_ (_03073_, _03072_, _03069_);
  nand _35817_ (_03074_, _01919_, _25195_);
  nor _35818_ (_03075_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor _35819_ (_03076_, _03075_, _25631_);
  nand _35820_ (_03077_, _03076_, _03074_);
  nand _35821_ (_03079_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nand _35822_ (_03080_, _03079_, _03077_);
  nor _35823_ (_03081_, _03080_, rst);
  nand _35824_ (_23768_, _03081_, _03073_);
  nor _35825_ (_03082_, _25159_, _24059_);
  nand _35826_ (_03083_, _03082_, _25099_);
  not _35827_ (_03085_, _03082_);
  nand _35828_ (_03086_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand _35829_ (_23769_, _03086_, _03083_);
  nand _35830_ (_03088_, _03082_, _25203_);
  nand _35831_ (_03089_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nand _35832_ (_23770_, _03089_, _03088_);
  nand _35833_ (_03090_, _03082_, _25039_);
  nand _35834_ (_03091_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nand _35835_ (_23771_, _03091_, _03090_);
  nand _35836_ (_03092_, _03082_, _25150_);
  nand _35837_ (_03093_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nand _35838_ (_23772_, _03093_, _03092_);
  nor _35839_ (_03094_, _25627_, _01549_);
  nand _35840_ (_03095_, _03094_, _24717_);
  nor _35841_ (_03097_, _03094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _35842_ (_03098_, _03097_, _26245_);
  nand _35843_ (_03099_, _03098_, _03095_);
  nand _35844_ (_03100_, _03094_, _24820_);
  nand _35845_ (_03101_, _03100_, _25630_);
  nor _35846_ (_03103_, _03101_, _03097_);
  nand _35847_ (_03104_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand _35848_ (_03105_, _03104_, _26487_);
  nor _35849_ (_03106_, _03105_, _03103_);
  nand _35850_ (_23773_, _03106_, _03099_);
  nor _35851_ (_03107_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _35852_ (_03108_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _35853_ (_03109_, _03108_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _35854_ (_03110_, _03109_, _26487_);
  nor _35855_ (_28221_[0], _03110_, _03107_);
  nor _35856_ (_03111_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _35857_ (_03112_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _35858_ (_03113_, _03112_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _35859_ (_03114_, _03113_, _26487_);
  nor _35860_ (_28221_[1], _03114_, _03111_);
  nor _35861_ (_03115_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _35862_ (_03116_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _35863_ (_03117_, _03116_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _35864_ (_03119_, _03117_, _26487_);
  nor _35865_ (_28221_[2], _03119_, _03115_);
  nor _35866_ (_03120_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _35867_ (_03122_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand _35868_ (_03123_, _03122_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _35869_ (_03124_, _03123_, _26487_);
  nor _35870_ (_28221_[3], _03124_, _03120_);
  nor _35871_ (_03125_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _35872_ (_03126_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand _35873_ (_03127_, _03126_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _35874_ (_03128_, _03127_, _26487_);
  nor _35875_ (_28221_[4], _03128_, _03125_);
  nor _35876_ (_03130_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _35877_ (_03131_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _35878_ (_03132_, _03131_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _35879_ (_03134_, _03132_, _26487_);
  nor _35880_ (_28221_[5], _03134_, _03130_);
  nor _35881_ (_03135_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _35882_ (_03136_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _35883_ (_03137_, _03136_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand _35884_ (_03138_, _03137_, _26487_);
  nor _35885_ (_28221_[6], _03138_, _03135_);
  nor _35886_ (_03139_, _25159_, _25057_);
  nand _35887_ (_03140_, _03139_, _25099_);
  not _35888_ (_03141_, _03139_);
  nand _35889_ (_03142_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nand _35890_ (_23774_, _03142_, _03140_);
  nor _35891_ (_28224_[0], _28027_, rst);
  nor _35892_ (_28224_[1], _28040_, rst);
  nor _35893_ (_28224_[2], _28035_, rst);
  nand _35894_ (_03145_, _03139_, _28096_);
  nand _35895_ (_03146_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nand _35896_ (_23775_, _03146_, _03145_);
  nor _35897_ (_03147_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand _35898_ (_03148_, _27586_, _25443_);
  nand _35899_ (_03149_, _03148_, _26487_);
  nor _35900_ (_28226_[0], _03149_, _03147_);
  nor _35901_ (_03150_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand _35902_ (_03151_, _27586_, _25248_);
  nand _35903_ (_03152_, _03151_, _26487_);
  nor _35904_ (_28226_[1], _03152_, _03150_);
  nor _35905_ (_03153_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand _35906_ (_03154_, _27586_, _25269_);
  nand _35907_ (_03155_, _03154_, _26487_);
  nor _35908_ (_28226_[2], _03155_, _03153_);
  nor _35909_ (_03156_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand _35910_ (_03157_, _27586_, _25218_);
  nand _35911_ (_03158_, _03157_, _26487_);
  nor _35912_ (_28226_[3], _03158_, _03156_);
  nor _35913_ (_03160_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand _35914_ (_03162_, _27586_, _25309_);
  nand _35915_ (_03163_, _03162_, _26487_);
  nor _35916_ (_28226_[4], _03163_, _03160_);
  nor _35917_ (_03164_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand _35918_ (_03165_, _27586_, _25373_);
  nand _35919_ (_03166_, _03165_, _26487_);
  nor _35920_ (_28226_[5], _03166_, _03164_);
  nor _35921_ (_03168_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand _35922_ (_03169_, _27586_, _24956_);
  nand _35923_ (_03170_, _03169_, _26487_);
  nor _35924_ (_28226_[6], _03170_, _03168_);
  nor _35925_ (_03171_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand _35926_ (_03172_, _27586_, _25341_);
  nand _35927_ (_03173_, _03172_, _26487_);
  nor _35928_ (_28226_[7], _03173_, _03171_);
  nor _35929_ (_03174_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _35930_ (_03175_, _27586_, _25434_);
  nand _35931_ (_03176_, _03175_, _26487_);
  nor _35932_ (_28226_[8], _03176_, _03174_);
  nor _35933_ (_03177_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _35934_ (_03178_, _27586_, _25250_);
  nand _35935_ (_03179_, _03178_, _26487_);
  nor _35936_ (_28226_[9], _03179_, _03177_);
  nor _35937_ (_03180_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand _35938_ (_03181_, _27586_, _25282_);
  nand _35939_ (_03182_, _03181_, _26487_);
  nor _35940_ (_28226_[10], _03182_, _03180_);
  nor _35941_ (_03183_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _35942_ (_03184_, _27586_, _25210_);
  nand _35943_ (_03185_, _03184_, _26487_);
  nor _35944_ (_28226_[11], _03185_, _03183_);
  nor _35945_ (_03186_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand _35946_ (_03187_, _27586_, _25311_);
  nand _35947_ (_03188_, _03187_, _26487_);
  nor _35948_ (_28226_[12], _03188_, _03186_);
  nor _35949_ (_03189_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _35950_ (_03190_, _27586_, _25364_);
  nand _35951_ (_03191_, _03190_, _26487_);
  nor _35952_ (_28226_[13], _03191_, _03189_);
  nor _35953_ (_03192_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _35954_ (_03193_, _27586_, _24935_);
  nand _35955_ (_03194_, _03193_, _26487_);
  nor _35956_ (_28226_[14], _03194_, _03192_);
  nor _35957_ (_03195_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _35958_ (_03197_, _27586_, _25330_);
  nand _35959_ (_03198_, _03197_, _26487_);
  nor _35960_ (_28226_[15], _03198_, _03195_);
  nor _35961_ (_03199_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _35962_ (_03200_, _27586_, _25432_);
  nand _35963_ (_03201_, _03200_, _26487_);
  nor _35964_ (_28226_[16], _03201_, _03199_);
  nor _35965_ (_03203_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _35966_ (_03204_, _27586_, _25253_);
  nand _35967_ (_03205_, _03204_, _26487_);
  nor _35968_ (_28226_[17], _03205_, _03203_);
  nor _35969_ (_03206_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _35970_ (_03207_, _27586_, _25271_);
  nand _35971_ (_03208_, _03207_, _26487_);
  nor _35972_ (_28226_[18], _03208_, _03206_);
  nor _35973_ (_03209_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _35974_ (_03210_, _27586_, _25903_);
  nand _35975_ (_03211_, _03210_, _26487_);
  nor _35976_ (_28226_[19], _03211_, _03209_);
  nor _35977_ (_03213_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand _35978_ (_03214_, _27586_, _25314_);
  nand _35979_ (_03215_, _03214_, _26487_);
  nor _35980_ (_28226_[20], _03215_, _03213_);
  nor _35981_ (_03216_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _35982_ (_03217_, _27586_, _25362_);
  nand _35983_ (_03218_, _03217_, _26487_);
  nor _35984_ (_28226_[21], _03218_, _03216_);
  nor _35985_ (_03220_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _35986_ (_03221_, _27586_, _24959_);
  nand _35987_ (_03222_, _03221_, _26487_);
  nor _35988_ (_28226_[22], _03222_, _03220_);
  nor _35989_ (_03223_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _35990_ (_03224_, _27586_, _25332_);
  nand _35991_ (_03225_, _03224_, _26487_);
  nor _35992_ (_28226_[23], _03225_, _03223_);
  nor _35993_ (_03226_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand _35994_ (_03227_, _27586_, _26314_);
  nand _35995_ (_03228_, _03227_, _26487_);
  nor _35996_ (_28226_[24], _03228_, _03226_);
  nor _35997_ (_03229_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _35998_ (_03230_, _27586_, _25242_);
  nand _35999_ (_03231_, _03230_, _26487_);
  nor _36000_ (_28226_[25], _03231_, _03229_);
  nor _36001_ (_03232_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _36002_ (_03233_, _27586_, _26370_);
  nand _36003_ (_03234_, _03233_, _26487_);
  nor _36004_ (_28226_[26], _03234_, _03232_);
  nor _36005_ (_03235_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _36006_ (_03236_, _27586_, _25897_);
  nand _36007_ (_03237_, _03236_, _26487_);
  nor _36008_ (_28226_[27], _03237_, _03235_);
  nor _36009_ (_03238_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand _36010_ (_03239_, _27586_, _25304_);
  nand _36011_ (_03240_, _03239_, _26487_);
  nor _36012_ (_28226_[28], _03240_, _03238_);
  nor _36013_ (_03242_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _36014_ (_03243_, _27586_, _26102_);
  nand _36015_ (_03244_, _03243_, _26487_);
  nor _36016_ (_28226_[29], _03244_, _03242_);
  nor _36017_ (_03246_, _27586_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand _36018_ (_03248_, _27586_, _25971_);
  nand _36019_ (_03249_, _03248_, _26487_);
  nor _36020_ (_28226_[30], _03249_, _03246_);
  nand _36021_ (_03250_, _03139_, _25039_);
  nand _36022_ (_03251_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nand _36023_ (_23776_, _03251_, _03250_);
  not _36024_ (_03252_, _26239_);
  nor _36025_ (_03253_, _03252_, _00617_);
  not _36026_ (_03254_, _03253_);
  nor _36027_ (_03255_, _00263_, _03254_);
  nand _36028_ (_03256_, _03255_, _24717_);
  nor _36029_ (_03257_, _03255_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor _36030_ (_03258_, _03257_, _26245_);
  nand _36031_ (_03259_, _03258_, _03256_);
  not _36032_ (_03260_, _03094_);
  nor _36033_ (_03261_, _03260_, _25194_);
  not _36034_ (_03262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nand _36035_ (_03263_, _03260_, _03262_);
  nand _36036_ (_03264_, _03263_, _25630_);
  nor _36037_ (_03265_, _03264_, _03261_);
  nand _36038_ (_03266_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nand _36039_ (_03267_, _03266_, _26487_);
  nor _36040_ (_03268_, _03267_, _03265_);
  nand _36041_ (_23777_, _03268_, _03259_);
  nand _36042_ (_03269_, _03139_, _25150_);
  nand _36043_ (_03270_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nand _36044_ (_23778_, _03270_, _03269_);
  nor _36045_ (_03271_, _01666_, _03254_);
  nand _36046_ (_03272_, _03271_, _24717_);
  nor _36047_ (_03273_, _03271_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _36048_ (_03274_, _03273_, _26245_);
  nand _36049_ (_03275_, _03274_, _03272_);
  nand _36050_ (_03276_, _03094_, _25140_);
  nor _36051_ (_03277_, _03094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _36052_ (_03278_, _03277_, _25631_);
  nand _36053_ (_03279_, _03278_, _03276_);
  nand _36054_ (_03280_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nand _36055_ (_03281_, _03280_, _03279_);
  nor _36056_ (_03282_, _03281_, rst);
  nand _36057_ (_23779_, _03282_, _03275_);
  nor _36058_ (_03283_, _00135_, _03254_);
  nand _36059_ (_03284_, _03283_, _24717_);
  nor _36060_ (_03285_, _03283_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor _36061_ (_03286_, _03285_, _26245_);
  nand _36062_ (_03287_, _03286_, _03284_);
  nand _36063_ (_03288_, _03094_, _26096_);
  nor _36064_ (_03289_, _03094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor _36065_ (_03290_, _03289_, _25631_);
  nand _36066_ (_03291_, _03290_, _03288_);
  nand _36067_ (_03292_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand _36068_ (_03293_, _03292_, _03291_);
  nor _36069_ (_03294_, _03293_, rst);
  nand _36070_ (_23780_, _03294_, _03287_);
  nor _36071_ (_03295_, _01974_, _28052_);
  not _36072_ (_03296_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nand _36073_ (_03297_, _28052_, _03296_);
  nand _36074_ (_03298_, _03297_, _26487_);
  nor _36075_ (_28230_[0], _03298_, _03295_);
  nor _36076_ (_03299_, _02509_, _28052_);
  not _36077_ (_03300_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nand _36078_ (_03301_, _28052_, _03300_);
  nand _36079_ (_03302_, _03301_, _26487_);
  nor _36080_ (_28230_[1], _03302_, _03299_);
  nor _36081_ (_03303_, _02096_, _28052_);
  not _36082_ (_03304_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nand _36083_ (_03305_, _28052_, _03304_);
  nand _36084_ (_03306_, _03305_, _26487_);
  nor _36085_ (_28230_[2], _03306_, _03303_);
  nor _36086_ (_03307_, _02620_, _28052_);
  not _36087_ (_03308_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nand _36088_ (_03309_, _28052_, _03308_);
  nand _36089_ (_03310_, _03309_, _26487_);
  nor _36090_ (_28230_[3], _03310_, _03307_);
  nand _36091_ (_03311_, _00377_, _03253_);
  nand _36092_ (_03312_, _03311_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand _36093_ (_03313_, _00384_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand _36094_ (_03314_, _03313_, _00381_);
  nand _36095_ (_03315_, _03314_, _03253_);
  nand _36096_ (_03316_, _03315_, _03312_);
  nand _36097_ (_03317_, _03316_, _26244_);
  nand _36098_ (_03318_, _03260_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand _36099_ (_03319_, _03094_, _25028_);
  nand _36100_ (_03320_, _03319_, _03318_);
  nand _36101_ (_03321_, _03320_, _25630_);
  nand _36102_ (_03322_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand _36103_ (_03323_, _03322_, _03321_);
  nor _36104_ (_03324_, _03323_, rst);
  nand _36105_ (_23781_, _03324_, _03317_);
  nor _36106_ (_03325_, _00276_, _03254_);
  nand _36107_ (_03326_, _03325_, _24717_);
  nor _36108_ (_03327_, _03325_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor _36109_ (_03328_, _03327_, _26245_);
  nand _36110_ (_03329_, _03328_, _03326_);
  nand _36111_ (_03330_, _03094_, _25703_);
  nor _36112_ (_03331_, _03094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor _36113_ (_03332_, _03331_, _25631_);
  nand _36114_ (_03333_, _03332_, _03330_);
  nand _36115_ (_03334_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nand _36116_ (_03335_, _03334_, _03333_);
  nor _36117_ (_03336_, _03335_, rst);
  nand _36118_ (_23782_, _03336_, _03329_);
  nand _36119_ (_03337_, _25160_, _25099_);
  nand _36120_ (_03338_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand _36121_ (_23783_, _03338_, _03337_);
  nand _36122_ (_03340_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nand _36123_ (_03341_, _01520_, _25203_);
  nand _36124_ (_23784_, _03341_, _03340_);
  nand _36125_ (_03343_, _28096_, _25160_);
  nand _36126_ (_03344_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand _36127_ (_23785_, _03344_, _03343_);
  nand _36128_ (_03345_, _25160_, _25039_);
  nand _36129_ (_03346_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand _36130_ (_23786_, _03346_, _03345_);
  nand _36131_ (_03347_, _01278_, _01665_);
  nor _36132_ (_03348_, _03347_, _24717_);
  not _36133_ (_03349_, _01287_);
  nand _36134_ (_03350_, _03347_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _36135_ (_03351_, _03350_, _03349_);
  nor _36136_ (_03352_, _03351_, _03348_);
  nand _36137_ (_03353_, _01287_, _25140_);
  nand _36138_ (_03354_, _03353_, _26487_);
  nor _36139_ (_23787_, _03354_, _03352_);
  not _36140_ (_03355_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  not _36141_ (_03356_, _00135_);
  nand _36142_ (_03357_, _01278_, _03356_);
  nand _36143_ (_03358_, _03357_, _03355_);
  nand _36144_ (_03359_, _03358_, _01293_);
  nor _36145_ (_03360_, _03357_, _24716_);
  nor _36146_ (_03361_, _03360_, _03359_);
  nor _36147_ (_03362_, _01293_, _26096_);
  nor _36148_ (_03363_, _03362_, _03361_);
  nor _36149_ (_23788_, _03363_, rst);
  nor _36150_ (_03364_, _00265_, _25627_);
  nand _36151_ (_03365_, _03364_, _26244_);
  nor _36152_ (_03366_, _03365_, _24716_);
  nor _36153_ (_03367_, _00786_, _00651_);
  nor _36154_ (_03368_, _03367_, _00540_);
  nand _36155_ (_03369_, _03368_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nand _36156_ (_03370_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _00535_);
  nand _36157_ (_03371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _36158_ (_03372_, _03371_, _03370_);
  nand _36159_ (_03373_, _03372_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _36160_ (_03374_, _03373_);
  nor _36161_ (_03375_, _00742_, _00701_);
  nor _36162_ (_03376_, _03375_, _00540_);
  not _36163_ (_03377_, _03376_);
  nor _36164_ (_03378_, _03377_, _03374_);
  not _36165_ (_03380_, _03378_);
  nor _36166_ (_03381_, _03380_, _03369_);
  nor _36167_ (_03382_, _03381_, _00562_);
  nand _36168_ (_03383_, _03382_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _36169_ (_03384_, _03365_, _03383_);
  nand _36170_ (_03385_, _03384_, _00622_);
  nor _36171_ (_03387_, _03385_, _03366_);
  nor _36172_ (_03388_, _00622_, _25195_);
  nor _36173_ (_03389_, _03388_, _03387_);
  nor _36174_ (_23789_, _03389_, rst);
  nand _36175_ (_03390_, _00429_, _01665_);
  nor _36176_ (_03391_, _03390_, _24716_);
  not _36177_ (_03392_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand _36178_ (_03393_, _03390_, _03392_);
  nand _36179_ (_03394_, _03393_, _00438_);
  nor _36180_ (_03395_, _03394_, _03391_);
  nor _36181_ (_03396_, _00438_, _25140_);
  nor _36182_ (_03397_, _03396_, _03395_);
  nor _36183_ (_23790_, _03397_, rst);
  nand _36184_ (_03398_, _00494_, _03356_);
  nor _36185_ (_03399_, _03398_, _24716_);
  nand _36186_ (_03400_, _03398_, _00578_);
  nand _36187_ (_03402_, _03400_, _00503_);
  nor _36188_ (_03404_, _03402_, _03399_);
  nor _36189_ (_03405_, _00503_, _26096_);
  nor _36190_ (_03407_, _03405_, _03404_);
  nor _36191_ (_23791_, _03407_, rst);
  nor _36192_ (_03408_, _01277_, _00219_);
  nand _36193_ (_03409_, _03408_, _00146_);
  nand _36194_ (_03410_, _03409_, _01582_);
  nand _36195_ (_03411_, _03410_, _00622_);
  nor _36196_ (_03412_, _03409_, _24716_);
  nor _36197_ (_03413_, _03412_, _03411_);
  nor _36198_ (_03414_, _00622_, _25029_);
  nor _36199_ (_03415_, _03414_, _03413_);
  nor _36200_ (_23792_, _03415_, rst);
  nand _36201_ (_03416_, _00991_, _24830_);
  nand _36202_ (_03417_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  nand _36203_ (_23793_, _03417_, _03416_);
  nand _36204_ (_03418_, _00683_, _00698_);
  not _36205_ (_03420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _36206_ (_03421_, _00598_, _03420_);
  nor _36207_ (_03422_, _03421_, _03418_);
  nor _36208_ (_03423_, _03422_, _00607_);
  nand _36209_ (_03424_, _03423_, _00668_);
  nand _36210_ (_03426_, _00794_, _00661_);
  nand _36211_ (_03427_, _00722_, _00656_);
  nor _36212_ (_03428_, _00584_, _03420_);
  nor _36213_ (_03429_, _03428_, _03427_);
  nor _36214_ (_03431_, _03429_, _03426_);
  nand _36215_ (_03432_, _03431_, _00590_);
  nand _36216_ (_03433_, _03432_, _03424_);
  nor _36217_ (_03434_, _03433_, _00537_);
  nand _36218_ (_03436_, _00537_, _03420_);
  nand _36219_ (_03437_, _03436_, _26487_);
  nor _36220_ (_23794_, _03437_, _03434_);
  nand _36221_ (_03439_, _25160_, _25150_);
  nand _36222_ (_03440_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand _36223_ (_23795_, _03440_, _03439_);
  nor _36224_ (_03442_, _00393_, _24889_);
  nand _36225_ (_03443_, _03442_, _24927_);
  not _36226_ (_03444_, _03442_);
  nand _36227_ (_03445_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  nand _36228_ (_23796_, _03445_, _03443_);
  nor _36229_ (_03446_, _25159_, _24978_);
  nand _36230_ (_03447_, _03446_, _24830_);
  not _36231_ (_03449_, _03446_);
  nand _36232_ (_03450_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nand _36233_ (_23797_, _03450_, _03447_);
  nand _36234_ (_03451_, _00494_, _01665_);
  nor _36235_ (_03453_, _03451_, _24716_);
  not _36236_ (_03454_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  nand _36237_ (_03455_, _03451_, _03454_);
  nand _36238_ (_03456_, _03455_, _00503_);
  nor _36239_ (_03457_, _03456_, _03453_);
  nor _36240_ (_03458_, _00503_, _25140_);
  nor _36241_ (_03459_, _03458_, _03457_);
  nor _36242_ (_23798_, _03459_, rst);
  nand _36243_ (_03460_, _03446_, _28096_);
  nand _36244_ (_03461_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand _36245_ (_23799_, _03461_, _03460_);
  nand _36246_ (_03462_, _03446_, _25039_);
  nand _36247_ (_03463_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand _36248_ (_23800_, _03463_, _03462_);
  nand _36249_ (_03464_, _03446_, _25150_);
  nand _36250_ (_03465_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nand _36251_ (_23801_, _03465_, _03464_);
  nand _36252_ (_03466_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nand _36253_ (_03467_, _01520_, _28096_);
  nand _36254_ (_23802_, _03467_, _03466_);
  nand _36255_ (_03468_, _00955_, _25039_);
  nand _36256_ (_03469_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nand _36257_ (_23803_, _03469_, _03468_);
  nand _36258_ (_03470_, _03082_, _24830_);
  nand _36259_ (_03471_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand _36260_ (_23804_, _03471_, _03470_);
  not _36261_ (_03472_, _00811_);
  nor _36262_ (_03473_, _00596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _36263_ (_03474_, _03473_, _00595_);
  nor _36264_ (_03475_, _03474_, _00599_);
  nor _36265_ (_03476_, _03475_, _00608_);
  nor _36266_ (_03477_, _03476_, _00604_);
  nor _36267_ (_03478_, _03477_, _03472_);
  nor _36268_ (_03479_, _00591_, _00554_);
  not _36269_ (_03480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nand _36270_ (_03481_, _00744_, _03480_);
  nand _36271_ (_03482_, _03481_, _00645_);
  nand _36272_ (_03483_, _03482_, _00722_);
  nand _36273_ (_03484_, _03483_, _00656_);
  nand _36274_ (_03485_, _03484_, _00794_);
  nand _36275_ (_03486_, _03485_, _03479_);
  nand _36276_ (_03487_, _03486_, _00536_);
  nor _36277_ (_03488_, _03487_, _03478_);
  nand _36278_ (_03489_, _00537_, _03480_);
  nand _36279_ (_03490_, _03489_, _26487_);
  nor _36280_ (_23805_, _03490_, _03488_);
  not _36281_ (_03491_, _00840_);
  nor _36282_ (_03492_, _03491_, _00669_);
  nand _36283_ (_03493_, _00840_, _00590_);
  nand _36284_ (_03494_, _03493_, _00541_);
  nand _36285_ (_03495_, _03494_, _26487_);
  nor _36286_ (_23806_, _03495_, _03492_);
  not _36287_ (_03496_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _36288_ (_03497_, _03408_, _00275_);
  nand _36289_ (_03498_, _03497_, _03496_);
  nand _36290_ (_03499_, _03498_, _00622_);
  nor _36291_ (_03500_, _03497_, _24716_);
  nor _36292_ (_03501_, _03500_, _03499_);
  nor _36293_ (_03502_, _00622_, _25703_);
  nor _36294_ (_03503_, _03502_, _03501_);
  nor _36295_ (_23807_, _03503_, rst);
  nor _36296_ (_03504_, _00385_, _00571_);
  nor _36297_ (_03505_, _03504_, _00382_);
  nor _36298_ (_03506_, _03505_, _00495_);
  nand _36299_ (_03507_, _00494_, _00377_);
  nand _36300_ (_03508_, _03507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _36301_ (_03509_, _03508_, _00503_);
  nor _36302_ (_03510_, _03509_, _03506_);
  nand _36303_ (_03511_, _00506_, _25029_);
  nand _36304_ (_03512_, _03511_, _26487_);
  nor _36305_ (_23808_, _03512_, _03510_);
  nand _36306_ (_03513_, _00429_, _03356_);
  nor _36307_ (_03514_, _03513_, _24716_);
  nand _36308_ (_03515_, _03513_, _00577_);
  nand _36309_ (_03516_, _03515_, _00438_);
  nor _36310_ (_03517_, _03516_, _03514_);
  nor _36311_ (_03518_, _00438_, _26096_);
  nor _36312_ (_03519_, _03518_, _03517_);
  nor _36313_ (_23809_, _03519_, rst);
  nor _36314_ (_03520_, _25159_, _24795_);
  nand _36315_ (_03521_, _03520_, _25099_);
  not _36316_ (_03522_, _03520_);
  nand _36317_ (_03523_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nand _36318_ (_23810_, _03523_, _03521_);
  nand _36319_ (_03524_, _03520_, _25203_);
  nand _36320_ (_03525_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nand _36321_ (_23811_, _03525_, _03524_);
  nand _36322_ (_03526_, _03520_, _24927_);
  nand _36323_ (_03527_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nand _36324_ (_23812_, _03527_, _03526_);
  nand _36325_ (_03528_, _03520_, _25039_);
  nand _36326_ (_03529_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nand _36327_ (_23813_, _03529_, _03528_);
  nand _36328_ (_03530_, _03520_, _24789_);
  nand _36329_ (_03531_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand _36330_ (_23814_, _03531_, _03530_);
  nand _36331_ (_03532_, _01178_, _25099_);
  nand _36332_ (_03533_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand _36333_ (_23815_, _03533_, _03532_);
  nand _36334_ (_03534_, _01178_, _25203_);
  nand _36335_ (_03535_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand _36336_ (_23816_, _03535_, _03534_);
  nand _36337_ (_03536_, _01178_, _25150_);
  nand _36338_ (_03537_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand _36339_ (_23817_, _03537_, _03536_);
  nand _36340_ (_03538_, _01178_, _24789_);
  nand _36341_ (_03539_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nand _36342_ (_23818_, _03539_, _03538_);
  nor _36343_ (_03540_, _00114_, _24993_);
  nand _36344_ (_03541_, _03540_, _25099_);
  not _36345_ (_03542_, _03540_);
  nand _36346_ (_03543_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nand _36347_ (_23819_, _03543_, _03541_);
  nor _36348_ (_03545_, _24982_, _24071_);
  not _36349_ (_03546_, _03545_);
  nor _36350_ (_03547_, _03546_, _00926_);
  not _36351_ (_03548_, _03547_);
  nand _36352_ (_03549_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  nand _36353_ (_03550_, _03547_, _25099_);
  nand _36354_ (_23820_, _03550_, _03549_);
  nand _36355_ (_03551_, _03540_, _25203_);
  nand _36356_ (_03552_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  nand _36357_ (_23821_, _03552_, _03551_);
  nand _36358_ (_03553_, _03540_, _24927_);
  nand _36359_ (_03554_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  nand _36360_ (_23822_, _03554_, _03553_);
  nand _36361_ (_03555_, _00479_, _28096_);
  nand _36362_ (_03556_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nand _36363_ (_23823_, _03556_, _03555_);
  nand _36364_ (_03557_, _03540_, _24789_);
  nand _36365_ (_03558_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  nand _36366_ (_23824_, _03558_, _03557_);
  nand _36367_ (_03559_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  nand _36368_ (_03560_, _03547_, _24830_);
  nand _36369_ (_23825_, _03560_, _03559_);
  nor _36370_ (_03561_, _00629_, _24993_);
  nand _36371_ (_03562_, _03561_, _24830_);
  not _36372_ (_03563_, _03561_);
  nand _36373_ (_03564_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nand _36374_ (_23826_, _03564_, _03562_);
  nand _36375_ (_03565_, _03561_, _25203_);
  nand _36376_ (_03566_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nand _36377_ (_23827_, _03566_, _03565_);
  nand _36378_ (_03567_, _03561_, _24927_);
  nand _36379_ (_03568_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  nand _36380_ (_23828_, _03568_, _03567_);
  nand _36381_ (_03569_, _03561_, _24789_);
  nand _36382_ (_03570_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  nand _36383_ (_23829_, _03570_, _03569_);
  nor _36384_ (_03571_, _24882_, _24993_);
  nand _36385_ (_03572_, _03571_, _24830_);
  not _36386_ (_03573_, _03571_);
  nand _36387_ (_03575_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  nand _36388_ (_23830_, _03575_, _03572_);
  nand _36389_ (_03576_, _03571_, _28096_);
  nand _36390_ (_03577_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  nand _36391_ (_23831_, _03577_, _03576_);
  nand _36392_ (_03578_, _03571_, _25039_);
  nand _36393_ (_03579_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nand _36394_ (_23832_, _03579_, _03578_);
  nand _36395_ (_03581_, _03571_, _25150_);
  nand _36396_ (_03582_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nand _36397_ (_23833_, _03582_, _03581_);
  not _36398_ (_03583_, _00376_);
  nand _36399_ (_03584_, _01278_, _03583_);
  nand _36400_ (_03585_, _03584_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _36401_ (_03586_, _03585_, _01293_);
  not _36402_ (_03587_, _01278_);
  nor _36403_ (_03588_, _26402_, _01426_);
  nor _36404_ (_03589_, _03588_, _00382_);
  nor _36405_ (_03591_, _03589_, _03587_);
  nor _36406_ (_03592_, _03591_, _03586_);
  nand _36407_ (_03593_, _01287_, _25029_);
  nand _36408_ (_03595_, _03593_, _26487_);
  nor _36409_ (_23834_, _03595_, _03592_);
  nor _36410_ (_03596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nand _36411_ (_03597_, _03596_, _01241_);
  not _36412_ (_03598_, _03597_);
  nand _36413_ (_03599_, _03598_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _36414_ (_03600_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand _36415_ (_03601_, _03600_, _03599_);
  nor _36416_ (_03602_, _03601_, _01278_);
  nand _36417_ (_03603_, _00275_, _24716_);
  not _36418_ (_03604_, _03603_);
  nand _36419_ (_03605_, _00276_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand _36420_ (_03607_, _03605_, _01278_);
  nor _36421_ (_03609_, _03607_, _03604_);
  nor _36422_ (_03611_, _03609_, _03602_);
  nor _36423_ (_03612_, _03611_, _01287_);
  nand _36424_ (_03613_, _01287_, _25703_);
  nand _36425_ (_03614_, _03613_, _26487_);
  nor _36426_ (_23835_, _03614_, _03612_);
  nor _36427_ (_03615_, _01253_, _01347_);
  not _36428_ (_03616_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _36429_ (_03617_, _01254_, _03616_);
  nor _36430_ (_03618_, _03617_, _03615_);
  nor _36431_ (_03619_, _03618_, _01261_);
  nand _36432_ (_03620_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand _36433_ (_03621_, _03620_, _01241_);
  nor _36434_ (_03623_, _03621_, _01260_);
  nor _36435_ (_03624_, _03623_, _03619_);
  nor _36436_ (_23836_, _03624_, rst);
  nor _36437_ (_03626_, _01303_, _25625_);
  nand _36438_ (_03627_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nand _36439_ (_03628_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nand _36440_ (_03629_, _03628_, _03627_);
  nand _36441_ (_03630_, _03629_, _01260_);
  nand _36442_ (_03631_, _01309_, _25139_);
  nand _36443_ (_03632_, _03631_, _03630_);
  nor _36444_ (_03633_, _03632_, _03626_);
  nor _36445_ (_23837_, _03633_, rst);
  not _36446_ (_03634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  nand _36447_ (_03635_, _00434_, _25628_);
  nand _36448_ (_03637_, _03635_, _03634_);
  nand _36449_ (_03638_, _03637_, _26487_);
  nor _36450_ (_03639_, _03635_, _25194_);
  nor _36451_ (_23838_, _03639_, _03638_);
  not _36452_ (_03640_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  nand _36453_ (_03641_, _03635_, _03640_);
  nand _36454_ (_03642_, _03641_, _26487_);
  nor _36455_ (_03643_, _03635_, _25089_);
  nor _36456_ (_23839_, _03643_, _03642_);
  not _36457_ (_03644_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  nand _36458_ (_03645_, _03635_, _03644_);
  nand _36459_ (_03646_, _03645_, _26487_);
  nor _36460_ (_03647_, _03635_, _24920_);
  nor _36461_ (_23840_, _03647_, _03646_);
  not _36462_ (_03649_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _36463_ (_03650_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _03355_);
  nand _36464_ (_03651_, _03650_, _01241_);
  nand _36465_ (_03652_, _03651_, _03596_);
  nand _36466_ (_03653_, _03652_, _03649_);
  nor _36467_ (_03654_, _03653_, _01278_);
  nand _36468_ (_03655_, _25722_, _24716_);
  not _36469_ (_03656_, _03655_);
  nand _36470_ (_03657_, _25723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _36471_ (_03658_, _03657_, _01278_);
  nor _36472_ (_03659_, _03658_, _03656_);
  nor _36473_ (_03660_, _03659_, _03654_);
  nor _36474_ (_03662_, _03660_, _01287_);
  nand _36475_ (_03664_, _01290_, _24820_);
  nand _36476_ (_03665_, _03664_, _26487_);
  nor _36477_ (_23841_, _03665_, _03662_);
  not _36478_ (_03666_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  nand _36479_ (_03667_, _03635_, _03666_);
  nand _36480_ (_03668_, _03667_, _26487_);
  nor _36481_ (_03669_, _03635_, _25028_);
  nor _36482_ (_23842_, _03669_, _03668_);
  nor _36483_ (_03670_, _03635_, _24821_);
  not _36484_ (_03671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand _36485_ (_03672_, _03635_, _03671_);
  nand _36486_ (_03673_, _03672_, _26487_);
  nor _36487_ (_23843_, _03673_, _03670_);
  nor _36488_ (_03674_, _01303_, _25140_);
  nand _36489_ (_03675_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nand _36490_ (_03676_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand _36491_ (_03678_, _03676_, _03675_);
  nand _36492_ (_03679_, _03678_, _01260_);
  nand _36493_ (_03680_, _01309_, _24920_);
  nand _36494_ (_03682_, _03680_, _03679_);
  nor _36495_ (_03684_, _03682_, _03674_);
  nor _36496_ (_23844_, _03684_, rst);
  not _36497_ (_03685_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand _36498_ (_03686_, _03635_, _03685_);
  nand _36499_ (_03687_, _03686_, _26487_);
  nor _36500_ (_03688_, _03635_, _25139_);
  nor _36501_ (_23845_, _03688_, _03687_);
  not _36502_ (_03689_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  nand _36503_ (_03690_, _03635_, _03689_);
  nand _36504_ (_03691_, _03690_, _26487_);
  nor _36505_ (_03692_, _03635_, _25680_);
  nor _36506_ (_23846_, _03692_, _03691_);
  nor _36507_ (_03693_, _01314_, _24782_);
  not _36508_ (_03694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nand _36509_ (_03695_, _01253_, _03694_);
  nand _36510_ (_03697_, _01254_, _03616_);
  nand _36511_ (_03698_, _03697_, _03695_);
  nand _36512_ (_03699_, _03698_, _01260_);
  nand _36513_ (_03701_, _03699_, _26487_);
  nor _36514_ (_23847_, _03701_, _03693_);
  nand _36515_ (_03702_, _03571_, _24789_);
  nand _36516_ (_03703_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  nand _36517_ (_23848_, _03703_, _03702_);
  nor _36518_ (_03704_, _00393_, _24993_);
  nand _36519_ (_03705_, _03704_, _28096_);
  not _36520_ (_03706_, _03704_);
  nand _36521_ (_03707_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nand _36522_ (_23849_, _03707_, _03705_);
  nand _36523_ (_03708_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  nand _36524_ (_23850_, _03708_, _01490_);
  nand _36525_ (_03709_, _01467_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not _36526_ (_03710_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  not _36527_ (_03711_, _01440_);
  nand _36528_ (_03713_, _03711_, _01430_);
  nand _36529_ (_03714_, _03713_, _03710_);
  nor _36530_ (_03715_, _01452_, _03711_);
  nor _36531_ (_03716_, _03715_, _01456_);
  nand _36532_ (_03717_, _03716_, _03714_);
  nand _36533_ (_03718_, _03717_, _03709_);
  nand _36534_ (_03719_, _03718_, _01415_);
  nand _36535_ (_23851_, _03719_, _01418_);
  nor _36536_ (_03720_, _01481_, _01445_);
  nor _36537_ (_03722_, _01479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _36538_ (_03724_, _03722_, _03720_);
  nor _36539_ (_23852_, _03724_, rst);
  nand _36540_ (_03725_, _00979_, _24789_);
  nand _36541_ (_03726_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  nand _36542_ (_23853_, _03726_, _03725_);
  nand _36543_ (_03727_, _25152_, _24830_);
  nand _36544_ (_03728_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  nand _36545_ (_23854_, _03728_, _03727_);
  nand _36546_ (_03729_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nand _36547_ (_03731_, _28074_, _25150_);
  nand _36548_ (_23855_, _03731_, _03729_);
  nor _36549_ (_03732_, _01445_, _01476_);
  nand _36550_ (_03734_, _03732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor _36551_ (_03735_, _03734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nand _36552_ (_03736_, _03735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _36553_ (_03737_, _03736_, _01435_);
  nor _36554_ (_03738_, _03737_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not _36555_ (_03739_, rxd_i);
  nand _36556_ (_03740_, _03737_, _03739_);
  nand _36557_ (_03741_, _03740_, _26487_);
  nor _36558_ (_23856_, _03741_, _03738_);
  nand _36559_ (_03742_, _03704_, _25203_);
  nand _36560_ (_03743_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nand _36561_ (_23857_, _03743_, _03742_);
  nor _36562_ (_03744_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  nand _36563_ (_03746_, _03744_, _01454_);
  nor _36564_ (_03748_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor _36565_ (_03749_, _03748_, _01460_);
  nand _36566_ (_03750_, _03749_, _03746_);
  nand _36567_ (_23858_, _03750_, _01420_);
  nand _36568_ (_03751_, _03732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nand _36569_ (_03752_, _03734_, _01434_);
  nor _36570_ (_03753_, _03752_, _03751_);
  nor _36571_ (_03755_, _03753_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nand _36572_ (_03756_, _03752_, _01481_);
  nand _36573_ (_03757_, _03756_, _26487_);
  nor _36574_ (_23859_, _03757_, _03755_);
  nand _36575_ (_03759_, _03704_, _24927_);
  nand _36576_ (_03760_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  nand _36577_ (_23860_, _03760_, _03759_);
  nand _36578_ (_03761_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand _36579_ (_03762_, _01467_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _36580_ (_03763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor _36581_ (_03764_, _01456_, _03763_);
  nand _36582_ (_03765_, _03764_, _01454_);
  nand _36583_ (_03766_, _03765_, _03762_);
  nand _36584_ (_03767_, _03766_, _01415_);
  nand _36585_ (_23861_, _03767_, _03761_);
  nor _36586_ (_03768_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  nand _36587_ (_03769_, _03768_, _01454_);
  nor _36588_ (_03770_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  nor _36589_ (_03771_, _03770_, _01460_);
  nand _36590_ (_03772_, _03771_, _03769_);
  nand _36591_ (_23862_, _03772_, _01422_);
  nand _36592_ (_03773_, _00479_, _25039_);
  nand _36593_ (_03774_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  nand _36594_ (_23863_, _03774_, _03773_);
  nand _36595_ (_03775_, _25166_, _25099_);
  nand _36596_ (_03777_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nand _36597_ (_23864_, _03777_, _03775_);
  nand _36598_ (_03778_, _28096_, _25166_);
  nand _36599_ (_03779_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nand _36600_ (_23865_, _03779_, _03778_);
  nand _36601_ (_03780_, _03704_, _24789_);
  nand _36602_ (_03781_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  nand _36603_ (_23866_, _03781_, _03780_);
  nor _36604_ (_03782_, _00954_, _24993_);
  nand _36605_ (_03783_, _03782_, _25099_);
  not _36606_ (_03785_, _03782_);
  nand _36607_ (_03786_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nand _36608_ (_23867_, _03786_, _03783_);
  nand _36609_ (_03787_, _01182_, _28096_);
  nand _36610_ (_03788_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  nand _36611_ (_23868_, _03788_, _03787_);
  nand _36612_ (_03789_, _03782_, _28096_);
  nand _36613_ (_03790_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  nand _36614_ (_23869_, _03790_, _03789_);
  nand _36615_ (_03791_, _03782_, _25039_);
  nand _36616_ (_03792_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  nand _36617_ (_23930_, _03792_, _03791_);
  nand _36618_ (_03793_, _03782_, _25150_);
  nand _36619_ (_03794_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nand _36620_ (_23947_, _03794_, _03793_);
  nand _36621_ (_03795_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nand _36622_ (_03796_, _03547_, _24927_);
  nand _36623_ (_23949_, _03796_, _03795_);
  nand _36624_ (_03797_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nand _36625_ (_03798_, _03547_, _25039_);
  nand _36626_ (_23983_, _03798_, _03797_);
  nand _36627_ (_03800_, _01905_, _24927_);
  nand _36628_ (_03801_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nand _36629_ (_24008_, _03801_, _03800_);
  nand _36630_ (_03803_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nand _36631_ (_03804_, _03547_, _25203_);
  nand _36632_ (_24011_, _03804_, _03803_);
  nand _36633_ (_03805_, _01905_, _25039_);
  nand _36634_ (_03806_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nand _36635_ (_24022_, _03806_, _03805_);
  nand _36636_ (_03807_, _24852_, _24789_);
  nand _36637_ (_03808_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  nand _36638_ (_24101_, _03808_, _03807_);
  nand _36639_ (_03809_, _00991_, _28096_);
  nand _36640_ (_03810_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  nand _36641_ (_24107_, _03810_, _03809_);
  nor _36642_ (_03811_, _00629_, _25159_);
  nand _36643_ (_03812_, _03811_, _24789_);
  not _36644_ (_03813_, _03811_);
  nand _36645_ (_03814_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand _36646_ (_24134_, _03814_, _03812_);
  nand _36647_ (_03815_, _03811_, _25150_);
  nand _36648_ (_03816_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nand _36649_ (_24141_, _03816_, _03815_);
  nand _36650_ (_03817_, _03811_, _24927_);
  nand _36651_ (_03818_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nand _36652_ (_24168_, _03818_, _03817_);
  nand _36653_ (_03819_, _03811_, _25039_);
  nand _36654_ (_03820_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nand _36655_ (_24219_, _03820_, _03819_);
  nor _36656_ (_03822_, _00631_, _24999_);
  nand _36657_ (_03824_, _03822_, _28096_);
  not _36658_ (_03825_, _03822_);
  nand _36659_ (_03826_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nand _36660_ (_24233_, _03826_, _03824_);
  nand _36661_ (_03827_, _03822_, _25039_);
  nand _36662_ (_03828_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  nand _36663_ (_24238_, _03828_, _03827_);
  nor _36664_ (_03829_, _03546_, _24795_);
  not _36665_ (_03830_, _03829_);
  nand _36666_ (_03831_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  nand _36667_ (_03832_, _03829_, _25039_);
  nand _36668_ (_24246_, _03832_, _03831_);
  nor _36669_ (_03834_, _00629_, _25059_);
  nand _36670_ (_03835_, _03834_, _24789_);
  not _36671_ (_03836_, _03834_);
  nand _36672_ (_03837_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  nand _36673_ (_24291_, _03837_, _03835_);
  nand _36674_ (_03838_, _25203_, _25166_);
  nand _36675_ (_03839_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nand _36676_ (_24307_, _03839_, _03838_);
  nor _36677_ (_03840_, _00631_, _24882_);
  nand _36678_ (_03841_, _03840_, _24830_);
  not _36679_ (_03842_, _03840_);
  nand _36680_ (_03843_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nand _36681_ (_24341_, _03843_, _03841_);
  nand _36682_ (_03844_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nand _36683_ (_03845_, _03829_, _25203_);
  nand _36684_ (_24399_, _03845_, _03844_);
  nand _36685_ (_03846_, _03822_, _24830_);
  nand _36686_ (_03847_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nand _36687_ (_24487_, _03847_, _03846_);
  nand _36688_ (_03848_, _00955_, _25150_);
  nand _36689_ (_03849_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nand _36690_ (_24503_, _03849_, _03848_);
  nor _36691_ (_03850_, _25165_, _28080_);
  nand _36692_ (_03851_, _03850_, _25203_);
  not _36693_ (_03852_, _03850_);
  nand _36694_ (_03853_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  nand _36695_ (_24526_, _03853_, _03851_);
  nand _36696_ (_03854_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  nand _36697_ (_03855_, _03829_, _24927_);
  nand _36698_ (_24572_, _03855_, _03854_);
  nand _36699_ (_03856_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  nand _36700_ (_03857_, _03829_, _24789_);
  nand _36701_ (_24587_, _03857_, _03856_);
  nor _36702_ (_03858_, _00631_, _28073_);
  nand _36703_ (_03859_, _03858_, _25099_);
  not _36704_ (_03861_, _03858_);
  nand _36705_ (_03862_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  nand _36706_ (_24596_, _03862_, _03859_);
  nand _36707_ (_03865_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  nand _36708_ (_03866_, _03829_, _25150_);
  nand _36709_ (_24598_, _03866_, _03865_);
  nor _36710_ (_03867_, _00629_, _25051_);
  not _36711_ (_03868_, _03867_);
  nand _36712_ (_03869_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  nand _36713_ (_03870_, _03867_, _24830_);
  nand _36714_ (_24608_, _03870_, _03869_);
  nand _36715_ (_03871_, _03811_, _24830_);
  nand _36716_ (_03872_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand _36717_ (_24615_, _03872_, _03871_);
  nand _36718_ (_03873_, _00115_, _24830_);
  nand _36719_ (_03874_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nand _36720_ (_24652_, _03874_, _03873_);
  nor _36721_ (_03876_, _00393_, _25165_);
  nand _36722_ (_03877_, _03876_, _25203_);
  not _36723_ (_03878_, _03876_);
  nand _36724_ (_03879_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  nand _36725_ (_24660_, _03879_, _03877_);
  nand _36726_ (_03880_, _00632_, _24927_);
  nand _36727_ (_03881_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  nand _36728_ (_24662_, _03881_, _03880_);
  nand _36729_ (_03882_, _03876_, _25039_);
  nand _36730_ (_03883_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nand _36731_ (_24800_, _03883_, _03882_);
  nor _36732_ (_03884_, _03546_, _24059_);
  not _36733_ (_03886_, _03884_);
  nand _36734_ (_03888_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  nand _36735_ (_03889_, _03884_, _24927_);
  nand _36736_ (_24825_, _03889_, _03888_);
  nand _36737_ (_03890_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  nand _36738_ (_03891_, _03884_, _24789_);
  nand _36739_ (_24828_, _03891_, _03890_);
  nand _36740_ (_03892_, _03811_, _25203_);
  nand _36741_ (_03893_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nand _36742_ (_24834_, _03893_, _03892_);
  nor _36743_ (_03894_, _24984_, _24059_);
  nand _36744_ (_03895_, _03894_, _24927_);
  not _36745_ (_03896_, _03894_);
  nand _36746_ (_03897_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  nand _36747_ (_24841_, _03897_, _03895_);
  nand _36748_ (_03898_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nand _36749_ (_03900_, _03884_, _25150_);
  nand _36750_ (_24844_, _03900_, _03898_);
  nand _36751_ (_03902_, _03811_, _28096_);
  nand _36752_ (_03903_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand _36753_ (_24851_, _03903_, _03902_);
  nand _36754_ (_03904_, _03811_, _25099_);
  nand _36755_ (_03905_, _03813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand _36756_ (_24854_, _03905_, _03904_);
  nand _36757_ (_03906_, _00394_, _25203_);
  nand _36758_ (_03907_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  nand _36759_ (_24857_, _03907_, _03906_);
  nand _36760_ (_03908_, _03822_, _25203_);
  nand _36761_ (_03910_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  nand _36762_ (_24875_, _03910_, _03908_);
  nor _36763_ (_03911_, _28073_, _25165_);
  nand _36764_ (_03912_, _03911_, _24830_);
  not _36765_ (_03913_, _03911_);
  nand _36766_ (_03914_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nand _36767_ (_24880_, _03914_, _03912_);
  not _36768_ (_03915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _36769_ (_03916_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _03915_);
  not _36770_ (_03917_, _03368_);
  nand _36771_ (_03918_, _03917_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor _36772_ (_03919_, _03918_, _03380_);
  nor _36773_ (_03920_, _03919_, _00556_);
  nor _36774_ (_03921_, _03920_, _03916_);
  nor _36775_ (_03923_, _00135_, _23938_);
  nand _36776_ (_03924_, _03923_, _25628_);
  not _36777_ (_03925_, _03924_);
  nand _36778_ (_03926_, _03925_, _26244_);
  nand _36779_ (_03928_, _03926_, _03921_);
  nand _36780_ (_03929_, _03928_, _00622_);
  nor _36781_ (_03930_, _03926_, _24716_);
  nor _36782_ (_03931_, _03930_, _03929_);
  nor _36783_ (_03932_, _00622_, _26096_);
  nor _36784_ (_03933_, _03932_, _03931_);
  nor _36785_ (_24915_, _03933_, rst);
  nor _36786_ (_03934_, _00131_, _24836_);
  not _36787_ (_03935_, _03934_);
  nor _36788_ (_03936_, _03935_, _01549_);
  nand _36789_ (_03937_, _03936_, _24849_);
  nor _36790_ (_03938_, _03937_, _25194_);
  not _36791_ (_03939_, _03937_);
  nor _36792_ (_03940_, _03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _36793_ (_24937_, _03940_, _03938_);
  nor _36794_ (_03942_, _03937_, _24920_);
  nor _36795_ (_03943_, _03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _36796_ (_24943_, _03943_, _03942_);
  not _36797_ (_03944_, _00297_);
  nor _36798_ (_03945_, _00287_, _25194_);
  nand _36799_ (_03946_, _00272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand _36800_ (_03947_, _00271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nand _36801_ (_03948_, _03947_, _03946_);
  nor _36802_ (_03949_, _03948_, _00279_);
  nor _36803_ (_03951_, _03949_, _03945_);
  nor _36804_ (_03952_, _03951_, _03944_);
  not _36805_ (_03953_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand _36806_ (_03954_, _03944_, _03953_);
  nand _36807_ (_03955_, _03954_, _26487_);
  nor _36808_ (_24948_, _03955_, _03952_);
  nor _36809_ (_03956_, _03937_, _25028_);
  nor _36810_ (_03957_, _03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _36811_ (_24952_, _03957_, _03956_);
  nor _36812_ (_03958_, _00415_, _28057_);
  nand _36813_ (_03959_, _03958_, _24927_);
  not _36814_ (_03960_, _03958_);
  nand _36815_ (_03961_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  nand _36816_ (_24967_, _03961_, _03959_);
  nand _36817_ (_03962_, _00991_, _25099_);
  nand _36818_ (_03964_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  nand _36819_ (_24974_, _03964_, _03962_);
  nand _36820_ (_03966_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nand _36821_ (_03967_, _03829_, _25099_);
  nand _36822_ (_24980_, _03967_, _03966_);
  nand _36823_ (_03968_, _00115_, _28096_);
  nand _36824_ (_03969_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nand _36825_ (_25016_, _03969_, _03968_);
  nor _36826_ (_03971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _36827_ (_03973_, _03971_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _36828_ (_03974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand _36829_ (_03975_, _03375_, _03374_);
  nor _36830_ (_03976_, _03975_, _03918_);
  nor _36831_ (_03977_, _03976_, _03974_);
  nor _36832_ (_03978_, _03977_, _03973_);
  nor _36833_ (_03979_, _26245_, _23938_);
  nand _36834_ (_03980_, _03979_, _25628_);
  not _36835_ (_03981_, _03980_);
  nand _36836_ (_03983_, _03981_, _26135_);
  nand _36837_ (_03985_, _03983_, _03978_);
  nand _36838_ (_03986_, _03985_, _00622_);
  nor _36839_ (_03987_, _03983_, _24716_);
  nor _36840_ (_03988_, _03987_, _03986_);
  nor _36841_ (_03989_, _00622_, _25625_);
  nor _36842_ (_03990_, _03989_, _03988_);
  nor _36843_ (_25019_, _03990_, rst);
  nand _36844_ (_03991_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  nand _36845_ (_03992_, _03829_, _24830_);
  nand _36846_ (_25035_, _03992_, _03991_);
  nand _36847_ (_03994_, _28063_, _25150_);
  nand _36848_ (_03995_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  nand _36849_ (_25041_, _03995_, _03994_);
  nor _36850_ (_03998_, _03937_, _24782_);
  nor _36851_ (_03999_, _03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _36852_ (_25060_, _03999_, _03998_);
  nand _36853_ (_04000_, _03834_, _25150_);
  nand _36854_ (_04001_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nand _36855_ (_25064_, _04001_, _04000_);
  nor _36856_ (_04003_, _03937_, _25139_);
  nor _36857_ (_04005_, _03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _36858_ (_25077_, _04005_, _04003_);
  nor _36859_ (_04006_, _00954_, _24889_);
  nand _36860_ (_04007_, _04006_, _25150_);
  not _36861_ (_04008_, _04006_);
  nand _36862_ (_04009_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nand _36863_ (_25090_, _04009_, _04007_);
  nand _36864_ (_04011_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  nand _36865_ (_04012_, _03884_, _25099_);
  nand _36866_ (_25100_, _04012_, _04011_);
  nand _36867_ (_04013_, _25000_, _24789_);
  nand _36868_ (_04014_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  nand _36869_ (_25105_, _04014_, _04013_);
  nor _36870_ (_04015_, _25051_, _28080_);
  not _36871_ (_04016_, _04015_);
  nand _36872_ (_04017_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nand _36873_ (_04018_, _04015_, _25150_);
  nand _36874_ (_25117_, _04018_, _04017_);
  nand _36875_ (_04019_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nand _36876_ (_04020_, _03884_, _24830_);
  nand _36877_ (_25120_, _04020_, _04019_);
  nor _36878_ (_04021_, _25051_, _24882_);
  not _36879_ (_04022_, _04021_);
  nand _36880_ (_04023_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nand _36881_ (_04024_, _04021_, _28096_);
  nand _36882_ (_25124_, _04024_, _04023_);
  nand _36883_ (_04025_, _00479_, _24830_);
  nand _36884_ (_04026_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  nand _36885_ (_25142_, _04026_, _04025_);
  nand _36886_ (_04027_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nand _36887_ (_04028_, _03867_, _25099_);
  nand _36888_ (_25184_, _04028_, _04027_);
  nor _36889_ (_04030_, _03937_, _24820_);
  not _36890_ (_04031_, _04030_);
  nand _36891_ (_04033_, _03937_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nand _36892_ (_25211_, _04033_, _04031_);
  nand _36893_ (_04034_, _03850_, _28096_);
  nand _36894_ (_04035_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  nand _36895_ (_25221_, _04035_, _04034_);
  nor _36896_ (_04036_, _25395_, _25235_);
  nor _36897_ (_04037_, _25395_, _25298_);
  nor _36898_ (_04038_, _26195_, _25416_);
  nor _36899_ (_04040_, _04038_, _04037_);
  not _36900_ (_04041_, _04040_);
  nor _36901_ (_04042_, _04041_, _04036_);
  nor _36902_ (_04043_, _26202_, _25395_);
  nor _36903_ (_04044_, _04043_, _25417_);
  nand _36904_ (_04045_, _04044_, _04042_);
  nor _36905_ (_04046_, _26202_, _25470_);
  nor _36906_ (_04047_, _04046_, _04045_);
  nor _36907_ (_04048_, _04047_, _24864_);
  not _36908_ (_04050_, _25804_);
  nor _36909_ (_04052_, _04050_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _36910_ (_04053_, _25805_);
  nor _36911_ (_04054_, _04053_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _36912_ (_04055_, _04054_, _04052_);
  nand _36913_ (_04056_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _36914_ (_04057_, _04056_, _04055_);
  nor _36915_ (_04058_, _04057_, _04048_);
  nor _36916_ (_28194_[1], _04058_, rst);
  nand _36917_ (_04059_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  nand _36918_ (_04060_, _03884_, _25203_);
  nand _36919_ (_25247_, _04060_, _04059_);
  nand _36920_ (_04061_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nand _36921_ (_04062_, _03884_, _28096_);
  nand _36922_ (_25257_, _04062_, _04061_);
  nand _36923_ (_04063_, _03894_, _25203_);
  nand _36924_ (_04065_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  nand _36925_ (_25302_, _04065_, _04063_);
  nand _36926_ (_04066_, _28063_, _24789_);
  nand _36927_ (_04067_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  nand _36928_ (_25429_, _04067_, _04066_);
  not _36929_ (_04068_, _25579_);
  nor _36930_ (_04069_, _01022_, _04068_);
  not _36931_ (_04070_, _04069_);
  not _36932_ (_04071_, _25602_);
  nor _36933_ (_04072_, _25426_, _25482_);
  nor _36934_ (_04074_, _04072_, _04071_);
  not _36935_ (_04076_, _25567_);
  nor _36936_ (_04078_, _25565_, _25327_);
  nor _36937_ (_04079_, _04078_, _04076_);
  nand _36938_ (_04080_, _04079_, _04074_);
  nor _36939_ (_04081_, _04080_, _04070_);
  not _36940_ (_04082_, _04081_);
  nand _36941_ (_04083_, _25544_, _25535_);
  nor _36942_ (_04084_, _04083_, _04082_);
  nor _36943_ (_04085_, _04084_, _25530_);
  not _36944_ (_04086_, _25541_);
  nor _36945_ (_04087_, _04086_, _25537_);
  nor _36946_ (_04088_, _04087_, _25505_);
  nor _36947_ (_04089_, _04088_, _04085_);
  nor _36948_ (_28234_, _04089_, rst);
  nand _36949_ (_04090_, _03937_, _25769_);
  nand _36950_ (_04091_, _04090_, _26487_);
  nor _36951_ (_28196_[7], _04091_, _03998_);
  nor _36952_ (_04093_, _03935_, _25629_);
  not _36953_ (_04094_, _04093_);
  nor _36954_ (_04095_, _04094_, _25625_);
  nand _36955_ (_04096_, _04094_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nand _36956_ (_04097_, _04096_, _24849_);
  nor _36957_ (_04098_, _04097_, _04095_);
  nand _36958_ (_04099_, _24850_, _25764_);
  nand _36959_ (_04101_, _04099_, _26487_);
  nor _36960_ (_28197_[7], _04101_, _04098_);
  nor _36961_ (_04103_, _03935_, _00233_);
  nand _36962_ (_04104_, _04103_, _24849_);
  nor _36963_ (_04105_, _04104_, _24782_);
  nand _36964_ (_04106_, _04104_, _25759_);
  nand _36965_ (_04107_, _04106_, _26487_);
  nor _36966_ (_28198_[7], _04107_, _04105_);
  nor _36967_ (_04109_, _03935_, _24845_);
  not _36968_ (_04110_, _04109_);
  nor _36969_ (_04111_, _04110_, _24850_);
  not _36970_ (_04113_, _04111_);
  nor _36971_ (_04114_, _04113_, _25625_);
  nor _36972_ (_04116_, _04111_, _25789_);
  nor _36973_ (_04117_, _04116_, _04114_);
  nor _36974_ (_28199_[7], _04117_, rst);
  nor _36975_ (_04118_, _01549_, _24838_);
  nor _36976_ (_04119_, _04093_, _03936_);
  nor _36977_ (_04120_, _04109_, _04103_);
  nand _36978_ (_04121_, _04120_, _04119_);
  nor _36979_ (_04122_, _04121_, _04118_);
  nor _36980_ (_04123_, _04122_, _24850_);
  not _36981_ (_04125_, _04123_);
  nor _36982_ (_04127_, _04125_, _03936_);
  nor _36983_ (_04129_, _04127_, _25778_);
  not _36984_ (_04130_, _04118_);
  nor _36985_ (_04131_, _04130_, _25625_);
  not _36986_ (_04132_, _04120_);
  nor _36987_ (_04133_, _04132_, _04093_);
  nor _36988_ (_04134_, _04133_, _25778_);
  nor _36989_ (_04136_, _04134_, _04131_);
  nor _36990_ (_04138_, _04136_, _24850_);
  nor _36991_ (_04139_, _04138_, _04129_);
  nor _36992_ (_28200_[7], _04139_, rst);
  nor _36993_ (_04140_, _25629_, _24838_);
  nand _36994_ (_04141_, _04140_, _24849_);
  nor _36995_ (_04142_, _04141_, _25625_);
  not _36996_ (_04144_, _04122_);
  nor _36997_ (_04145_, _04144_, _04140_);
  nor _36998_ (_04146_, _04145_, _24850_);
  nand _36999_ (_04148_, _04146_, _04119_);
  nor _37000_ (_04149_, _04132_, _04118_);
  nor _37001_ (_04150_, _04149_, _24850_);
  nor _37002_ (_04151_, _04150_, _04148_);
  nor _37003_ (_04152_, _04151_, _25773_);
  nor _37004_ (_04153_, _04152_, _04142_);
  nor _37005_ (_28201_[7], _04153_, rst);
  nor _37006_ (_04154_, _00233_, _24838_);
  not _37007_ (_04155_, _04154_);
  nor _37008_ (_04156_, _04155_, _24850_);
  not _37009_ (_04157_, _04156_);
  nor _37010_ (_04158_, _04157_, _25625_);
  nor _37011_ (_04159_, _04156_, _25786_);
  nor _37012_ (_04160_, _04159_, _04158_);
  nor _37013_ (_28202_[7], _04160_, rst);
  nor _37014_ (_04162_, _24855_, _25625_);
  nor _37015_ (_04163_, _24852_, _25781_);
  nor _37016_ (_04165_, _04163_, _04162_);
  nor _37017_ (_28203_[7], _04165_, rst);
  nor _37018_ (_04166_, _03546_, _24978_);
  not _37019_ (_04167_, _04166_);
  nand _37020_ (_04168_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nand _37021_ (_04169_, _04166_, _28096_);
  nand _37022_ (_25525_, _04169_, _04168_);
  nand _37023_ (_04170_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  nand _37024_ (_04171_, _04166_, _25099_);
  nand _37025_ (_25536_, _04171_, _04170_);
  nor _37026_ (_04172_, _00149_, _25627_);
  not _37027_ (_04173_, _04172_);
  nor _37028_ (_04174_, _04173_, _25139_);
  not _37029_ (_04175_, _01573_);
  not _37030_ (_04176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _37031_ (_04177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _37032_ (_04178_, _04177_, _04176_);
  not _37033_ (_04180_, _04178_);
  not _37034_ (_04181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _37035_ (_04182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  not _37036_ (_04183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _37037_ (_04185_, _01575_, _04183_);
  not _37038_ (_04186_, _04185_);
  nor _37039_ (_04187_, _04186_, _04182_);
  not _37040_ (_04188_, _04187_);
  nor _37041_ (_04189_, _04188_, _04181_);
  not _37042_ (_04191_, _04189_);
  nor _37043_ (_04192_, _04191_, _01605_);
  not _37044_ (_04193_, _04192_);
  nor _37045_ (_04194_, _04193_, _04180_);
  not _37046_ (_04195_, _04194_);
  nor _37047_ (_04196_, _04195_, _01608_);
  nor _37048_ (_04198_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _37049_ (_04199_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _37050_ (_04201_, _04199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _37051_ (_04203_, _04201_, _04198_);
  nor _37052_ (_04204_, _04191_, _04180_);
  not _37053_ (_04205_, _04204_);
  nor _37054_ (_04206_, _04205_, _01597_);
  nand _37055_ (_04207_, _04206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _37056_ (_04208_, _01574_);
  nor _37057_ (_04209_, _04206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _37058_ (_04210_, _04209_, _04208_);
  nand _37059_ (_04212_, _04210_, _04207_);
  not _37060_ (_04214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _37061_ (_04215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _37062_ (_04217_, _01597_, _01619_);
  not _37063_ (_04219_, _04217_);
  nor _37064_ (_04220_, _04219_, _04215_);
  nand _37065_ (_04221_, _04220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _37066_ (_04222_, _04221_);
  nand _37067_ (_04223_, _04222_, _04204_);
  nand _37068_ (_04225_, _04223_, _04214_);
  not _37069_ (_04226_, _01615_);
  nor _37070_ (_04228_, _04215_, _01618_);
  nand _37071_ (_04230_, _04217_, _04228_);
  nor _37072_ (_04231_, _04205_, _04214_);
  not _37073_ (_04232_, _04231_);
  nor _37074_ (_04233_, _04232_, _04230_);
  nor _37075_ (_04234_, _04233_, _04226_);
  nand _37076_ (_04235_, _04234_, _04225_);
  nand _37077_ (_04236_, _04235_, _04212_);
  nor _37078_ (_04237_, _04236_, _04203_);
  nand _37079_ (_04238_, _04237_, _04173_);
  nand _37080_ (_04240_, _04238_, _04175_);
  nor _37081_ (_04242_, _04240_, _04174_);
  nor _37082_ (_04243_, _04175_, _04214_);
  nor _37083_ (_04244_, _04243_, _04242_);
  nor _37084_ (_25539_, _04244_, rst);
  nand _37085_ (_04245_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nand _37086_ (_04246_, _04166_, _24830_);
  nand _37087_ (_25543_, _04246_, _04245_);
  nand _37088_ (_04247_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  nand _37089_ (_04248_, _04166_, _25039_);
  nand _37090_ (_25667_, _04248_, _04247_);
  nand _37091_ (_04249_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  nand _37092_ (_04250_, _04166_, _24927_);
  nand _37093_ (_25763_, _04250_, _04249_);
  nor _37094_ (_04251_, _00926_, _24984_);
  nand _37095_ (_04252_, _04251_, _25150_);
  not _37096_ (_04253_, _04251_);
  nand _37097_ (_04254_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  nand _37098_ (_25875_, _04254_, _04252_);
  nor _37099_ (_04255_, _03546_, _24999_);
  not _37100_ (_04257_, _04255_);
  nand _37101_ (_04258_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  nand _37102_ (_04259_, _04255_, _24927_);
  nand _37103_ (_25878_, _04259_, _04258_);
  nand _37104_ (_04261_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  nand _37105_ (_04262_, _04255_, _24789_);
  nand _37106_ (_26022_, _04262_, _04261_);
  nor _37107_ (_04264_, _00122_, _25051_);
  not _37108_ (_04265_, _04264_);
  nand _37109_ (_04266_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nand _37110_ (_04267_, _04264_, _25099_);
  nand _37111_ (_26116_, _04267_, _04266_);
  nor _37112_ (_04269_, _24972_, _24862_);
  not _37113_ (_04270_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nand _37114_ (_04271_, _24862_, _04270_);
  nand _37115_ (_04273_, _04271_, _26487_);
  nor _37116_ (_28186_[6], _04273_, _04269_);
  nand _37117_ (_04274_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  nand _37118_ (_04275_, _04255_, _24830_);
  nand _37119_ (_26128_, _04275_, _04274_);
  nor _37120_ (_04276_, _25470_, _25482_);
  nor _37121_ (_04277_, _04276_, _25467_);
  not _37122_ (_04279_, _04277_);
  nor _37123_ (_04280_, _26202_, _25577_);
  not _37124_ (_04282_, _04280_);
  nand _37125_ (_04283_, _04282_, _01051_);
  nor _37126_ (_04285_, _04283_, _04279_);
  nor _37127_ (_04286_, _04285_, _24864_);
  not _37128_ (_04288_, _00101_);
  nand _37129_ (_04289_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _37130_ (_04290_, _04289_, _04288_);
  nor _37131_ (_04291_, _04290_, _04286_);
  nor _37132_ (_28188_[1], _04291_, rst);
  nand _37133_ (_04292_, _25166_, _25150_);
  nand _37134_ (_04293_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  nand _37135_ (_26181_, _04293_, _04292_);
  nand _37136_ (_04296_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  nand _37137_ (_04298_, _04255_, _28096_);
  nand _37138_ (_26219_, _04298_, _04296_);
  nor _37139_ (_04299_, _03546_, _25057_);
  not _37140_ (_04301_, _04299_);
  nand _37141_ (_04302_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  nand _37142_ (_04303_, _04299_, _25039_);
  nand _37143_ (_26280_, _04303_, _04302_);
  nand _37144_ (_04304_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  nand _37145_ (_04305_, _04299_, _24927_);
  nand _37146_ (_26297_, _04305_, _04304_);
  nand _37147_ (_04306_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nand _37148_ (_04307_, _01388_, _25099_);
  nand _37149_ (_26308_, _04307_, _04306_);
  nor _37150_ (_04308_, _00631_, _25057_);
  nand _37151_ (_04309_, _04308_, _24789_);
  not _37152_ (_04310_, _04308_);
  nand _37153_ (_04311_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  nand _37154_ (_26316_, _04311_, _04309_);
  nor _37155_ (_04312_, _25057_, _24993_);
  nand _37156_ (_04313_, _04312_, _25039_);
  not _37157_ (_04314_, _04312_);
  nand _37158_ (_04315_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  nand _37159_ (_26321_, _04315_, _04313_);
  nand _37160_ (_04316_, _01153_, _24789_);
  nand _37161_ (_04317_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  nand _37162_ (_26327_, _04317_, _04316_);
  nand _37163_ (_04318_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  nand _37164_ (_04319_, _04299_, _25150_);
  nand _37165_ (_26336_, _04319_, _04318_);
  nand _37166_ (_04320_, _00394_, _24927_);
  nand _37167_ (_04321_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  nand _37168_ (_26446_, _04321_, _04320_);
  nor _37169_ (_04322_, _03546_, _28080_);
  not _37170_ (_04323_, _04322_);
  nand _37171_ (_04324_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  nand _37172_ (_04325_, _04322_, _24789_);
  nand _37173_ (_26462_, _04325_, _04324_);
  nand _37174_ (_04326_, _25203_, _25000_);
  nand _37175_ (_04327_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nand _37176_ (_26479_, _04327_, _04326_);
  nand _37177_ (_04328_, _00115_, _25203_);
  nand _37178_ (_04329_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  nand _37179_ (_26497_, _04329_, _04328_);
  nand _37180_ (_04331_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  nand _37181_ (_04332_, _04299_, _25099_);
  nand _37182_ (_26516_, _04332_, _04331_);
  nor _37183_ (_04333_, _03939_, _26287_);
  nor _37184_ (_04335_, _04333_, _04030_);
  nor _37185_ (_28196_[0], _04335_, rst);
  nor _37186_ (_04336_, _03937_, _25089_);
  nand _37187_ (_04337_, _03937_, _26448_);
  nand _37188_ (_04338_, _04337_, _26487_);
  nor _37189_ (_28196_[1], _04338_, _04336_);
  nor _37190_ (_04340_, _03937_, _25680_);
  nand _37191_ (_04341_, _03937_, _26354_);
  nand _37192_ (_04342_, _04341_, _26487_);
  nor _37193_ (_28196_[2], _04342_, _04340_);
  nand _37194_ (_04344_, _03937_, _25858_);
  nand _37195_ (_04346_, _04344_, _26487_);
  nor _37196_ (_28196_[3], _04346_, _03938_);
  nand _37197_ (_04347_, _03937_, _26020_);
  nand _37198_ (_04348_, _04347_, _26487_);
  nor _37199_ (_28196_[4], _04348_, _03956_);
  nand _37200_ (_04350_, _03937_, _26079_);
  nand _37201_ (_04352_, _04350_, _26487_);
  nor _37202_ (_28196_[5], _04352_, _03942_);
  nand _37203_ (_04354_, _03937_, _25953_);
  nand _37204_ (_04356_, _04354_, _26487_);
  nor _37205_ (_28196_[6], _04356_, _04003_);
  nand _37206_ (_04358_, _24849_, _24821_);
  nor _37207_ (_04360_, _04358_, _04094_);
  nor _37208_ (_04362_, _04094_, _24850_);
  nor _37209_ (_04363_, _04362_, _26284_);
  nor _37210_ (_04366_, _04363_, _04360_);
  nor _37211_ (_28197_[0], _04366_, rst);
  nor _37212_ (_04367_, _25088_, _04094_);
  nand _37213_ (_04369_, _04094_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand _37214_ (_04370_, _04369_, _24849_);
  nor _37215_ (_04371_, _04370_, _04367_);
  nand _37216_ (_04372_, _24850_, _26444_);
  nand _37217_ (_04373_, _04372_, _26487_);
  nor _37218_ (_28197_[1], _04373_, _04371_);
  nor _37219_ (_04375_, _25703_, _04094_);
  nand _37220_ (_04376_, _04094_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nand _37221_ (_04377_, _04376_, _24849_);
  nor _37222_ (_04378_, _04377_, _04375_);
  nand _37223_ (_04379_, _24850_, _26352_);
  nand _37224_ (_04380_, _04379_, _26487_);
  nor _37225_ (_28197_[2], _04380_, _04378_);
  nor _37226_ (_04382_, _25195_, _04094_);
  nand _37227_ (_04383_, _04094_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nand _37228_ (_04384_, _04383_, _24849_);
  nor _37229_ (_04385_, _04384_, _04382_);
  nand _37230_ (_04386_, _24850_, _25864_);
  nand _37231_ (_04387_, _04386_, _26487_);
  nor _37232_ (_28197_[3], _04387_, _04385_);
  nor _37233_ (_04389_, _25029_, _04094_);
  nand _37234_ (_04390_, _04094_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nand _37235_ (_04391_, _04390_, _24849_);
  nor _37236_ (_04392_, _04391_, _04389_);
  nand _37237_ (_04393_, _24850_, _26037_);
  nand _37238_ (_04394_, _04393_, _26487_);
  nor _37239_ (_28197_[4], _04394_, _04392_);
  nor _37240_ (_04395_, _26096_, _04094_);
  nand _37241_ (_04396_, _04094_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nand _37242_ (_04397_, _04396_, _24849_);
  nor _37243_ (_04398_, _04397_, _04395_);
  nand _37244_ (_04399_, _24850_, _26077_);
  nand _37245_ (_04400_, _04399_, _26487_);
  nor _37246_ (_28197_[5], _04400_, _04398_);
  nor _37247_ (_04401_, _25140_, _04094_);
  nand _37248_ (_04402_, _04094_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nand _37249_ (_04403_, _04402_, _24849_);
  nor _37250_ (_04405_, _04403_, _04401_);
  nand _37251_ (_04407_, _24850_, _25951_);
  nand _37252_ (_04409_, _04407_, _26487_);
  nor _37253_ (_28197_[6], _04409_, _04405_);
  not _37254_ (_04410_, _04104_);
  nor _37255_ (_04411_, _04410_, _26282_);
  nor _37256_ (_04412_, _04104_, _24820_);
  nor _37257_ (_04413_, _04412_, _04411_);
  nor _37258_ (_28198_[0], _04413_, rst);
  nor _37259_ (_04415_, _04104_, _25088_);
  nor _37260_ (_04416_, _04410_, _26442_);
  nor _37261_ (_04418_, _04416_, _04415_);
  nor _37262_ (_28198_[1], _04418_, rst);
  nor _37263_ (_04419_, _04104_, _25680_);
  nand _37264_ (_04420_, _04104_, _26359_);
  nand _37265_ (_04421_, _04420_, _26487_);
  nor _37266_ (_28198_[2], _04421_, _04419_);
  nor _37267_ (_04423_, _04104_, _25194_);
  nand _37268_ (_04424_, _04104_, _25869_);
  nand _37269_ (_04425_, _04424_, _26487_);
  nor _37270_ (_28198_[3], _04425_, _04423_);
  nor _37271_ (_04426_, _04104_, _25028_);
  nand _37272_ (_04427_, _04104_, _26018_);
  nand _37273_ (_04428_, _04427_, _26487_);
  nor _37274_ (_28198_[4], _04428_, _04426_);
  nor _37275_ (_04429_, _04104_, _26096_);
  nor _37276_ (_04430_, _04410_, _26072_);
  nor _37277_ (_04431_, _04430_, _04429_);
  nor _37278_ (_28198_[5], _04431_, rst);
  nor _37279_ (_04434_, _04104_, _25140_);
  nor _37280_ (_04435_, _04410_, _25958_);
  nor _37281_ (_04437_, _04435_, _04434_);
  nor _37282_ (_28198_[6], _04437_, rst);
  nor _37283_ (_04440_, _04111_, _26301_);
  nor _37284_ (_04442_, _04358_, _04110_);
  nor _37285_ (_04443_, _04442_, _04440_);
  nor _37286_ (_28199_[0], _04443_, rst);
  nor _37287_ (_04444_, _04111_, _26461_);
  nor _37288_ (_04445_, _04113_, _25088_);
  nor _37289_ (_04446_, _04445_, _04444_);
  nor _37290_ (_28199_[1], _04446_, rst);
  nor _37291_ (_04447_, _04111_, _26348_);
  nor _37292_ (_04449_, _04113_, _25703_);
  nor _37293_ (_04450_, _04449_, _04447_);
  nor _37294_ (_28199_[2], _04450_, rst);
  nor _37295_ (_04451_, _04113_, _25195_);
  nor _37296_ (_04452_, _04111_, _25866_);
  nor _37297_ (_04453_, _04452_, _04451_);
  nor _37298_ (_28199_[3], _04453_, rst);
  nor _37299_ (_04454_, _04113_, _25029_);
  nor _37300_ (_04455_, _04111_, _26030_);
  nor _37301_ (_04456_, _04455_, _04454_);
  nor _37302_ (_28199_[4], _04456_, rst);
  nor _37303_ (_04457_, _04113_, _26096_);
  nor _37304_ (_04458_, _04111_, _26074_);
  nor _37305_ (_04459_, _04458_, _04457_);
  nor _37306_ (_28199_[5], _04459_, rst);
  nor _37307_ (_04460_, _04113_, _25140_);
  nor _37308_ (_04461_, _04111_, _25947_);
  nor _37309_ (_04462_, _04461_, _04460_);
  nor _37310_ (_28199_[6], _04462_, rst);
  nor _37311_ (_04464_, _04123_, _26289_);
  nor _37312_ (_04465_, _24850_, _26289_);
  nand _37313_ (_04466_, _04465_, _04121_);
  nor _37314_ (_04467_, _04130_, _24850_);
  nand _37315_ (_04468_, _04467_, _24821_);
  nand _37316_ (_04470_, _04468_, _04466_);
  nor _37317_ (_04471_, _04470_, _04464_);
  nor _37318_ (_28200_[0], _04471_, rst);
  nor _37319_ (_04473_, _04127_, _26454_);
  nor _37320_ (_04475_, _25088_, _04130_);
  nor _37321_ (_04476_, _04133_, _26454_);
  nor _37322_ (_04477_, _04476_, _04475_);
  nor _37323_ (_04478_, _04477_, _24850_);
  nor _37324_ (_04479_, _04478_, _04473_);
  nor _37325_ (_28200_[1], _04479_, rst);
  not _37326_ (_04480_, _04467_);
  nor _37327_ (_04482_, _04480_, _25703_);
  nor _37328_ (_04484_, _04467_, _26341_);
  nor _37329_ (_04485_, _04484_, _04482_);
  nor _37330_ (_28200_[2], _04485_, rst);
  nor _37331_ (_04486_, _04127_, _25860_);
  nor _37332_ (_04487_, _25195_, _04130_);
  nor _37333_ (_04488_, _04133_, _25860_);
  nor _37334_ (_04490_, _04488_, _04487_);
  nor _37335_ (_04491_, _04490_, _24850_);
  nor _37336_ (_04492_, _04491_, _04486_);
  nor _37337_ (_28200_[3], _04492_, rst);
  nor _37338_ (_04493_, _04127_, _26024_);
  nor _37339_ (_04494_, _25029_, _04130_);
  nor _37340_ (_04495_, _04133_, _26024_);
  nor _37341_ (_04496_, _04495_, _04494_);
  nor _37342_ (_04497_, _04496_, _24850_);
  nor _37343_ (_04498_, _04497_, _04493_);
  nor _37344_ (_28200_[4], _04498_, rst);
  nor _37345_ (_04499_, _04480_, _26096_);
  nand _37346_ (_04500_, _04125_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor _37347_ (_04502_, _24850_, _26088_);
  nand _37348_ (_04503_, _04502_, _04121_);
  nand _37349_ (_04505_, _04503_, _04500_);
  nor _37350_ (_04508_, _04505_, _04499_);
  nor _37351_ (_28200_[5], _04508_, rst);
  nor _37352_ (_04509_, _04127_, _25940_);
  nor _37353_ (_04510_, _25140_, _04130_);
  nor _37354_ (_04511_, _04133_, _25940_);
  nor _37355_ (_04513_, _04511_, _04510_);
  nor _37356_ (_04514_, _04513_, _24850_);
  nor _37357_ (_04515_, _04514_, _04509_);
  nor _37358_ (_28200_[6], _04515_, rst);
  not _37359_ (_04517_, _04140_);
  nor _37360_ (_04518_, _04358_, _04517_);
  nor _37361_ (_04520_, _04151_, _26293_);
  nor _37362_ (_04521_, _04520_, _04518_);
  nor _37363_ (_28201_[0], _04521_, rst);
  nor _37364_ (_04522_, _04141_, _25088_);
  nor _37365_ (_04523_, _04151_, _26450_);
  nor _37366_ (_04524_, _04523_, _04522_);
  nor _37367_ (_28201_[1], _04524_, rst);
  nor _37368_ (_04525_, _04141_, _25703_);
  nor _37369_ (_04526_, _04151_, _26343_);
  nor _37370_ (_04528_, _04526_, _04525_);
  nor _37371_ (_28201_[2], _04528_, rst);
  nor _37372_ (_04529_, _04141_, _25195_);
  nor _37373_ (_04530_, _04151_, _25871_);
  nor _37374_ (_04531_, _04530_, _04529_);
  nor _37375_ (_28201_[3], _04531_, rst);
  nor _37376_ (_04532_, _04141_, _25029_);
  not _37377_ (_04533_, _04149_);
  nor _37378_ (_04534_, _04533_, _04148_);
  nor _37379_ (_04536_, _04534_, _26032_);
  nor _37380_ (_04537_, _04536_, _04532_);
  nor _37381_ (_28201_[4], _04537_, rst);
  nor _37382_ (_04538_, _04534_, _26085_);
  nor _37383_ (_04539_, _04141_, _26096_);
  nor _37384_ (_04541_, _04539_, _04538_);
  nor _37385_ (_28201_[5], _04541_, rst);
  nor _37386_ (_04542_, _04141_, _25140_);
  nor _37387_ (_04543_, _04151_, _25942_);
  nor _37388_ (_04544_, _04543_, _04542_);
  nor _37389_ (_28201_[6], _04544_, rst);
  nor _37390_ (_04545_, _04156_, _26299_);
  nor _37391_ (_04546_, _04358_, _04155_);
  nor _37392_ (_04547_, _04546_, _04545_);
  nor _37393_ (_28202_[0], _04547_, rst);
  nor _37394_ (_04548_, _04157_, _25088_);
  nor _37395_ (_04549_, _04156_, _26459_);
  nor _37396_ (_04550_, _04549_, _04548_);
  nor _37397_ (_28202_[1], _04550_, rst);
  nor _37398_ (_04552_, _04157_, _25703_);
  nor _37399_ (_04553_, _04156_, _26357_);
  nor _37400_ (_04554_, _04553_, _04552_);
  nor _37401_ (_28202_[2], _04554_, rst);
  nor _37402_ (_04555_, _04157_, _25195_);
  nor _37403_ (_04556_, _04156_, _25855_);
  nor _37404_ (_04557_, _04556_, _04555_);
  nor _37405_ (_28202_[3], _04557_, rst);
  nor _37406_ (_04558_, _04157_, _25029_);
  nor _37407_ (_04559_, _04156_, _26035_);
  nor _37408_ (_04560_, _04559_, _04558_);
  nor _37409_ (_28202_[4], _04560_, rst);
  nor _37410_ (_04562_, _04156_, _26083_);
  nor _37411_ (_04563_, _04157_, _26096_);
  nor _37412_ (_04564_, _04563_, _04562_);
  nor _37413_ (_28202_[5], _04564_, rst);
  nor _37414_ (_04566_, _04157_, _25140_);
  nor _37415_ (_04567_, _04156_, _25956_);
  nor _37416_ (_04569_, _04567_, _04566_);
  nor _37417_ (_28202_[6], _04569_, rst);
  nand _37418_ (_04570_, _03958_, _25203_);
  nand _37419_ (_04571_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nand _37420_ (_26617_, _04571_, _04570_);
  nor _37421_ (_04573_, _24848_, _24820_);
  nor _37422_ (_04575_, _24852_, _26295_);
  nor _37423_ (_04576_, _04575_, _04573_);
  nand _37424_ (_04577_, _24850_, _26295_);
  nand _37425_ (_04579_, _04577_, _26487_);
  nor _37426_ (_28203_[0], _04579_, _04576_);
  nor _37427_ (_04580_, _25088_, _24855_);
  nor _37428_ (_04581_, _24852_, _26456_);
  nor _37429_ (_04583_, _04581_, _04580_);
  nor _37430_ (_28203_[1], _04583_, rst);
  nor _37431_ (_04584_, _24852_, _26346_);
  nor _37432_ (_04585_, _25703_, _24855_);
  nor _37433_ (_04586_, _04585_, _04584_);
  nor _37434_ (_28203_[2], _04586_, rst);
  nor _37435_ (_04587_, _25195_, _24855_);
  nor _37436_ (_04588_, _24852_, _25853_);
  nor _37437_ (_04589_, _04588_, _04587_);
  nor _37438_ (_28203_[3], _04589_, rst);
  nor _37439_ (_04590_, _24852_, _26026_);
  nor _37440_ (_04591_, _25029_, _24855_);
  nor _37441_ (_04592_, _04591_, _04590_);
  nor _37442_ (_28203_[4], _04592_, rst);
  nor _37443_ (_04594_, _24852_, _26090_);
  nor _37444_ (_04596_, _26096_, _24855_);
  nor _37445_ (_04597_, _04596_, _04594_);
  nor _37446_ (_28203_[5], _04597_, rst);
  nor _37447_ (_04598_, _25140_, _24855_);
  nor _37448_ (_04599_, _24852_, _25945_);
  nor _37449_ (_04600_, _04599_, _04598_);
  nor _37450_ (_28203_[6], _04600_, rst);
  nor _37451_ (_04601_, _00114_, _25051_);
  not _37452_ (_04602_, _04601_);
  nand _37453_ (_04603_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nand _37454_ (_04604_, _04601_, _25099_);
  nand _37455_ (_26631_, _04604_, _04603_);
  nand _37456_ (_04606_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  nand _37457_ (_04607_, _24927_, _24796_);
  nand _37458_ (_27085_, _04607_, _04606_);
  nand _37459_ (_04608_, _04251_, _28096_);
  nand _37460_ (_04609_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  nand _37461_ (_27110_, _04609_, _04608_);
  nor _37462_ (_04610_, _00954_, _25051_);
  not _37463_ (_04611_, _04610_);
  nand _37464_ (_04613_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  nand _37465_ (_04614_, _04610_, _25150_);
  nand _37466_ (_27128_, _04614_, _04613_);
  nand _37467_ (_04615_, _03958_, _24830_);
  nand _37468_ (_04616_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  nand _37469_ (_27156_, _04616_, _04615_);
  nand _37470_ (_04617_, _00632_, _25150_);
  nand _37471_ (_04618_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  nand _37472_ (_27162_, _04618_, _04617_);
  nand _37473_ (_04620_, _01398_, _25150_);
  nand _37474_ (_04621_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  nand _37475_ (_27165_, _04621_, _04620_);
  nand _37476_ (_04622_, _03876_, _28096_);
  nand _37477_ (_04623_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  nand _37478_ (_27170_, _04623_, _04622_);
  nor _37479_ (_04624_, _00114_, _25059_);
  nand _37480_ (_04625_, _04624_, _24789_);
  not _37481_ (_04626_, _04624_);
  nand _37482_ (_04627_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  nand _37483_ (_27257_, _04627_, _04625_);
  nand _37484_ (_04628_, _03377_, _03373_);
  nor _37485_ (_04629_, _04628_, _03369_);
  nor _37486_ (_04630_, _04629_, _00551_);
  nor _37487_ (_04631_, _04630_, _00615_);
  nor _37488_ (_04632_, _25627_, _24845_);
  nand _37489_ (_04633_, _04632_, _26244_);
  nand _37490_ (_04634_, _04633_, _04631_);
  nand _37491_ (_04635_, _04634_, _00622_);
  nor _37492_ (_04637_, _04633_, _24716_);
  nor _37493_ (_04638_, _04637_, _04635_);
  nor _37494_ (_04639_, _00622_, _25088_);
  nor _37495_ (_04640_, _04639_, _04638_);
  nor _37496_ (_27260_, _04640_, rst);
  nand _37497_ (_04642_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor _37498_ (_04643_, _04642_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  nand _37499_ (_04644_, _04643_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor _37500_ (_28377_, _04644_, rst);
  not _37501_ (_04646_, _04643_);
  nand _37502_ (_04647_, _04646_, _26487_);
  not _37503_ (_04648_, _04642_);
  nand _37504_ (_04650_, _04648_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  not _37505_ (_04652_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand _37506_ (_04653_, _04642_, _04652_);
  nand _37507_ (_04654_, _04653_, _04650_);
  nor _37508_ (_28378_[3], _04654_, _04647_);
  nand _37509_ (_04655_, _26124_, _25993_);
  nor _37510_ (_04656_, _26059_, _25843_);
  not _37511_ (_04657_, _04656_);
  nor _37512_ (_04659_, _04657_, _25919_);
  not _37513_ (_04660_, _04659_);
  nor _37514_ (_04662_, _04660_, _04655_);
  not _37515_ (_04664_, _04662_);
  nand _37516_ (_04666_, _02685_, _26234_);
  not _37517_ (_04667_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _37518_ (_04668_, _26250_, _04667_);
  not _37519_ (_04669_, _04668_);
  nor _37520_ (_04670_, _00146_, _04667_);
  not _37521_ (_04671_, _04670_);
  nand _37522_ (_04672_, _04671_, _00381_);
  nor _37523_ (_04673_, _26247_, _26236_);
  nand _37524_ (_04675_, _04673_, _04672_);
  nand _37525_ (_04676_, _04675_, _04669_);
  nor _37526_ (_04678_, _04676_, _26226_);
  nand _37527_ (_04679_, _04678_, _04666_);
  nor _37528_ (_04680_, _02727_, _26225_);
  not _37529_ (_04681_, _04680_);
  nand _37530_ (_04682_, _04681_, _04679_);
  nand _37531_ (_04683_, _02761_, _26234_);
  not _37532_ (_04684_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _37533_ (_04685_, _26250_, _04684_);
  not _37534_ (_04686_, _04685_);
  nand _37535_ (_04687_, _03356_, _24716_);
  nor _37536_ (_04689_, _03356_, _04684_);
  not _37537_ (_04690_, _04689_);
  nand _37538_ (_04692_, _04690_, _04687_);
  nand _37539_ (_04693_, _04692_, _04673_);
  nand _37540_ (_04694_, _04693_, _04686_);
  nor _37541_ (_04695_, _04694_, _26226_);
  nand _37542_ (_04696_, _04695_, _04683_);
  nand _37543_ (_04697_, _02802_, _26226_);
  nand _37544_ (_04698_, _04697_, _04696_);
  nand _37545_ (_04700_, _04698_, _04682_);
  nor _37546_ (_04701_, _02229_, _26233_);
  not _37547_ (_04702_, _04678_);
  nor _37548_ (_04703_, _04702_, _04701_);
  nor _37549_ (_04704_, _04680_, _04703_);
  nor _37550_ (_04706_, _02307_, _26233_);
  not _37551_ (_04707_, _04695_);
  nor _37552_ (_04708_, _04707_, _04706_);
  not _37553_ (_04710_, _04697_);
  nor _37554_ (_04711_, _04710_, _04708_);
  nand _37555_ (_04712_, _04711_, _04704_);
  nand _37556_ (_04713_, _04712_, _04700_);
  not _37557_ (_04714_, _02369_);
  nor _37558_ (_04715_, _04714_, _02330_);
  nand _37559_ (_04716_, _04715_, _02341_);
  nor _37560_ (_04717_, _04716_, _02337_);
  nor _37561_ (_04718_, _04717_, _26233_);
  nor _37562_ (_04719_, _26250_, _24541_);
  not _37563_ (_04720_, _04719_);
  nand _37564_ (_04721_, _01665_, _24716_);
  nor _37565_ (_04722_, _01665_, _24541_);
  not _37566_ (_04723_, _04722_);
  nand _37567_ (_04724_, _04723_, _04721_);
  nand _37568_ (_04725_, _04724_, _04673_);
  nand _37569_ (_04726_, _04725_, _04720_);
  nor _37570_ (_04727_, _04726_, _26226_);
  not _37571_ (_04728_, _04727_);
  nor _37572_ (_04729_, _04728_, _04718_);
  nor _37573_ (_04730_, _02861_, _26225_);
  nor _37574_ (_04731_, _04730_, _04729_);
  nor _37575_ (_04732_, _27460_, _26233_);
  nor _37576_ (_04733_, _26250_, _24124_);
  not _37577_ (_04734_, _04733_);
  nor _37578_ (_04736_, _26135_, _24124_);
  not _37579_ (_04737_, _04736_);
  nand _37580_ (_04738_, _04737_, _00225_);
  nand _37581_ (_04739_, _04738_, _04673_);
  nand _37582_ (_04740_, _04739_, _04734_);
  nor _37583_ (_04742_, _04740_, _26226_);
  not _37584_ (_04744_, _04742_);
  nor _37585_ (_04745_, _04744_, _04732_);
  nor _37586_ (_04746_, _27564_, _26225_);
  nor _37587_ (_04747_, _04746_, _04745_);
  nor _37588_ (_04749_, _04747_, _04731_);
  nand _37589_ (_04750_, _02373_, _26234_);
  nand _37590_ (_04751_, _04727_, _04750_);
  not _37591_ (_04752_, _04730_);
  nand _37592_ (_04753_, _04752_, _04751_);
  nand _37593_ (_04754_, _02415_, _26234_);
  nand _37594_ (_04755_, _04742_, _04754_);
  not _37595_ (_04756_, _27503_);
  nor _37596_ (_04757_, _04756_, _27500_);
  nor _37597_ (_04759_, _04757_, _24089_);
  nor _37598_ (_04760_, _27561_, _04759_);
  nand _37599_ (_04761_, _04760_, _26226_);
  nand _37600_ (_04762_, _04761_, _04755_);
  nor _37601_ (_04763_, _04762_, _04753_);
  nor _37602_ (_04764_, _04763_, _04749_);
  nand _37603_ (_04766_, _04764_, _04713_);
  nor _37604_ (_04767_, _04711_, _04704_);
  nor _37605_ (_04768_, _04698_, _04682_);
  nor _37606_ (_04769_, _04768_, _04767_);
  nand _37607_ (_04770_, _04762_, _04753_);
  nand _37608_ (_04771_, _04747_, _04731_);
  nand _37609_ (_04772_, _04771_, _04770_);
  nand _37610_ (_04773_, _04772_, _04769_);
  nand _37611_ (_04774_, _04773_, _04766_);
  nor _37612_ (_04775_, _02448_, _26233_);
  nor _37613_ (_04776_, _26250_, _24404_);
  not _37614_ (_04777_, _04776_);
  nor _37615_ (_04778_, _25722_, _24404_);
  not _37616_ (_04779_, _04778_);
  nand _37617_ (_04780_, _04779_, _03655_);
  nand _37618_ (_04781_, _04780_, _04673_);
  nand _37619_ (_04782_, _04781_, _04777_);
  nor _37620_ (_04783_, _04782_, _26226_);
  not _37621_ (_04784_, _04783_);
  nor _37622_ (_04785_, _04784_, _04775_);
  nand _37623_ (_04786_, _02478_, _26226_);
  not _37624_ (_04787_, _04786_);
  nor _37625_ (_04788_, _04787_, _04785_);
  nor _37626_ (_04789_, _02041_, _26233_);
  not _37627_ (_04790_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _37628_ (_04791_, _26250_, _04790_);
  not _37629_ (_04792_, _04791_);
  nor _37630_ (_04793_, _24840_, _04790_);
  not _37631_ (_04794_, _04793_);
  nand _37632_ (_04795_, _04794_, _01280_);
  nand _37633_ (_04796_, _04795_, _04673_);
  nand _37634_ (_04797_, _04796_, _04792_);
  nor _37635_ (_04799_, _04797_, _26226_);
  not _37636_ (_04800_, _04799_);
  nor _37637_ (_04801_, _04800_, _04789_);
  nand _37638_ (_04802_, _02540_, _26226_);
  not _37639_ (_04803_, _04802_);
  nor _37640_ (_04804_, _04803_, _04801_);
  nand _37641_ (_04805_, _04804_, _04788_);
  nand _37642_ (_04806_, _01974_, _26234_);
  nand _37643_ (_04807_, _04783_, _04806_);
  nand _37644_ (_04808_, _04786_, _04807_);
  nand _37645_ (_04809_, _02509_, _26234_);
  nand _37646_ (_04810_, _04799_, _04809_);
  nand _37647_ (_04811_, _04802_, _04810_);
  nand _37648_ (_04812_, _04811_, _04808_);
  nand _37649_ (_04813_, _04812_, _04805_);
  nand _37650_ (_04814_, _02096_, _26234_);
  nor _37651_ (_04815_, _26250_, _24302_);
  not _37652_ (_04817_, _04815_);
  nor _37653_ (_04818_, _00275_, _24302_);
  not _37654_ (_04819_, _04818_);
  nand _37655_ (_04820_, _04819_, _03603_);
  nand _37656_ (_04821_, _04820_, _04673_);
  nand _37657_ (_04822_, _04821_, _04817_);
  nor _37658_ (_04823_, _04822_, _26226_);
  nand _37659_ (_04824_, _04823_, _04814_);
  nor _37660_ (_04826_, _02599_, _26225_);
  not _37661_ (_04827_, _04826_);
  nand _37662_ (_04828_, _04827_, _04824_);
  nor _37663_ (_04829_, _02160_, _26233_);
  nor _37664_ (_04830_, _26250_, _24271_);
  not _37665_ (_04831_, _04830_);
  nor _37666_ (_04833_, _00444_, _24271_);
  not _37667_ (_04834_, _04833_);
  nand _37668_ (_04835_, _04834_, _00489_);
  nand _37669_ (_04836_, _04835_, _04673_);
  nand _37670_ (_04837_, _04836_, _04831_);
  nor _37671_ (_04839_, _04837_, _26226_);
  not _37672_ (_04841_, _04839_);
  nor _37673_ (_04842_, _04841_, _04829_);
  nand _37674_ (_04844_, _02652_, _26226_);
  not _37675_ (_04845_, _04844_);
  nor _37676_ (_04847_, _04845_, _04842_);
  nor _37677_ (_04848_, _04847_, _04828_);
  nor _37678_ (_04849_, _02564_, _26233_);
  not _37679_ (_04850_, _04823_);
  nor _37680_ (_04851_, _04850_, _04849_);
  nor _37681_ (_04852_, _04826_, _04851_);
  nand _37682_ (_04853_, _02620_, _26234_);
  nand _37683_ (_04854_, _04839_, _04853_);
  nand _37684_ (_04855_, _04844_, _04854_);
  nor _37685_ (_04856_, _04855_, _04852_);
  nor _37686_ (_04858_, _04856_, _04848_);
  nand _37687_ (_04860_, _04858_, _04813_);
  nor _37688_ (_04861_, _04811_, _04808_);
  nor _37689_ (_04862_, _04804_, _04788_);
  nor _37690_ (_04864_, _04862_, _04861_);
  nand _37691_ (_04865_, _04855_, _04852_);
  nand _37692_ (_04867_, _04847_, _04828_);
  nand _37693_ (_04868_, _04867_, _04865_);
  nand _37694_ (_04870_, _04868_, _04864_);
  nand _37695_ (_04871_, _04870_, _04860_);
  nand _37696_ (_04872_, _04871_, _04774_);
  nor _37697_ (_04873_, _04772_, _04769_);
  nor _37698_ (_04874_, _04764_, _04713_);
  nor _37699_ (_04875_, _04874_, _04873_);
  nor _37700_ (_04876_, _04868_, _04864_);
  nor _37701_ (_04877_, _04858_, _04813_);
  nor _37702_ (_04878_, _04877_, _04876_);
  nand _37703_ (_04879_, _04878_, _04875_);
  nand _37704_ (_04880_, _04879_, _04872_);
  nor _37705_ (_04881_, _04880_, _26400_);
  nor _37706_ (_04882_, _26472_, _26338_);
  nand _37707_ (_04883_, _26400_, _25720_);
  nand _37708_ (_04884_, _04883_, _04882_);
  nor _37709_ (_04885_, _04884_, _04881_);
  nor _37710_ (_04886_, _26472_, _26407_);
  nand _37711_ (_04887_, _04886_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor _37712_ (_04888_, _26473_, _26407_);
  nand _37713_ (_04889_, _04888_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand _37714_ (_04891_, _04889_, _04887_);
  nand _37715_ (_04892_, _04891_, _26400_);
  nor _37716_ (_04893_, _26473_, _26338_);
  not _37717_ (_04894_, _04893_);
  nor _37718_ (_04895_, _26403_, _02078_);
  not _37719_ (_04897_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _37720_ (_04898_, _26400_, _04897_);
  nor _37721_ (_04899_, _04898_, _04895_);
  nor _37722_ (_04900_, _04899_, _04894_);
  not _37723_ (_04901_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  not _37724_ (_04902_, _04886_);
  nor _37725_ (_04903_, _04902_, _04901_);
  not _37726_ (_04904_, _04888_);
  nor _37727_ (_04905_, _04904_, _25738_);
  nor _37728_ (_04906_, _04905_, _04903_);
  nor _37729_ (_04907_, _04906_, _26400_);
  nor _37730_ (_04908_, _04907_, _04900_);
  nand _37731_ (_04909_, _04908_, _04892_);
  nor _37732_ (_04910_, _04909_, _04885_);
  nor _37733_ (_04911_, _04910_, _04664_);
  nand _37734_ (_04912_, _04659_, _04655_);
  nor _37735_ (_04913_, _26058_, _25843_);
  not _37736_ (_04914_, _04913_);
  nor _37737_ (_04915_, _04914_, _04655_);
  not _37738_ (_04916_, _04915_);
  nor _37739_ (_04917_, _04916_, _25916_);
  nor _37740_ (_04919_, _26124_, _25993_);
  not _37741_ (_04920_, _04919_);
  nor _37742_ (_04922_, _04920_, _04914_);
  not _37743_ (_04923_, _04922_);
  nor _37744_ (_04924_, _04923_, _25919_);
  nor _37745_ (_04926_, _04924_, _04917_);
  nand _37746_ (_04927_, _04926_, _04912_);
  nor _37747_ (_04928_, _25993_, _25843_);
  nand _37748_ (_04929_, _04928_, _25919_);
  nand _37749_ (_04930_, _04929_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _37750_ (_04931_, _04930_, _04662_);
  nor _37751_ (_04932_, _26124_, _25991_);
  not _37752_ (_04933_, _04932_);
  nor _37753_ (_04934_, _04933_, _04914_);
  not _37754_ (_04936_, _04934_);
  nor _37755_ (_04937_, _04936_, _25919_);
  nand _37756_ (_04939_, _26124_, _25991_);
  nor _37757_ (_04940_, _04939_, _04914_);
  nand _37758_ (_04941_, _04940_, _25916_);
  not _37759_ (_04942_, _04941_);
  nor _37760_ (_04944_, _04942_, _04937_);
  nand _37761_ (_04945_, _04944_, _04931_);
  nor _37762_ (_04947_, _04945_, _04927_);
  nand _37763_ (_04948_, _26481_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not _37764_ (_04949_, _25393_);
  nor _37765_ (_04950_, _26202_, _04949_);
  nor _37766_ (_04952_, _04950_, _25604_);
  not _37767_ (_04953_, _01064_);
  nor _37768_ (_04954_, _04949_, _25298_);
  nor _37769_ (_04955_, _04954_, _04953_);
  not _37770_ (_04957_, _04955_);
  nor _37771_ (_04958_, _25392_, _25235_);
  nor _37772_ (_04959_, _04958_, _25408_);
  nor _37773_ (_04960_, _25583_, _25554_);
  nand _37774_ (_04961_, _04960_, _04959_);
  nor _37775_ (_04962_, _04961_, _04957_);
  nand _37776_ (_04964_, _04962_, _04952_);
  nor _37777_ (_04965_, _01049_, _25473_);
  nor _37778_ (_04967_, _04965_, _25491_);
  not _37779_ (_04968_, _04967_);
  nor _37780_ (_04969_, _25556_, _25424_);
  nand _37781_ (_04971_, _04969_, _25533_);
  nor _37782_ (_04972_, _04971_, _04968_);
  nand _37783_ (_04973_, _04972_, _25581_);
  nor _37784_ (_04974_, _04973_, _04964_);
  nor _37785_ (_04976_, _04974_, _25530_);
  nor _37786_ (_04977_, _04976_, p3_in[7]);
  not _37787_ (_04978_, _04976_);
  nor _37788_ (_04979_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor _37789_ (_04980_, _04979_, _04977_);
  nand _37790_ (_04982_, _04980_, _26400_);
  nor _37791_ (_04984_, _04976_, p3_in[3]);
  nor _37792_ (_04985_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor _37793_ (_04986_, _04985_, _04984_);
  nand _37794_ (_04988_, _04986_, _26403_);
  nand _37795_ (_04989_, _04988_, _04982_);
  nand _37796_ (_04990_, _04989_, _04888_);
  nor _37797_ (_04991_, _04976_, p3_in[4]);
  nor _37798_ (_04992_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor _37799_ (_04994_, _04992_, _04991_);
  nand _37800_ (_04995_, _04994_, _26400_);
  nor _37801_ (_04996_, _04976_, p3_in[0]);
  nor _37802_ (_04998_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _37803_ (_04999_, _04998_, _04996_);
  nand _37804_ (_05000_, _04999_, _26403_);
  nand _37805_ (_05001_, _05000_, _04995_);
  nand _37806_ (_05002_, _05001_, _04882_);
  nand _37807_ (_05003_, _05002_, _04990_);
  nor _37808_ (_05004_, _04976_, p3_in[5]);
  nor _37809_ (_05005_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor _37810_ (_05006_, _05005_, _05004_);
  nand _37811_ (_05007_, _05006_, _26400_);
  nor _37812_ (_05008_, _04976_, p3_in[1]);
  nor _37813_ (_05009_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor _37814_ (_05010_, _05009_, _05008_);
  nand _37815_ (_05011_, _05010_, _26403_);
  nand _37816_ (_05012_, _05011_, _05007_);
  nand _37817_ (_05013_, _05012_, _04886_);
  nor _37818_ (_05014_, _04976_, p3_in[6]);
  nor _37819_ (_05015_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _37820_ (_05017_, _05015_, _05014_);
  nand _37821_ (_05019_, _05017_, _26400_);
  nor _37822_ (_05020_, _04976_, p3_in[2]);
  nor _37823_ (_05021_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor _37824_ (_05022_, _05021_, _05020_);
  nand _37825_ (_05023_, _05022_, _26403_);
  nand _37826_ (_05025_, _05023_, _05019_);
  nand _37827_ (_05026_, _05025_, _04893_);
  nand _37828_ (_05027_, _05026_, _05013_);
  nor _37829_ (_05029_, _05027_, _05003_);
  nor _37830_ (_05030_, _05029_, _04660_);
  nand _37831_ (_05031_, _05030_, _04919_);
  nor _37832_ (_05032_, _26403_, _24541_);
  nor _37833_ (_05034_, _26400_, _24302_);
  nor _37834_ (_05035_, _05034_, _05032_);
  nor _37835_ (_05036_, _05035_, _04894_);
  not _37836_ (_05037_, _04882_);
  nor _37837_ (_05038_, _26403_, _04667_);
  nor _37838_ (_05039_, _26400_, _24404_);
  nor _37839_ (_05041_, _05039_, _05038_);
  nor _37840_ (_05043_, _05041_, _05037_);
  nor _37841_ (_05044_, _05043_, _05036_);
  nor _37842_ (_05046_, _26403_, _24124_);
  nor _37843_ (_05047_, _26400_, _24271_);
  nor _37844_ (_05048_, _05047_, _05046_);
  nor _37845_ (_05049_, _05048_, _04904_);
  nor _37846_ (_05050_, _26403_, _04684_);
  nor _37847_ (_05051_, _26400_, _04790_);
  nor _37848_ (_05052_, _05051_, _05050_);
  nor _37849_ (_05053_, _05052_, _04902_);
  nor _37850_ (_05055_, _05053_, _05049_);
  nand _37851_ (_05056_, _05055_, _05044_);
  nand _37852_ (_05058_, _05056_, _04937_);
  nand _37853_ (_05059_, _05058_, _05031_);
  not _37854_ (_05060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _37855_ (_05061_, _26403_, _05060_);
  nor _37856_ (_05062_, _26400_, _00163_);
  nor _37857_ (_05063_, _05062_, _05061_);
  nor _37858_ (_05064_, _05063_, _04894_);
  nor _37859_ (_05065_, _26403_, _00383_);
  nor _37860_ (_05066_, _26400_, _00154_);
  nor _37861_ (_05067_, _05066_, _05065_);
  nor _37862_ (_05069_, _05067_, _05037_);
  nor _37863_ (_05070_, _05069_, _05064_);
  nor _37864_ (_05071_, _26403_, _00215_);
  not _37865_ (_05072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _37866_ (_05073_, _26400_, _05072_);
  nor _37867_ (_05074_, _05073_, _05071_);
  nor _37868_ (_05075_, _05074_, _04904_);
  not _37869_ (_05076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _37870_ (_05077_, _26403_, _05076_);
  nor _37871_ (_05079_, _26400_, _01200_);
  nor _37872_ (_05080_, _05079_, _05077_);
  nor _37873_ (_05081_, _05080_, _04902_);
  nor _37874_ (_05082_, _05081_, _05075_);
  nand _37875_ (_05083_, _05082_, _05070_);
  nand _37876_ (_05084_, _05083_, _04917_);
  not _37877_ (_05085_, _04939_);
  nor _37878_ (_05087_, _04976_, p1_in[7]);
  nor _37879_ (_05088_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor _37880_ (_05089_, _05088_, _05087_);
  nand _37881_ (_05090_, _05089_, _26400_);
  nor _37882_ (_05091_, _04976_, p1_in[3]);
  nor _37883_ (_05092_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor _37884_ (_05093_, _05092_, _05091_);
  nand _37885_ (_05094_, _05093_, _26403_);
  nand _37886_ (_05095_, _05094_, _05090_);
  nand _37887_ (_05097_, _05095_, _04888_);
  nor _37888_ (_05098_, _04976_, p1_in[6]);
  nor _37889_ (_05100_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _37890_ (_05101_, _05100_, _05098_);
  nand _37891_ (_05102_, _05101_, _26400_);
  nor _37892_ (_05103_, _04976_, p1_in[2]);
  nor _37893_ (_05104_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor _37894_ (_05106_, _05104_, _05103_);
  nand _37895_ (_05108_, _05106_, _26403_);
  nand _37896_ (_05109_, _05108_, _05102_);
  nand _37897_ (_05111_, _05109_, _04893_);
  nand _37898_ (_05112_, _05111_, _05097_);
  nor _37899_ (_05113_, _04976_, p1_in[4]);
  nor _37900_ (_05114_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor _37901_ (_05115_, _05114_, _05113_);
  nand _37902_ (_05116_, _05115_, _26400_);
  nor _37903_ (_05117_, _04976_, p1_in[0]);
  nor _37904_ (_05118_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _37905_ (_05119_, _05118_, _05117_);
  nand _37906_ (_05120_, _05119_, _26403_);
  nand _37907_ (_05121_, _05120_, _05116_);
  nand _37908_ (_05122_, _05121_, _04882_);
  nor _37909_ (_05123_, _04976_, p1_in[5]);
  nor _37910_ (_05124_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor _37911_ (_05125_, _05124_, _05123_);
  nand _37912_ (_05126_, _05125_, _26400_);
  nor _37913_ (_05127_, _04976_, p1_in[1]);
  nor _37914_ (_05128_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor _37915_ (_05129_, _05128_, _05127_);
  nand _37916_ (_05130_, _05129_, _26403_);
  nand _37917_ (_05131_, _05130_, _05126_);
  nand _37918_ (_05132_, _05131_, _04886_);
  nand _37919_ (_05133_, _05132_, _05122_);
  nor _37920_ (_05134_, _05133_, _05112_);
  nor _37921_ (_05135_, _05134_, _04660_);
  nand _37922_ (_05136_, _05135_, _05085_);
  nand _37923_ (_05137_, _05136_, _05084_);
  nor _37924_ (_05138_, _05137_, _05059_);
  nand _37925_ (_05139_, _05138_, _04948_);
  nor _37926_ (_05140_, _05139_, _04947_);
  nand _37927_ (_05141_, _04656_, _25919_);
  nor _37928_ (_05143_, _05141_, _04920_);
  nor _37929_ (_05145_, _26403_, _03392_);
  nor _37930_ (_05146_, _26400_, _00561_);
  nor _37931_ (_05148_, _05146_, _05145_);
  nor _37932_ (_05149_, _05148_, _04894_);
  nor _37933_ (_05151_, _26403_, _00422_);
  nor _37934_ (_05152_, _26400_, _00473_);
  nor _37935_ (_05153_, _05152_, _05151_);
  nor _37936_ (_05155_, _05153_, _05037_);
  nor _37937_ (_05156_, _05155_, _05149_);
  nor _37938_ (_05157_, _26403_, _00577_);
  nor _37939_ (_05158_, _26400_, _00555_);
  nor _37940_ (_05159_, _05158_, _05157_);
  nor _37941_ (_05160_, _05159_, _04902_);
  not _37942_ (_05161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor _37943_ (_05162_, _26403_, _05161_);
  nor _37944_ (_05164_, _26400_, _00447_);
  nor _37945_ (_05166_, _05164_, _05162_);
  nor _37946_ (_05167_, _05166_, _04904_);
  nor _37947_ (_05169_, _05167_, _05160_);
  nand _37948_ (_05170_, _05169_, _05156_);
  nand _37949_ (_05171_, _05170_, _05143_);
  nor _37950_ (_05172_, _04976_, p2_in[5]);
  nor _37951_ (_05173_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor _37952_ (_05174_, _05173_, _05172_);
  nand _37953_ (_05175_, _05174_, _26400_);
  nor _37954_ (_05176_, _04976_, p2_in[1]);
  nor _37955_ (_05177_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor _37956_ (_05178_, _05177_, _05176_);
  nand _37957_ (_05179_, _05178_, _26403_);
  nand _37958_ (_05180_, _05179_, _05175_);
  nand _37959_ (_05181_, _05180_, _26473_);
  nor _37960_ (_05183_, _04976_, p2_in[7]);
  nor _37961_ (_05184_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor _37962_ (_05185_, _05184_, _05183_);
  nand _37963_ (_05186_, _05185_, _26400_);
  nor _37964_ (_05187_, _04976_, p2_in[3]);
  nor _37965_ (_05188_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor _37966_ (_05189_, _05188_, _05187_);
  nand _37967_ (_05190_, _05189_, _26403_);
  nand _37968_ (_05191_, _05190_, _05186_);
  nand _37969_ (_05192_, _05191_, _26472_);
  nand _37970_ (_05193_, _05192_, _05181_);
  nand _37971_ (_05194_, _05193_, _26338_);
  nor _37972_ (_05195_, _04976_, p2_in[4]);
  nor _37973_ (_05196_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _37974_ (_05197_, _05196_, _05195_);
  nand _37975_ (_05198_, _05197_, _26400_);
  nor _37976_ (_05199_, _04976_, p2_in[0]);
  nor _37977_ (_05201_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _37978_ (_05202_, _05201_, _05199_);
  nand _37979_ (_05203_, _05202_, _26403_);
  nand _37980_ (_05205_, _05203_, _05198_);
  nand _37981_ (_05206_, _05205_, _26473_);
  nor _37982_ (_05207_, _04976_, p2_in[6]);
  nor _37983_ (_05208_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor _37984_ (_05209_, _05208_, _05207_);
  nand _37985_ (_05210_, _05209_, _26400_);
  nor _37986_ (_05211_, _04976_, p2_in[2]);
  nor _37987_ (_05212_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor _37988_ (_05213_, _05212_, _05211_);
  nand _37989_ (_05214_, _05213_, _26403_);
  nand _37990_ (_05215_, _05214_, _05210_);
  nand _37991_ (_05216_, _05215_, _26472_);
  nand _37992_ (_05217_, _05216_, _05206_);
  nand _37993_ (_05218_, _05217_, _26407_);
  nand _37994_ (_05219_, _05218_, _05194_);
  nand _37995_ (_05220_, _05219_, _04924_);
  nand _37996_ (_05221_, _05220_, _05171_);
  nor _37997_ (_05222_, _04914_, _25916_);
  nand _37998_ (_05223_, _26400_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand _37999_ (_05225_, _26403_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nand _38000_ (_05226_, _05225_, _05223_);
  nand _38001_ (_05227_, _05226_, _04886_);
  nand _38002_ (_05228_, _26400_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  nand _38003_ (_05229_, _26403_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nand _38004_ (_05230_, _05229_, _05228_);
  nand _38005_ (_05231_, _05230_, _04893_);
  nand _38006_ (_05232_, _26400_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _38007_ (_05233_, _26403_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _38008_ (_05234_, _05233_, _05232_);
  nand _38009_ (_05235_, _05234_, _04882_);
  nand _38010_ (_05236_, _05235_, _05231_);
  nor _38011_ (_05237_, _26403_, _00543_);
  not _38012_ (_05238_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor _38013_ (_05239_, _26400_, _05238_);
  nor _38014_ (_05240_, _05239_, _05237_);
  nor _38015_ (_05241_, _05240_, _04904_);
  nor _38016_ (_05242_, _05241_, _05236_);
  nand _38017_ (_05243_, _05242_, _05227_);
  nand _38018_ (_05244_, _05243_, _04919_);
  nor _38019_ (_05245_, _26403_, _01603_);
  nor _38020_ (_05246_, _26400_, _03496_);
  nor _38021_ (_05247_, _05246_, _05245_);
  nor _38022_ (_05248_, _05247_, _04894_);
  nor _38023_ (_05249_, _26403_, _01582_);
  nor _38024_ (_05250_, _26400_, _00615_);
  nor _38025_ (_05252_, _05250_, _05249_);
  nor _38026_ (_05253_, _05252_, _05037_);
  nor _38027_ (_05255_, _05253_, _05248_);
  nand _38028_ (_05257_, _04886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nor _38029_ (_05258_, _04904_, _00562_);
  nor _38030_ (_05259_, _05258_, _26400_);
  nand _38031_ (_05260_, _05259_, _05257_);
  nand _38032_ (_05261_, _04886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nor _38033_ (_05263_, _04904_, _03974_);
  nor _38034_ (_05264_, _05263_, _26403_);
  nand _38035_ (_05266_, _05264_, _05261_);
  nand _38036_ (_05267_, _05266_, _05260_);
  nand _38037_ (_05269_, _05267_, _05255_);
  nand _38038_ (_05270_, _05269_, _05085_);
  nand _38039_ (_05271_, _05270_, _05244_);
  nand _38040_ (_05273_, _05271_, _05222_);
  nand _38041_ (_05274_, _04932_, _04659_);
  not _38042_ (_05275_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor _38043_ (_05276_, _26403_, _05275_);
  not _38044_ (_05277_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _38045_ (_05278_, _26400_, _05277_);
  nor _38046_ (_05279_, _05278_, _05276_);
  nor _38047_ (_05281_, _05279_, _04902_);
  not _38048_ (_05282_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor _38049_ (_05284_, _26403_, _05282_);
  not _38050_ (_05285_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor _38051_ (_05286_, _26400_, _05285_);
  nor _38052_ (_05287_, _05286_, _05284_);
  nor _38053_ (_05288_, _05287_, _04894_);
  not _38054_ (_05290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor _38055_ (_05291_, _26403_, _05290_);
  not _38056_ (_05292_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor _38057_ (_05293_, _26400_, _05292_);
  nor _38058_ (_05295_, _05293_, _05291_);
  nor _38059_ (_05296_, _05295_, _05037_);
  nor _38060_ (_05297_, _05296_, _05288_);
  nand _38061_ (_05298_, _26400_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _38062_ (_05299_, _26403_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _38063_ (_05300_, _05299_, _05298_);
  nand _38064_ (_05301_, _05300_, _04888_);
  nand _38065_ (_05302_, _05301_, _05297_);
  nor _38066_ (_05304_, _05302_, _05281_);
  nor _38067_ (_05305_, _05304_, _05274_);
  nor _38068_ (_05306_, _05141_, _04939_);
  nand _38069_ (_05307_, _26400_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nand _38070_ (_05308_, _26403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _38071_ (_05309_, _05308_, _05307_);
  nand _38072_ (_05311_, _05309_, _04886_);
  nand _38073_ (_05313_, _26400_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _38074_ (_05314_, _26403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _38075_ (_05316_, _05314_, _05313_);
  nand _38076_ (_05318_, _05316_, _04882_);
  nand _38077_ (_05319_, _26400_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _38078_ (_05320_, _26403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand _38079_ (_05322_, _05320_, _05319_);
  nand _38080_ (_05323_, _05322_, _04893_);
  nand _38081_ (_05325_, _05323_, _05318_);
  not _38082_ (_05327_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _38083_ (_05328_, _26403_, _05327_);
  nor _38084_ (_05329_, _26400_, _01294_);
  nor _38085_ (_05331_, _05329_, _05328_);
  nor _38086_ (_05333_, _05331_, _04904_);
  nor _38087_ (_05334_, _05333_, _05325_);
  nand _38088_ (_05336_, _05334_, _05311_);
  nand _38089_ (_05337_, _05336_, _05306_);
  nor _38090_ (_05338_, _04976_, p0_in[5]);
  nor _38091_ (_05339_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor _38092_ (_05340_, _05339_, _05338_);
  nand _38093_ (_05341_, _05340_, _26400_);
  nor _38094_ (_05342_, _04976_, p0_in[1]);
  nor _38095_ (_05343_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor _38096_ (_05344_, _05343_, _05342_);
  nand _38097_ (_05345_, _05344_, _26403_);
  nand _38098_ (_05346_, _05345_, _05341_);
  nand _38099_ (_05347_, _05346_, _26473_);
  nor _38100_ (_05348_, _04976_, p0_in[7]);
  nor _38101_ (_05349_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor _38102_ (_05350_, _05349_, _05348_);
  nand _38103_ (_05351_, _05350_, _26400_);
  nor _38104_ (_05352_, _04976_, p0_in[3]);
  nor _38105_ (_05354_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor _38106_ (_05355_, _05354_, _05352_);
  nand _38107_ (_05356_, _05355_, _26403_);
  nand _38108_ (_05357_, _05356_, _05351_);
  nand _38109_ (_05359_, _05357_, _26472_);
  nand _38110_ (_05361_, _05359_, _05347_);
  nand _38111_ (_05362_, _05361_, _26338_);
  nor _38112_ (_05364_, _04976_, p0_in[4]);
  nor _38113_ (_05365_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor _38114_ (_05367_, _05365_, _05364_);
  nand _38115_ (_05368_, _05367_, _26400_);
  nor _38116_ (_05370_, _04976_, p0_in[0]);
  nor _38117_ (_05371_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _38118_ (_05372_, _05371_, _05370_);
  nand _38119_ (_05374_, _05372_, _26403_);
  nand _38120_ (_05376_, _05374_, _05368_);
  nand _38121_ (_05378_, _05376_, _26473_);
  nor _38122_ (_05379_, _04976_, p0_in[6]);
  nor _38123_ (_05380_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _38124_ (_05382_, _05380_, _05379_);
  nand _38125_ (_05383_, _05382_, _26400_);
  nor _38126_ (_05384_, _04976_, p0_in[2]);
  nor _38127_ (_05386_, _04978_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor _38128_ (_05388_, _05386_, _05384_);
  nand _38129_ (_05390_, _05388_, _26403_);
  nand _38130_ (_05392_, _05390_, _05383_);
  nand _38131_ (_05393_, _05392_, _26472_);
  nand _38132_ (_05394_, _05393_, _05378_);
  nand _38133_ (_05396_, _05394_, _26407_);
  nand _38134_ (_05398_, _05396_, _05362_);
  nand _38135_ (_05399_, _05398_, _04942_);
  nand _38136_ (_05401_, _05399_, _05337_);
  nor _38137_ (_05403_, _05401_, _05305_);
  nand _38138_ (_05404_, _05403_, _05273_);
  nor _38139_ (_05405_, _05404_, _05221_);
  nand _38140_ (_05406_, _05405_, _05140_);
  nor _38141_ (_05407_, _05406_, _04911_);
  not _38142_ (_05408_, _26137_);
  not _38143_ (_05410_, _26229_);
  not _38144_ (_05411_, _04937_);
  nor _38145_ (_05413_, _05411_, _05410_);
  nor _38146_ (_05414_, _05413_, _05408_);
  not _38147_ (_05415_, _04948_);
  nand _38148_ (_05416_, _05415_, _24717_);
  nand _38149_ (_05417_, _05416_, _05414_);
  nor _38150_ (_05418_, _05417_, _05407_);
  nor _38151_ (_05419_, _26403_, _26096_);
  nor _38152_ (_05421_, _26400_, _25088_);
  nor _38153_ (_05423_, _05421_, _05419_);
  nor _38154_ (_05425_, _05423_, _04902_);
  nor _38155_ (_05426_, _26403_, _25029_);
  nor _38156_ (_05427_, _26400_, _24820_);
  nor _38157_ (_05428_, _05427_, _05426_);
  nor _38158_ (_05430_, _05428_, _05037_);
  nor _38159_ (_05431_, _26403_, _25140_);
  nor _38160_ (_05433_, _26400_, _25703_);
  nor _38161_ (_05435_, _05433_, _05431_);
  nor _38162_ (_05436_, _05435_, _04894_);
  nor _38163_ (_05437_, _05436_, _05430_);
  nand _38164_ (_05438_, _26400_, _24782_);
  nand _38165_ (_05439_, _26403_, _25194_);
  nand _38166_ (_05440_, _05439_, _05438_);
  nand _38167_ (_05441_, _05440_, _04888_);
  nand _38168_ (_05442_, _05441_, _05437_);
  nor _38169_ (_05443_, _05442_, _05425_);
  nor _38170_ (_05444_, _05443_, _05414_);
  nor _38171_ (_05445_, _05444_, _05418_);
  nor _38172_ (_28379_, _05445_, rst);
  nor _38173_ (_05446_, _26400_, _25919_);
  not _38174_ (_05447_, _05446_);
  nor _38175_ (_05448_, _05447_, _05037_);
  not _38176_ (_05450_, _05448_);
  nor _38177_ (_05452_, _05450_, _04936_);
  not _38178_ (_05453_, _05452_);
  nor _38179_ (_05454_, _05453_, _05410_);
  nor _38180_ (_05455_, _04904_, _26403_);
  nor _38181_ (_05456_, _05455_, _01275_);
  nand _38182_ (_05457_, _05456_, _26132_);
  not _38183_ (_05459_, _05457_);
  nor _38184_ (_05460_, _05459_, _05454_);
  nand _38185_ (_05461_, _05460_, _26483_);
  nor _38186_ (_05462_, _05453_, _26225_);
  nor _38187_ (_05463_, _05450_, _04657_);
  not _38188_ (_05464_, _05463_);
  nor _38189_ (_05465_, _05464_, _04655_);
  not _38190_ (_05466_, _05465_);
  nor _38191_ (_05467_, _05466_, _26252_);
  nor _38192_ (_05468_, _05467_, _05462_);
  nor _38193_ (_05469_, _26228_, _26223_);
  nor _38194_ (_05470_, _05447_, _04904_);
  nand _38195_ (_05472_, _05470_, _04940_);
  not _38196_ (_05473_, _05472_);
  nand _38197_ (_05475_, _05473_, _05469_);
  nand _38198_ (_05476_, _05475_, _05468_);
  nand _38199_ (_05478_, _05476_, _23870_);
  not _38200_ (_05479_, _05478_);
  nor _38201_ (_05480_, _05479_, _05461_);
  not _38202_ (_05481_, _05469_);
  nand _38203_ (_05482_, _04940_, _04893_);
  nor _38204_ (_05484_, _05482_, _05447_);
  not _38205_ (_05486_, _05484_);
  nor _38206_ (_05487_, _05486_, _05481_);
  not _38207_ (_05488_, _05487_);
  nand _38208_ (_05489_, _05488_, _26487_);
  nor _38209_ (_28380_, _05489_, _05480_);
  nor _38210_ (_05492_, _26400_, _25916_);
  not _38211_ (_05493_, _05492_);
  nor _38212_ (_05495_, _05493_, _05037_);
  not _38213_ (_05497_, _05495_);
  nor _38214_ (_05498_, _05497_, _04916_);
  nand _38215_ (_05499_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _38216_ (_05500_, _26403_, _25916_);
  not _38217_ (_05501_, _05500_);
  nor _38218_ (_05502_, _05501_, _05037_);
  not _38219_ (_05503_, _05502_);
  nor _38220_ (_05505_, _05503_, _04916_);
  nand _38221_ (_05506_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _38222_ (_05507_, _05506_, _05499_);
  nor _38223_ (_05508_, _05501_, _04902_);
  not _38224_ (_05509_, _05508_);
  nor _38225_ (_05511_, _05509_, _04916_);
  nand _38226_ (_05512_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor _38227_ (_05513_, _05493_, _04894_);
  not _38228_ (_05515_, _05513_);
  nor _38229_ (_05516_, _05515_, _04916_);
  nand _38230_ (_05517_, _05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand _38231_ (_05518_, _05517_, _05512_);
  nor _38232_ (_05520_, _05518_, _05507_);
  nand _38233_ (_05521_, _05495_, _04940_);
  not _38234_ (_05522_, _05521_);
  nand _38235_ (_05523_, _05522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor _38236_ (_05524_, _05493_, _04904_);
  nand _38237_ (_05526_, _05524_, _04915_);
  not _38238_ (_05528_, _05526_);
  nand _38239_ (_05530_, _05528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _38240_ (_05531_, _05530_, _05523_);
  nand _38241_ (_05533_, _05495_, _04922_);
  not _38242_ (_05534_, _05533_);
  nand _38243_ (_05535_, _05534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not _38244_ (_05536_, _05455_);
  nor _38245_ (_05537_, _05536_, _25919_);
  nor _38246_ (_05538_, _04920_, _04657_);
  nand _38247_ (_05539_, _05538_, _05537_);
  not _38248_ (_05540_, _05539_);
  nand _38249_ (_05541_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand _38250_ (_05542_, _05541_, _05535_);
  nor _38251_ (_05544_, _05542_, _05531_);
  nand _38252_ (_05546_, _05544_, _05520_);
  not _38253_ (_05547_, _04940_);
  nor _38254_ (_05548_, _05493_, _04902_);
  not _38255_ (_05550_, _05548_);
  nor _38256_ (_05551_, _05550_, _05547_);
  nand _38257_ (_05552_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nand _38258_ (_05553_, _05524_, _04940_);
  not _38259_ (_05554_, _05553_);
  nand _38260_ (_05555_, _05554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand _38261_ (_05556_, _05555_, _05552_);
  nor _38262_ (_05557_, _05509_, _05547_);
  nand _38263_ (_05558_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _38264_ (_05559_, _05515_, _05547_);
  nand _38265_ (_05560_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand _38266_ (_05561_, _05560_, _05558_);
  nor _38267_ (_05562_, _05561_, _05556_);
  nor _38268_ (_05563_, _04939_, _04657_);
  not _38269_ (_05564_, _05563_);
  nor _38270_ (_05565_, _05564_, _05550_);
  nand _38271_ (_05566_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nor _38272_ (_05567_, _05497_, _05564_);
  nand _38273_ (_05568_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand _38274_ (_05570_, _05568_, _05566_);
  nor _38275_ (_05571_, _05503_, _05547_);
  nand _38276_ (_05572_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _38277_ (_05574_, _05537_, _04940_);
  not _38278_ (_05575_, _05574_);
  nand _38279_ (_05577_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _38280_ (_05578_, _05577_, _05572_);
  nor _38281_ (_05579_, _05578_, _05570_);
  nand _38282_ (_05581_, _05579_, _05562_);
  nor _38283_ (_05582_, _05581_, _05546_);
  nand _38284_ (_05584_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand _38285_ (_05585_, _05473_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand _38286_ (_05586_, _05585_, _05584_);
  nand _38287_ (_05587_, _05463_, _04932_);
  not _38288_ (_05588_, _05587_);
  nand _38289_ (_05589_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor _38290_ (_05590_, _05447_, _04902_);
  nand _38291_ (_05592_, _05590_, _04940_);
  not _38292_ (_05593_, _05592_);
  nand _38293_ (_05595_, _05593_, _25927_);
  nand _38294_ (_05597_, _05595_, _05589_);
  nor _38295_ (_05599_, _05597_, _05586_);
  nor _38296_ (_05600_, _05564_, _05450_);
  nand _38297_ (_05601_, _05600_, _05089_);
  nor _38298_ (_05602_, _05450_, _05547_);
  nand _38299_ (_05604_, _05602_, _05350_);
  nand _38300_ (_05605_, _05604_, _05601_);
  nor _38301_ (_05606_, _05450_, _04923_);
  nand _38302_ (_05607_, _05606_, _05185_);
  not _38303_ (_05609_, _05538_);
  nor _38304_ (_05611_, _05609_, _05450_);
  nand _38305_ (_05612_, _05611_, _04980_);
  nand _38306_ (_05614_, _05612_, _05607_);
  nor _38307_ (_05616_, _05614_, _05605_);
  nand _38308_ (_05617_, _05616_, _05599_);
  nand _38309_ (_05618_, _05465_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand _38310_ (_05619_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand _38311_ (_05620_, _05619_, _05618_);
  nor _38312_ (_05621_, _05620_, _05617_);
  nand _38313_ (_05622_, _05621_, _05582_);
  nand _38314_ (_05624_, _05622_, _05480_);
  nor _38315_ (_05625_, _05505_, _05498_);
  nor _38316_ (_05627_, _05516_, _05511_);
  nand _38317_ (_05628_, _05627_, _05625_);
  not _38318_ (_05629_, _05628_);
  nor _38319_ (_05630_, _05528_, _05522_);
  not _38320_ (_05632_, _05630_);
  nand _38321_ (_05633_, _05539_, _05533_);
  nor _38322_ (_05634_, _05633_, _05632_);
  nand _38323_ (_05636_, _05634_, _05629_);
  nor _38324_ (_05637_, _05554_, _05551_);
  nor _38325_ (_05638_, _05559_, _05557_);
  nand _38326_ (_05639_, _05638_, _05637_);
  not _38327_ (_05640_, _05639_);
  not _38328_ (_05641_, _05571_);
  nand _38329_ (_05642_, _05574_, _05641_);
  nor _38330_ (_05643_, _05567_, _05565_);
  not _38331_ (_05644_, _05643_);
  nor _38332_ (_05645_, _05644_, _05642_);
  nand _38333_ (_05646_, _05645_, _05640_);
  nor _38334_ (_05648_, _05646_, _05636_);
  nand _38335_ (_05649_, _05448_, _04928_);
  nor _38336_ (_05650_, _05484_, _05473_);
  not _38337_ (_05651_, _05650_);
  nand _38338_ (_05652_, _05592_, _05587_);
  nor _38339_ (_05653_, _05652_, _05651_);
  nand _38340_ (_05654_, _05653_, _05649_);
  nor _38341_ (_05655_, _05465_, _05452_);
  not _38342_ (_05656_, _05655_);
  nor _38343_ (_05657_, _05656_, _05654_);
  nand _38344_ (_05658_, _05657_, _05648_);
  nand _38345_ (_05659_, _05658_, _05480_);
  nand _38346_ (_05660_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _38347_ (_05661_, _05660_, _05624_);
  nor _38348_ (_05662_, _05661_, _05487_);
  nand _38349_ (_05663_, _05487_, _27460_);
  nand _38350_ (_05664_, _05663_, _26487_);
  nor _38351_ (_28381_[7], _05664_, _05662_);
  nand _38352_ (_05665_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nand _38353_ (_05666_, _04322_, _25039_);
  nand _38354_ (_27337_, _05666_, _05665_);
  nand _38355_ (_05667_, _00955_, _24789_);
  nand _38356_ (_05668_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  nand _38357_ (_27341_, _05668_, _05667_);
  nand _38358_ (_05669_, _03834_, _25099_);
  nand _38359_ (_05670_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nand _38360_ (_27343_, _05670_, _05669_);
  nand _38361_ (_05671_, _01398_, _24927_);
  nand _38362_ (_05672_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  nand _38363_ (_27364_, _05672_, _05671_);
  nand _38364_ (_05675_, _01402_, _25039_);
  nand _38365_ (_05676_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  nand _38366_ (_27374_, _05676_, _05675_);
  nand _38367_ (_05678_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nand _38368_ (_05679_, _04322_, _24830_);
  nand _38369_ (_27419_, _05679_, _05678_);
  nand _38370_ (_05680_, _04312_, _25099_);
  nand _38371_ (_05682_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  nand _38372_ (_27422_, _05682_, _05680_);
  nand _38373_ (_05683_, _01398_, _25039_);
  nand _38374_ (_05684_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  nand _38375_ (_27428_, _05684_, _05683_);
  nor _38376_ (_05685_, _03546_, _28073_);
  not _38377_ (_05686_, _05685_);
  nand _38378_ (_05688_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  nand _38379_ (_05690_, _05685_, _24789_);
  nand _38380_ (_27435_, _05690_, _05688_);
  nand _38381_ (_05691_, _03834_, _24830_);
  nand _38382_ (_05693_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nand _38383_ (_27440_, _05693_, _05691_);
  nand _38384_ (_05695_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nand _38385_ (_05697_, _04322_, _25099_);
  nand _38386_ (_27490_, _05697_, _05695_);
  nand _38387_ (_05698_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nand _38388_ (_05699_, _05685_, _28096_);
  nand _38389_ (_27501_, _05699_, _05698_);
  nand _38390_ (_05700_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  nand _38391_ (_05701_, _05685_, _25203_);
  nand _38392_ (_27513_, _05701_, _05700_);
  nand _38393_ (_05702_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  nand _38394_ (_05704_, _05685_, _25099_);
  nand _38395_ (_27518_, _05704_, _05702_);
  nand _38396_ (_05705_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  nand _38397_ (_05706_, _05685_, _24927_);
  nand _38398_ (_27559_, _05706_, _05705_);
  nand _38399_ (_05708_, _03958_, _25099_);
  nand _38400_ (_05709_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nand _38401_ (_27562_, _05709_, _05708_);
  nand _38402_ (_05711_, _28105_, _28096_);
  nand _38403_ (_05712_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  nand _38404_ (_27585_, _05712_, _05711_);
  nand _38405_ (_05715_, _01371_, _24927_);
  nand _38406_ (_05716_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  nand _38407_ (_27588_, _05716_, _05715_);
  nand _38408_ (_05718_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  nand _38409_ (_05719_, _05685_, _25039_);
  nand _38410_ (_27593_, _05719_, _05718_);
  nand _38411_ (_05721_, _01278_, _26135_);
  nand _38412_ (_05722_, _05721_, _05327_);
  nand _38413_ (_05724_, _05722_, _01293_);
  nor _38414_ (_05725_, _05721_, _24716_);
  nor _38415_ (_05726_, _05725_, _05724_);
  nor _38416_ (_05727_, _01293_, _25625_);
  nor _38417_ (_05729_, _05727_, _05726_);
  nor _38418_ (_27621_, _05729_, rst);
  not _38419_ (_05730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _38420_ (_05731_, _03635_, _05730_);
  nand _38421_ (_05733_, _05731_, _26487_);
  nor _38422_ (_05734_, _03635_, _24782_);
  nor _38423_ (_27623_, _05734_, _05733_);
  nor _38424_ (_05735_, _03546_, _00122_);
  not _38425_ (_05736_, _05735_);
  nand _38426_ (_05737_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nand _38427_ (_05738_, _05735_, _25150_);
  nand _38428_ (_27627_, _05738_, _05737_);
  nor _38429_ (_05739_, _28057_, _24795_);
  nand _38430_ (_05740_, _05739_, _24830_);
  not _38431_ (_05741_, _05739_);
  nand _38432_ (_05742_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nand _38433_ (_27630_, _05742_, _05740_);
  nor _38434_ (_05743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _38435_ (_05744_, _05743_, _01241_);
  nand _38436_ (_05745_, _05744_, _01435_);
  nand _38437_ (_05746_, _01450_, _01524_);
  nand _38438_ (_05747_, _01479_, _01462_);
  nand _38439_ (_05748_, _05747_, _05746_);
  nand _38440_ (_05749_, _05748_, _05745_);
  nand _38441_ (_05750_, _01456_, _01524_);
  nand _38442_ (_05751_, _05750_, _05749_);
  nand _38443_ (_27655_, _05751_, _01415_);
  nand _38444_ (_05753_, _01415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _38445_ (_27658_, _05753_, _03761_);
  not _38446_ (_05754_, _03756_);
  nor _38447_ (_05756_, _05754_, _01443_);
  nor _38448_ (_05757_, _05756_, _03737_);
  nor _38449_ (_27661_, _05757_, rst);
  nor _38450_ (_05759_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nand _38451_ (_05761_, _05759_, _01444_);
  nor _38452_ (_05762_, _01479_, _05761_);
  nor _38453_ (_05763_, _05762_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _38454_ (_05764_, _05762_, _03739_);
  nand _38455_ (_05766_, _05764_, _26487_);
  nor _38456_ (_27665_, _05766_, _05763_);
  nor _38457_ (_05767_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _01426_);
  nor _38458_ (_05769_, _05767_, _01432_);
  nand _38459_ (_05770_, _05769_, _01477_);
  nand _38460_ (_05771_, _05770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor _38461_ (_05772_, _05770_, _03739_);
  nor _38462_ (_05774_, _05772_, rst);
  nand _38463_ (_27668_, _05774_, _05771_);
  not _38464_ (_05775_, _03973_);
  nor _38465_ (_05777_, _05775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor _38466_ (_05779_, _05327_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor _38467_ (_05780_, _00259_, _00383_);
  nor _38468_ (_05781_, _05780_, _05779_);
  not _38469_ (_05783_, _05781_);
  nor _38470_ (_05784_, _05783_, _05777_);
  not _38471_ (_05785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _38472_ (_05786_, _05730_, _05785_);
  nand _38473_ (_05788_, _05786_, _26487_);
  nor _38474_ (_27690_, _05788_, _05784_);
  not _38475_ (_05790_, _01346_);
  not _38476_ (_05791_, _01251_);
  not _38477_ (_05792_, _01339_);
  nor _38478_ (_05794_, _05792_, _01349_);
  nand _38479_ (_05795_, _05794_, _05791_);
  nor _38480_ (_05797_, _05795_, _05790_);
  nor _38481_ (_05798_, _05791_, _01272_);
  nor _38482_ (_05799_, _05798_, _05797_);
  nor _38483_ (_05800_, _05799_, _01248_);
  nand _38484_ (_05801_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _38485_ (_05802_, _05801_, _01247_);
  nor _38486_ (_05803_, _05802_, _05800_);
  nor _38487_ (_05805_, _05803_, _01245_);
  nor _38488_ (_05806_, _01351_, _01358_);
  nor _38489_ (_05808_, _05806_, _05805_);
  nor _38490_ (_27693_, _05808_, _01377_);
  not _38491_ (_05810_, _01246_);
  nand _38492_ (_05812_, _05797_, _05810_);
  nand _38493_ (_05813_, _05812_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _38494_ (_05815_, _05813_, _05806_);
  nor _38495_ (_05816_, _05815_, _01261_);
  nor _38496_ (_27697_, _05816_, rst);
  nor _38497_ (_05817_, _05784_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _38498_ (_05818_, _05817_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _38499_ (_05819_, _05817_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _38500_ (_05820_, _05819_, _26487_);
  nor _38501_ (_27702_, _05820_, _05818_);
  nand _38502_ (_05821_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  nand _38503_ (_05822_, _05735_, _24789_);
  nand _38504_ (_27706_, _05822_, _05821_);
  nand _38505_ (_05824_, _01259_, _25628_);
  nor _38506_ (_05825_, _05824_, _24920_);
  not _38507_ (_05826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand _38508_ (_05828_, _05824_, _05826_);
  nand _38509_ (_05829_, _05828_, _26487_);
  nor _38510_ (_27718_, _05829_, _05825_);
  nand _38511_ (_05830_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  nand _38512_ (_05831_, _05735_, _28096_);
  nand _38513_ (_27810_, _05831_, _05830_);
  nand _38514_ (_05832_, _01371_, _25039_);
  nand _38515_ (_05834_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  nand _38516_ (_27821_, _05834_, _05832_);
  nand _38517_ (_05836_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nand _38518_ (_05837_, _05735_, _25099_);
  nand _38519_ (_27842_, _05837_, _05836_);
  nand _38520_ (_05838_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nand _38521_ (_05840_, _05735_, _25039_);
  nand _38522_ (_27906_, _05840_, _05838_);
  nand _38523_ (_05841_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nand _38524_ (_05842_, _05735_, _25203_);
  nand _38525_ (_27913_, _05842_, _05841_);
  nand _38526_ (_05844_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  nand _38527_ (_05845_, _04610_, _28096_);
  nand _38528_ (_27985_, _05845_, _05844_);
  nor _38529_ (_05847_, _03546_, _25047_);
  not _38530_ (_05848_, _05847_);
  nand _38531_ (_05849_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  nand _38532_ (_05850_, _05847_, _25150_);
  nand _38533_ (_28018_, _05850_, _05849_);
  nand _38534_ (_05851_, _28096_, _25152_);
  nand _38535_ (_05852_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  nand _38536_ (_28058_, _05852_, _05851_);
  nand _38537_ (_05853_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  nand _38538_ (_05854_, _05847_, _24789_);
  nand _38539_ (_28067_, _05854_, _05853_);
  nand _38540_ (_05855_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nand _38541_ (_05856_, _01388_, _25039_);
  nand _38542_ (_28079_, _05856_, _05855_);
  nand _38543_ (_05857_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  nand _38544_ (_05858_, _05847_, _28096_);
  nand _38545_ (_28090_, _05858_, _05857_);
  nand _38546_ (_05859_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nand _38547_ (_05861_, _05847_, _25039_);
  nand _38548_ (_28112_, _05861_, _05859_);
  nand _38549_ (_05862_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  nand _38550_ (_05863_, _05847_, _25203_);
  nand _38551_ (_00003_, _05863_, _05862_);
  nor _38552_ (_05864_, _24882_, _24073_);
  not _38553_ (_05865_, _05864_);
  nand _38554_ (_05867_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  nand _38555_ (_05868_, _05864_, _25039_);
  nand _38556_ (_00020_, _05868_, _05867_);
  nor _38557_ (_28378_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  nor _38558_ (_05870_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nand _38559_ (_05871_, _04642_, _26487_);
  nor _38560_ (_28378_[1], _05871_, _05870_);
  nand _38561_ (_05872_, _04642_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  nand _38562_ (_05873_, _05872_, _04646_);
  nand _38563_ (_05874_, _05873_, _04644_);
  nor _38564_ (_28378_[2], _05874_, rst);
  not _38565_ (_05875_, _05480_);
  not _38566_ (_05876_, _04880_);
  nor _38567_ (_05877_, _05466_, _05876_);
  not _38568_ (_05879_, _05372_);
  not _38569_ (_05880_, _05602_);
  nor _38570_ (_05883_, _05880_, _05879_);
  nand _38571_ (_05884_, _05600_, _05119_);
  nand _38572_ (_05885_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nand _38573_ (_05886_, _05885_, _05884_);
  nor _38574_ (_05887_, _05886_, _05883_);
  nand _38575_ (_05889_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _38576_ (_05891_, _26277_);
  nand _38577_ (_05892_, _04940_, _04886_);
  nor _38578_ (_05894_, _05892_, _05447_);
  nand _38579_ (_05895_, _05894_, _05891_);
  nand _38580_ (_05896_, _05895_, _05889_);
  nand _38581_ (_05898_, _05606_, _05202_);
  nor _38582_ (_05899_, _05464_, _04920_);
  nand _38583_ (_05900_, _05899_, _04999_);
  nand _38584_ (_05901_, _05900_, _05898_);
  nor _38585_ (_05902_, _05901_, _05896_);
  nand _38586_ (_05903_, _05902_, _05887_);
  not _38587_ (_05904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not _38588_ (_05906_, _05516_);
  nor _38589_ (_05907_, _05906_, _05904_);
  nor _38590_ (_05908_, _05536_, _04941_);
  nand _38591_ (_05909_, _05908_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand _38592_ (_05910_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand _38593_ (_05911_, _05910_, _05909_);
  nor _38594_ (_05912_, _05911_, _05907_);
  nand _38595_ (_05914_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _38596_ (_05915_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _38597_ (_05917_, _05915_, _05914_);
  nand _38598_ (_05919_, _04940_, _04888_);
  nor _38599_ (_05920_, _05493_, _05919_);
  nand _38600_ (_05921_, _05920_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _38601_ (_05922_, _05493_, _05482_);
  nand _38602_ (_05924_, _05922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _38603_ (_05925_, _05924_, _05921_);
  nor _38604_ (_05926_, _05925_, _05917_);
  nand _38605_ (_05927_, _05926_, _05912_);
  nor _38606_ (_05928_, _05927_, _05903_);
  nand _38607_ (_05929_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  not _38608_ (_05931_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nor _38609_ (_05932_, _05919_, _05447_);
  not _38610_ (_05933_, _05932_);
  nor _38611_ (_05934_, _05933_, _05931_);
  nand _38612_ (_05935_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _38613_ (_05937_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _38614_ (_05939_, _05937_, _05935_);
  nor _38615_ (_05941_, _05939_, _05934_);
  nand _38616_ (_05942_, _05941_, _05929_);
  nor _38617_ (_05943_, _05533_, _00550_);
  nor _38618_ (_05944_, _05521_, _00615_);
  not _38619_ (_05946_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _38620_ (_05947_, _05526_, _05946_);
  nor _38621_ (_05949_, _05947_, _05944_);
  nand _38622_ (_05950_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _38623_ (_05952_, _05950_, _05949_);
  nor _38624_ (_05953_, _05952_, _05943_);
  not _38625_ (_05955_, _05511_);
  nor _38626_ (_05956_, _05955_, _00183_);
  nand _38627_ (_05958_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _38628_ (_05959_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _38629_ (_05961_, _05959_, _05958_);
  nor _38630_ (_05962_, _05961_, _05956_);
  nand _38631_ (_05963_, _05962_, _05953_);
  nor _38632_ (_05964_, _05963_, _05942_);
  nand _38633_ (_05965_, _05964_, _05928_);
  nor _38634_ (_05966_, _05965_, _05877_);
  nor _38635_ (_05967_, _05966_, _05875_);
  nand _38636_ (_05968_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _38637_ (_05969_, _05968_, _05488_);
  nor _38638_ (_05970_, _05969_, _05967_);
  nand _38639_ (_05971_, _05487_, _02448_);
  nand _38640_ (_05972_, _05971_, _26487_);
  nor _38641_ (_28381_[0], _05972_, _05970_);
  nand _38642_ (_05973_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nand _38643_ (_05974_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _38644_ (_05975_, _05974_, _05973_);
  nand _38645_ (_05977_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _38646_ (_05979_, _05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand _38647_ (_05980_, _05979_, _05977_);
  nor _38648_ (_05981_, _05980_, _05975_);
  nand _38649_ (_05982_, _05528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nand _38650_ (_05984_, _05522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand _38651_ (_05985_, _05984_, _05982_);
  nand _38652_ (_05986_, _05534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nand _38653_ (_05987_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nand _38654_ (_05988_, _05987_, _05986_);
  nor _38655_ (_05989_, _05988_, _05985_);
  nand _38656_ (_05990_, _05989_, _05981_);
  nand _38657_ (_05991_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand _38658_ (_05992_, _05554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _38659_ (_05994_, _05992_, _05991_);
  nand _38660_ (_05996_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _38661_ (_05997_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nand _38662_ (_05998_, _05997_, _05996_);
  nor _38663_ (_05999_, _05998_, _05994_);
  nand _38664_ (_06000_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  nand _38665_ (_06001_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _38666_ (_06002_, _06001_, _06000_);
  nand _38667_ (_06003_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _38668_ (_06005_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  nand _38669_ (_06006_, _06005_, _06003_);
  nor _38670_ (_06007_, _06006_, _06002_);
  nand _38671_ (_06009_, _06007_, _05999_);
  nor _38672_ (_06010_, _06009_, _05990_);
  nand _38673_ (_06011_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand _38674_ (_06012_, _05932_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand _38675_ (_06013_, _06012_, _06011_);
  nand _38676_ (_06015_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not _38677_ (_06016_, _26440_);
  nand _38678_ (_06017_, _05894_, _06016_);
  nand _38679_ (_06018_, _06017_, _06015_);
  nor _38680_ (_06020_, _06018_, _06013_);
  nand _38681_ (_06022_, _05602_, _05344_);
  nand _38682_ (_06024_, _05600_, _05129_);
  nand _38683_ (_06025_, _06024_, _06022_);
  nand _38684_ (_06026_, _05606_, _05178_);
  nand _38685_ (_06027_, _05611_, _05010_);
  nand _38686_ (_06029_, _06027_, _06026_);
  nor _38687_ (_06030_, _06029_, _06025_);
  nand _38688_ (_06031_, _06030_, _06020_);
  nand _38689_ (_06032_, _05465_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand _38690_ (_06033_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand _38691_ (_06035_, _06033_, _06032_);
  nor _38692_ (_06036_, _06035_, _06031_);
  nand _38693_ (_06037_, _06036_, _06010_);
  nand _38694_ (_06038_, _06037_, _05480_);
  nand _38695_ (_06039_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _38696_ (_06040_, _06039_, _06038_);
  nor _38697_ (_06042_, _06040_, _05487_);
  nand _38698_ (_06044_, _05487_, _02041_);
  nand _38699_ (_06045_, _06044_, _26487_);
  nor _38700_ (_28381_[1], _06045_, _06042_);
  nand _38701_ (_06047_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand _38702_ (_06048_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  nand _38703_ (_06049_, _06048_, _06047_);
  nand _38704_ (_06050_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _38705_ (_06051_, _05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand _38706_ (_06052_, _06051_, _06050_);
  nor _38707_ (_06053_, _06052_, _06049_);
  nand _38708_ (_06054_, _05522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _38709_ (_06055_, _05528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nand _38710_ (_06056_, _06055_, _06054_);
  nand _38711_ (_06057_, _05534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nand _38712_ (_06058_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand _38713_ (_06059_, _06058_, _06057_);
  nor _38714_ (_06060_, _06059_, _06056_);
  nand _38715_ (_06061_, _06060_, _06053_);
  nand _38716_ (_06062_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nand _38717_ (_06064_, _05554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand _38718_ (_06065_, _06064_, _06062_);
  nand _38719_ (_06067_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _38720_ (_06068_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand _38721_ (_06070_, _06068_, _06067_);
  nor _38722_ (_06072_, _06070_, _06065_);
  nand _38723_ (_06074_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  nand _38724_ (_06076_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand _38725_ (_06077_, _06076_, _06074_);
  nand _38726_ (_06078_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _38727_ (_06080_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  nand _38728_ (_06082_, _06080_, _06078_);
  nor _38729_ (_06084_, _06082_, _06077_);
  nand _38730_ (_06086_, _06084_, _06072_);
  nor _38731_ (_06087_, _06086_, _06061_);
  nand _38732_ (_06088_, _05465_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand _38733_ (_06089_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand _38734_ (_06090_, _06089_, _06088_);
  nand _38735_ (_06092_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _38736_ (_06093_, _26396_);
  nand _38737_ (_06095_, _05894_, _06093_);
  nand _38738_ (_06096_, _06095_, _06092_);
  nand _38739_ (_06098_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand _38740_ (_06100_, _05473_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand _38741_ (_06101_, _06100_, _06098_);
  nor _38742_ (_06102_, _06101_, _06096_);
  nand _38743_ (_06103_, _05600_, _05106_);
  nand _38744_ (_06104_, _05602_, _05388_);
  nand _38745_ (_06106_, _06104_, _06103_);
  nand _38746_ (_06107_, _05606_, _05213_);
  nand _38747_ (_06108_, _05611_, _05022_);
  nand _38748_ (_06109_, _06108_, _06107_);
  nor _38749_ (_06110_, _06109_, _06106_);
  nand _38750_ (_06111_, _06110_, _06102_);
  nor _38751_ (_06113_, _06111_, _06090_);
  nand _38752_ (_06114_, _06113_, _06087_);
  nand _38753_ (_06115_, _06114_, _05480_);
  nand _38754_ (_06116_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _38755_ (_06117_, _06116_, _06115_);
  nor _38756_ (_06119_, _06117_, _05487_);
  nand _38757_ (_06121_, _05487_, _02564_);
  nand _38758_ (_06122_, _06121_, _26487_);
  nor _38759_ (_28381_[2], _06122_, _06119_);
  nand _38760_ (_06124_, _05461_, _24261_);
  nand _38761_ (_06125_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nand _38762_ (_06126_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nand _38763_ (_06127_, _06126_, _06125_);
  nand _38764_ (_06128_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _38765_ (_06130_, _05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand _38766_ (_06131_, _06130_, _06128_);
  nor _38767_ (_06132_, _06131_, _06127_);
  nand _38768_ (_06133_, _05528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nand _38769_ (_06135_, _05522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand _38770_ (_06136_, _06135_, _06133_);
  nand _38771_ (_06138_, _05534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nand _38772_ (_06139_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand _38773_ (_06141_, _06139_, _06138_);
  nor _38774_ (_06142_, _06141_, _06136_);
  nand _38775_ (_06143_, _06142_, _06132_);
  nand _38776_ (_06144_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  nand _38777_ (_06145_, _05554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand _38778_ (_06146_, _06145_, _06144_);
  nand _38779_ (_06147_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _38780_ (_06148_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand _38781_ (_06149_, _06148_, _06147_);
  nor _38782_ (_06150_, _06149_, _06146_);
  nand _38783_ (_06152_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand _38784_ (_06153_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  nand _38785_ (_06154_, _06153_, _06152_);
  nand _38786_ (_06155_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _38787_ (_06157_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  nand _38788_ (_06159_, _06157_, _06155_);
  nor _38789_ (_06160_, _06159_, _06154_);
  nand _38790_ (_06161_, _06160_, _06150_);
  nor _38791_ (_06162_, _06161_, _06143_);
  nand _38792_ (_06163_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not _38793_ (_06164_, _25892_);
  nand _38794_ (_06166_, _05894_, _06164_);
  nand _38795_ (_06167_, _06166_, _06163_);
  nand _38796_ (_06169_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand _38797_ (_06171_, _05473_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nand _38798_ (_06172_, _06171_, _06169_);
  nor _38799_ (_06173_, _06172_, _06167_);
  nand _38800_ (_06175_, _05602_, _05355_);
  nand _38801_ (_06176_, _05600_, _05093_);
  nand _38802_ (_06177_, _06176_, _06175_);
  nand _38803_ (_06178_, _05606_, _05189_);
  nand _38804_ (_06179_, _05611_, _04986_);
  nand _38805_ (_06180_, _06179_, _06178_);
  nor _38806_ (_06182_, _06180_, _06177_);
  nand _38807_ (_06183_, _06182_, _06173_);
  nand _38808_ (_06184_, _05465_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand _38809_ (_06185_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand _38810_ (_06186_, _06185_, _06184_);
  nor _38811_ (_06187_, _06186_, _06183_);
  nand _38812_ (_06188_, _06187_, _06162_);
  nand _38813_ (_06189_, _06188_, _05478_);
  nand _38814_ (_06190_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _38815_ (_06191_, _06190_, _06189_);
  nand _38816_ (_06192_, _06191_, _06124_);
  nor _38817_ (_06193_, _06192_, _05487_);
  nor _38818_ (_06194_, _05488_, _02160_);
  nor _38819_ (_06195_, _06194_, _06193_);
  nor _38820_ (_28381_[3], _06195_, rst);
  nand _38821_ (_06196_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _38822_ (_06197_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _38823_ (_06199_, _06197_, _06196_);
  nand _38824_ (_06201_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand _38825_ (_06202_, _05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _38826_ (_06203_, _06202_, _06201_);
  nor _38827_ (_06204_, _06203_, _06199_);
  nand _38828_ (_06205_, _05528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand _38829_ (_06207_, _05522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand _38830_ (_06208_, _06207_, _06205_);
  nand _38831_ (_06209_, _05534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _38832_ (_06210_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nand _38833_ (_06212_, _06210_, _06209_);
  nor _38834_ (_06213_, _06212_, _06208_);
  nand _38835_ (_06215_, _06213_, _06204_);
  nand _38836_ (_06216_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand _38837_ (_06217_, _05554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _38838_ (_06218_, _06217_, _06216_);
  nand _38839_ (_06220_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _38840_ (_06221_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand _38841_ (_06222_, _06221_, _06220_);
  nor _38842_ (_06223_, _06222_, _06218_);
  nand _38843_ (_06224_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _38844_ (_06225_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand _38845_ (_06226_, _06225_, _06224_);
  nand _38846_ (_06228_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _38847_ (_06229_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  nand _38848_ (_06230_, _06229_, _06228_);
  nor _38849_ (_06231_, _06230_, _06226_);
  nand _38850_ (_06233_, _06231_, _06223_);
  nor _38851_ (_06234_, _06233_, _06215_);
  nand _38852_ (_06235_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand _38853_ (_06236_, _05473_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand _38854_ (_06237_, _06236_, _06235_);
  nand _38855_ (_06238_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not _38856_ (_06239_, _26052_);
  nand _38857_ (_06241_, _05593_, _06239_);
  nand _38858_ (_06242_, _06241_, _06238_);
  nor _38859_ (_06243_, _06242_, _06237_);
  nand _38860_ (_06245_, _05602_, _05367_);
  nand _38861_ (_06246_, _05600_, _05115_);
  nand _38862_ (_06247_, _06246_, _06245_);
  nand _38863_ (_06248_, _05606_, _05197_);
  nand _38864_ (_06249_, _05611_, _04994_);
  nand _38865_ (_06251_, _06249_, _06248_);
  nor _38866_ (_06252_, _06251_, _06247_);
  nand _38867_ (_06253_, _06252_, _06243_);
  nand _38868_ (_06254_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _38869_ (_06255_, _05465_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand _38870_ (_06256_, _06255_, _06254_);
  nor _38871_ (_06257_, _06256_, _06253_);
  nand _38872_ (_06258_, _06257_, _06234_);
  nand _38873_ (_06259_, _06258_, _05480_);
  nand _38874_ (_06260_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _38875_ (_06261_, _06260_, _06259_);
  nor _38876_ (_06263_, _06261_, _05487_);
  nand _38877_ (_06264_, _05487_, _02229_);
  nand _38878_ (_06266_, _06264_, _26487_);
  nor _38879_ (_28381_[4], _06266_, _06263_);
  nand _38880_ (_06268_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nand _38881_ (_06269_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand _38882_ (_06271_, _06269_, _06268_);
  nand _38883_ (_06272_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand _38884_ (_06273_, _05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand _38885_ (_06274_, _06273_, _06272_);
  nor _38886_ (_06276_, _06274_, _06271_);
  nand _38887_ (_06277_, _05528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand _38888_ (_06279_, _05522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand _38889_ (_06280_, _06279_, _06277_);
  nand _38890_ (_06281_, _05534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand _38891_ (_06282_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  nand _38892_ (_06283_, _06282_, _06281_);
  nor _38893_ (_06285_, _06283_, _06280_);
  nand _38894_ (_06287_, _06285_, _06276_);
  nand _38895_ (_06289_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand _38896_ (_06290_, _05554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand _38897_ (_06291_, _06290_, _06289_);
  nand _38898_ (_06292_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand _38899_ (_06293_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand _38900_ (_06294_, _06293_, _06292_);
  nor _38901_ (_06295_, _06294_, _06291_);
  nand _38902_ (_06296_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  nand _38903_ (_06297_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nand _38904_ (_06299_, _06297_, _06296_);
  nand _38905_ (_06300_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _38906_ (_06301_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  nand _38907_ (_06303_, _06301_, _06300_);
  nor _38908_ (_06304_, _06303_, _06299_);
  nand _38909_ (_06305_, _06304_, _06295_);
  nor _38910_ (_06306_, _06305_, _06287_);
  nand _38911_ (_06307_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand _38912_ (_06308_, _05473_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand _38913_ (_06309_, _06308_, _06307_);
  nand _38914_ (_06310_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not _38915_ (_06311_, _26070_);
  nand _38916_ (_06312_, _05593_, _06311_);
  nand _38917_ (_06313_, _06312_, _06310_);
  nor _38918_ (_06314_, _06313_, _06309_);
  nand _38919_ (_06315_, _05600_, _05125_);
  nand _38920_ (_06316_, _05602_, _05340_);
  nand _38921_ (_06317_, _06316_, _06315_);
  nand _38922_ (_06318_, _05606_, _05174_);
  nand _38923_ (_06319_, _05611_, _05006_);
  nand _38924_ (_06320_, _06319_, _06318_);
  nor _38925_ (_06321_, _06320_, _06317_);
  nand _38926_ (_06322_, _06321_, _06314_);
  nand _38927_ (_06323_, _05465_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand _38928_ (_06324_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _38929_ (_06325_, _06324_, _06323_);
  nor _38930_ (_06327_, _06325_, _06322_);
  nand _38931_ (_06328_, _06327_, _06306_);
  nand _38932_ (_06329_, _06328_, _05480_);
  nand _38933_ (_06331_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _38934_ (_06332_, _06331_, _06329_);
  nor _38935_ (_06333_, _06332_, _05487_);
  nand _38936_ (_06334_, _05487_, _02307_);
  nand _38937_ (_06335_, _06334_, _26487_);
  nor _38938_ (_28381_[5], _06335_, _06333_);
  nand _38939_ (_06336_, _05487_, _04717_);
  nand _38940_ (_06337_, _06336_, _26487_);
  nand _38941_ (_06338_, _05659_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _38942_ (_06339_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand _38943_ (_06340_, _05516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand _38944_ (_06341_, _06340_, _06339_);
  nand _38945_ (_06342_, _05498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _38946_ (_06344_, _05505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _38947_ (_06345_, _06344_, _06342_);
  nor _38948_ (_06346_, _06345_, _06341_);
  nand _38949_ (_06347_, _05522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nand _38950_ (_06348_, _05528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand _38951_ (_06349_, _06348_, _06347_);
  nand _38952_ (_06350_, _05534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  nand _38953_ (_06351_, _05540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand _38954_ (_06352_, _06351_, _06350_);
  nor _38955_ (_06353_, _06352_, _06349_);
  nand _38956_ (_06355_, _06353_, _06346_);
  nand _38957_ (_06356_, _05551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nand _38958_ (_06357_, _05554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _38959_ (_06358_, _06357_, _06356_);
  nand _38960_ (_06359_, _05557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _38961_ (_06360_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _38962_ (_06361_, _06360_, _06359_);
  nor _38963_ (_06362_, _06361_, _06358_);
  nand _38964_ (_06364_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  nand _38965_ (_06366_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _38966_ (_06367_, _06366_, _06364_);
  nand _38967_ (_06368_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _38968_ (_06369_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand _38969_ (_06370_, _06369_, _06368_);
  nor _38970_ (_06371_, _06370_, _06367_);
  nand _38971_ (_06372_, _06371_, _06362_);
  nor _38972_ (_06373_, _06372_, _06355_);
  nand _38973_ (_06375_, _05484_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand _38974_ (_06376_, _05473_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand _38975_ (_06377_, _06376_, _06375_);
  nand _38976_ (_06378_, _05588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not _38977_ (_06379_, _25938_);
  nand _38978_ (_06381_, _05593_, _06379_);
  nand _38979_ (_06382_, _06381_, _06378_);
  nor _38980_ (_06383_, _06382_, _06377_);
  nand _38981_ (_06384_, _05602_, _05382_);
  nand _38982_ (_06385_, _05600_, _05101_);
  nand _38983_ (_06386_, _06385_, _06384_);
  nand _38984_ (_06387_, _05606_, _05209_);
  nand _38985_ (_06388_, _05611_, _05017_);
  nand _38986_ (_06390_, _06388_, _06387_);
  nor _38987_ (_06392_, _06390_, _06386_);
  nand _38988_ (_06393_, _06392_, _06383_);
  nand _38989_ (_06395_, _05452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _38990_ (_06397_, _05465_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _38991_ (_06398_, _06397_, _06395_);
  nor _38992_ (_06400_, _06398_, _06393_);
  nand _38993_ (_06402_, _06400_, _06373_);
  not _38994_ (_06404_, _05461_);
  nor _38995_ (_06405_, _06404_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor _38996_ (_06406_, _06405_, _05479_);
  nand _38997_ (_06407_, _06406_, _06402_);
  nand _38998_ (_06409_, _06407_, _06338_);
  nor _38999_ (_06411_, _06409_, _05487_);
  nor _39000_ (_28381_[6], _06411_, _06337_);
  nor _39001_ (_06412_, _25383_, _24862_);
  not _39002_ (_06414_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nand _39003_ (_06416_, _24862_, _06414_);
  nand _39004_ (_06417_, _06416_, _26487_);
  nor _39005_ (_28186_[5], _06417_, _06412_);
  nor _39006_ (_06418_, _27754_, _24862_);
  not _39007_ (_06419_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nand _39008_ (_06420_, _24862_, _06419_);
  nand _39009_ (_06422_, _06420_, _26487_);
  nor _39010_ (_28186_[1], _06422_, _06418_);
  nand _39011_ (_06425_, _03840_, _25039_);
  nand _39012_ (_06426_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nand _39013_ (_00560_, _06426_, _06425_);
  nand _39014_ (_06427_, _03840_, _24927_);
  nand _39015_ (_06428_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  nand _39016_ (_00569_, _06428_, _06427_);
  nand _39017_ (_06429_, _03876_, _24830_);
  nand _39018_ (_06430_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  nand _39019_ (_00574_, _06430_, _06429_);
  nor _39020_ (_06431_, _00895_, \oc8051_top_1.oc8051_decoder1.state [1]);
  nor _39021_ (_06432_, _00904_, _00899_);
  nand _39022_ (_06433_, _06432_, _06431_);
  nand _39023_ (_06434_, _06433_, _00922_);
  nor _39024_ (_06435_, _00920_, _25517_);
  nor _39025_ (_06436_, _06435_, rst);
  nand _39026_ (_28185_[0], _06436_, _06434_);
  nor _39027_ (_28183_[1], _25620_, rst);
  nor _39028_ (_06437_, rst, _23870_);
  nand _39029_ (_06438_, _06437_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _39030_ (_06439_, _25394_);
  nor _39031_ (_06440_, _25465_, _06439_);
  not _39032_ (_06441_, _06440_);
  nor _39033_ (_06442_, _06441_, _25388_);
  not _39034_ (_06443_, _06442_);
  nor _39035_ (_06445_, _06443_, _25329_);
  nand _39036_ (_06446_, _25532_, _25458_);
  not _39037_ (_06447_, _04074_);
  nor _39038_ (_06449_, _06447_, _04046_);
  nand _39039_ (_06450_, _06449_, _06446_);
  nor _39040_ (_06451_, _06450_, _06445_);
  not _39041_ (_06452_, _04079_);
  nor _39042_ (_06454_, _26203_, _25531_);
  nand _39043_ (_06456_, _06454_, _26491_);
  nor _39044_ (_06457_, _06456_, _06452_);
  nor _39045_ (_06458_, _25577_, _25465_);
  not _39046_ (_06459_, _06458_);
  nor _39047_ (_06460_, _25465_, _25426_);
  nor _39048_ (_06461_, _25803_, _25483_);
  nor _39049_ (_06462_, _06461_, _06460_);
  nand _39050_ (_06463_, _06462_, _06459_);
  nand _39051_ (_06464_, _06440_, _25388_);
  nor _39052_ (_06465_, _06464_, _25329_);
  nor _39053_ (_06466_, _06465_, _06463_);
  nand _39054_ (_06468_, _06466_, _06457_);
  nor _39055_ (_06470_, _06468_, _04045_);
  nand _39056_ (_06472_, _06470_, _06451_);
  nand _39057_ (_06473_, _06472_, _00883_);
  nand _39058_ (_28194_[0], _06473_, _06438_);
  nand _39059_ (_06475_, _03876_, _25099_);
  nand _39060_ (_06476_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nand _39061_ (_00605_, _06476_, _06475_);
  nor _39062_ (_06477_, _01065_, _25424_);
  nand _39063_ (_06478_, _06477_, _04074_);
  nor _39064_ (_06479_, _06478_, _06442_);
  nor _39065_ (_06480_, _01052_, _25584_);
  nor _39066_ (_06481_, _04954_, _04950_);
  nand _39067_ (_06482_, _06481_, _06480_);
  nor _39068_ (_06483_, _06482_, _01030_);
  nand _39069_ (_06484_, _06483_, _06479_);
  nor _39070_ (_06485_, _25803_, _25553_);
  nor _39071_ (_06486_, _26202_, _25572_);
  not _39072_ (_06488_, _06486_);
  nor _39073_ (_06489_, _06488_, _25458_);
  nor _39074_ (_06490_, _06489_, _06461_);
  not _39075_ (_06491_, _06490_);
  nor _39076_ (_06492_, _06491_, _06485_);
  nand _39077_ (_06493_, _25462_, _25596_);
  nor _39078_ (_06494_, _26195_, _25392_);
  nand _39079_ (_06495_, _01033_, _25802_);
  not _39080_ (_06496_, _06495_);
  nor _39081_ (_06497_, _06496_, _06494_);
  nand _39082_ (_06498_, _06497_, _06493_);
  nor _39083_ (_06499_, _06498_, _04953_);
  nand _39084_ (_06500_, _06499_, _06492_);
  nor _39085_ (_06501_, _06500_, _06484_);
  nor _39086_ (_06503_, _06501_, _24864_);
  not _39087_ (_06504_, _04052_);
  nand _39088_ (_06505_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _39089_ (_06506_, _06505_, _06504_);
  nor _39090_ (_06509_, _06506_, _06503_);
  nor _39091_ (_28193_[2], _06509_, rst);
  nor _39092_ (_06511_, _04046_, _25424_);
  nand _39093_ (_06513_, _06511_, _25422_);
  nand _39094_ (_06515_, _06464_, _26491_);
  nor _39095_ (_06516_, _06515_, _06513_);
  not _39096_ (_06517_, _04952_);
  not _39097_ (_06518_, _04954_);
  nor _39098_ (_06519_, _04280_, _04078_);
  nand _39099_ (_06520_, _06519_, _06518_);
  nor _39100_ (_06521_, _06520_, _06517_);
  nand _39101_ (_06522_, _06521_, _06516_);
  nor _39102_ (_06523_, _26202_, _25423_);
  nor _39103_ (_06524_, _06523_, _25574_);
  not _39104_ (_06525_, _06524_);
  nor _39105_ (_06526_, _25803_, _25403_);
  nor _39106_ (_06528_, _06526_, _26203_);
  nor _39107_ (_06530_, _04038_, _01050_);
  nand _39108_ (_06532_, _06530_, _06528_);
  nor _39109_ (_06533_, _06532_, _06525_);
  nand _39110_ (_06534_, _06533_, _06499_);
  nor _39111_ (_06535_, _06534_, _06522_);
  nor _39112_ (_06536_, _06535_, _24864_);
  not _39113_ (_06537_, _04054_);
  nand _39114_ (_06538_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _39115_ (_06539_, _06538_, _06537_);
  nor _39116_ (_06540_, _06539_, _06536_);
  nor _39117_ (_28193_[1], _06540_, rst);
  nand _39118_ (_06541_, _25802_, _25561_);
  not _39119_ (_06542_, _06541_);
  nor _39120_ (_06543_, _06542_, _25569_);
  not _39121_ (_06544_, _06543_);
  not _39122_ (_06545_, _04950_);
  nor _39123_ (_06546_, _25397_, _25235_);
  nor _39124_ (_06547_, _26202_, _25511_);
  nor _39125_ (_06548_, _06547_, _06546_);
  nand _39126_ (_06550_, _06548_, _06545_);
  nor _39127_ (_06551_, _06550_, _06544_);
  nor _39128_ (_06553_, _06465_, _06445_);
  nand _39129_ (_06554_, _06553_, _06551_);
  not _39130_ (_06555_, _25483_);
  nand _39131_ (_06556_, _06555_, _25297_);
  nand _39132_ (_06557_, _06556_, _25407_);
  not _39133_ (_06558_, _25604_);
  not _39134_ (_06559_, _04043_);
  nor _39135_ (_06560_, _06559_, _25327_);
  nor _39136_ (_06562_, _06560_, _00874_);
  nand _39137_ (_06564_, _06562_, _06558_);
  nor _39138_ (_06565_, _06564_, _06557_);
  not _39139_ (_06566_, _25562_);
  nor _39140_ (_06568_, _06566_, _25476_);
  nor _39141_ (_06569_, _06461_, _04280_);
  nand _39142_ (_06570_, _06569_, _06568_);
  nor _39143_ (_06571_, _01049_, _25390_);
  nor _39144_ (_06573_, _06571_, _25467_);
  nand _39145_ (_06575_, _06573_, _25399_);
  nor _39146_ (_06576_, _06575_, _06570_);
  nand _39147_ (_06577_, _06576_, _06565_);
  nor _39148_ (_06579_, _06577_, _06554_);
  nor _39149_ (_06580_, _06579_, _24864_);
  nand _39150_ (_06581_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _39151_ (_06582_, _06581_, _06537_);
  nor _39152_ (_06584_, _06582_, _06580_);
  nor _39153_ (_28193_[0], _06584_, rst);
  not _39154_ (_06585_, _25405_);
  nor _39155_ (_06586_, _00879_, _06585_);
  nor _39156_ (_06587_, _06586_, _00874_);
  not _39157_ (_06588_, _06587_);
  nor _39158_ (_06589_, _25403_, _25482_);
  nor _39159_ (_06590_, _06589_, _06588_);
  not _39160_ (_06592_, _06590_);
  nand _39161_ (_28184_[0], _00883_, _06592_);
  not _39162_ (_06593_, _00877_);
  nand _39163_ (_28184_[1], _00883_, _06593_);
  nand _39164_ (_06594_, _06437_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _39165_ (_06596_, _06465_, _01028_);
  nand _39166_ (_06597_, _06596_, _06490_);
  not _39167_ (_06598_, _06530_);
  nor _39168_ (_06599_, _25467_, _25417_);
  nand _39169_ (_06600_, _06599_, _04079_);
  nor _39170_ (_06601_, _06600_, _06598_);
  nor _39171_ (_06603_, _25412_, _06439_);
  nor _39172_ (_06604_, _06603_, _06460_);
  nand _39173_ (_06605_, _25421_, _25329_);
  not _39174_ (_06606_, _06605_);
  nor _39175_ (_06607_, _26201_, _25236_);
  nor _39176_ (_06608_, _06607_, _25511_);
  nor _39177_ (_06609_, _06608_, _06606_);
  nand _39178_ (_06610_, _06609_, _06604_);
  not _39179_ (_06611_, _26206_);
  nand _39180_ (_06612_, _26194_, _01061_);
  nand _39181_ (_06613_, _06612_, _06611_);
  nor _39182_ (_06614_, _06613_, _01022_);
  nand _39183_ (_06615_, _06614_, _25575_);
  nor _39184_ (_06616_, _06615_, _06610_);
  nand _39185_ (_06617_, _06616_, _06601_);
  nor _39186_ (_06618_, _06617_, _06597_);
  nand _39187_ (_06619_, _06618_, _06451_);
  nand _39188_ (_06620_, _06619_, _00883_);
  nand _39189_ (_28192_[0], _06620_, _06594_);
  nand _39190_ (_06621_, _03840_, _28096_);
  nand _39191_ (_06622_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  nand _39192_ (_00673_, _06622_, _06621_);
  not _39193_ (_06623_, _06528_);
  nand _39194_ (_06624_, _06495_, _04050_);
  nor _39195_ (_06625_, _06624_, _06623_);
  nand _39196_ (_06626_, _06625_, _06492_);
  nor _39197_ (_06628_, _04954_, _04041_);
  not _39198_ (_06629_, _06628_);
  nor _39199_ (_06630_, _06440_, _04046_);
  nand _39200_ (_06632_, _04280_, _25459_);
  nand _39201_ (_06633_, _06632_, _06630_);
  nor _39202_ (_06635_, _06633_, _06629_);
  not _39203_ (_06636_, _01042_);
  nor _39204_ (_06637_, _06636_, _25400_);
  nor _39205_ (_06639_, _06637_, _06546_);
  not _39206_ (_06640_, _25417_);
  nand _39207_ (_06641_, _04053_, _06640_);
  nor _39208_ (_06642_, _25561_, _25489_);
  nor _39209_ (_06644_, _06642_, _25465_);
  nor _39210_ (_06645_, _06644_, _06641_);
  nand _39211_ (_06647_, _06645_, _06639_);
  nor _39212_ (_06648_, _26195_, _00875_);
  nor _39213_ (_06649_, _06648_, _01035_);
  nand _39214_ (_06651_, _06649_, _25603_);
  nor _39215_ (_06653_, _06651_, _04276_);
  not _39216_ (_06654_, _25477_);
  nor _39217_ (_06656_, _25586_, _06654_);
  nand _39218_ (_06657_, _06656_, _06653_);
  nor _39219_ (_06658_, _06657_, _06647_);
  nand _39220_ (_06659_, _06658_, _06635_);
  nor _39221_ (_06660_, _06659_, _06626_);
  nor _39222_ (_06662_, _06660_, _24864_);
  nand _39223_ (_06663_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _39224_ (_06664_, _06590_, _00100_);
  nor _39225_ (_06665_, _06664_, _25807_);
  nand _39226_ (_06667_, _06665_, _06663_);
  nor _39227_ (_06668_, _06667_, _06662_);
  nor _39228_ (_28191_[1], _06668_, rst);
  not _39229_ (_06671_, _01046_);
  nand _39230_ (_06672_, _06671_, _26796_);
  nor _39231_ (_06673_, _06672_, _06641_);
  nand _39232_ (_06675_, _01033_, _25550_);
  nand _39233_ (_06677_, _06636_, _06675_);
  nor _39234_ (_06678_, _25803_, _25473_);
  nor _39235_ (_06679_, _06678_, _01055_);
  nand _39236_ (_06680_, _06679_, _06541_);
  nor _39237_ (_06681_, _06680_, _06677_);
  nand _39238_ (_06682_, _06681_, _06673_);
  not _39239_ (_06683_, _06562_);
  nand _39240_ (_06685_, _25485_, _25393_);
  not _39241_ (_06686_, _01021_);
  nand _39242_ (_06687_, _06686_, _06685_);
  nor _39243_ (_06688_, _06687_, _06683_);
  nand _39244_ (_06689_, _06688_, _06628_);
  nor _39245_ (_06690_, _06689_, _06682_);
  not _39246_ (_06691_, _25592_);
  nor _39247_ (_06692_, _25803_, _25470_);
  nor _39248_ (_06693_, _06692_, _06691_);
  nor _39249_ (_06694_, _25803_, _25577_);
  nor _39250_ (_06695_, _06440_, _06694_);
  nand _39251_ (_06697_, _06695_, _06693_);
  nor _39252_ (_06698_, _06697_, _06550_);
  nand _39253_ (_06700_, _06698_, _06690_);
  nor _39254_ (_06701_, _06700_, _06626_);
  nor _39255_ (_06703_, _06701_, _24864_);
  nand _39256_ (_06704_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _39257_ (_06705_, _06704_, _06665_);
  nor _39258_ (_06706_, _06705_, _06703_);
  nor _39259_ (_28191_[0], _06706_, rst);
  nand _39260_ (_06709_, _03840_, _25203_);
  nand _39261_ (_06711_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  nand _39262_ (_00700_, _06711_, _06709_);
  not _39263_ (_06712_, _23998_);
  nor _39264_ (_06713_, _04089_, _25929_);
  nand _39265_ (_06714_, _06713_, _26058_);
  nand _39266_ (_06715_, _04089_, _26472_);
  nand _39267_ (_06716_, _06715_, _06714_);
  not _39268_ (_06717_, _06716_);
  nor _39269_ (_06718_, _06717_, _06712_);
  nor _39270_ (_06719_, _06716_, _23998_);
  nor _39271_ (_06720_, _06719_, _06718_);
  not _39272_ (_06721_, _06720_);
  nor _39273_ (_06723_, _06713_, _25991_);
  nor _39274_ (_06724_, _06723_, _24885_);
  nand _39275_ (_06726_, _06723_, _24885_);
  not _39276_ (_06728_, _06726_);
  nor _39277_ (_06730_, _06728_, _06724_);
  nor _39278_ (_06731_, _06713_, _26059_);
  nor _39279_ (_06732_, _06731_, _24065_);
  nor _39280_ (_06733_, _06713_, _26126_);
  not _39281_ (_06734_, _06733_);
  nand _39282_ (_06735_, _06734_, _24061_);
  not _39283_ (_06737_, _06735_);
  nor _39284_ (_06738_, _06737_, _06732_);
  nand _39285_ (_06739_, _06738_, _06730_);
  nor _39286_ (_06740_, _06739_, _06721_);
  not _39287_ (_06741_, _24053_);
  not _39288_ (_06743_, _04089_);
  nand _39289_ (_06744_, _06743_, _25843_);
  nor _39290_ (_06745_, _06744_, _26124_);
  nor _39291_ (_06747_, _06743_, _26403_);
  nor _39292_ (_06748_, _06747_, _06745_);
  nor _39293_ (_06749_, _06748_, _06741_);
  not _39294_ (_06751_, _06748_);
  nor _39295_ (_06753_, _06751_, _24053_);
  nor _39296_ (_06755_, _06753_, _06749_);
  not _39297_ (_06756_, _24019_);
  nor _39298_ (_06758_, _06744_, _25993_);
  nor _39299_ (_06759_, _06713_, _25919_);
  nor _39300_ (_06760_, _06759_, _06758_);
  not _39301_ (_06761_, _06760_);
  nor _39302_ (_06763_, _06761_, _06756_);
  nor _39303_ (_06764_, _06760_, _24019_);
  nor _39304_ (_06765_, _06764_, _06763_);
  nand _39305_ (_06766_, _06765_, _06755_);
  not _39306_ (_06767_, _23960_);
  nor _39307_ (_06768_, _06744_, _25916_);
  nand _39308_ (_06769_, _04089_, _26338_);
  not _39309_ (_06770_, _06769_);
  nor _39310_ (_06771_, _06770_, _06768_);
  nor _39311_ (_06772_, _06771_, _06767_);
  nand _39312_ (_06773_, _06713_, _25919_);
  nand _39313_ (_06774_, _06769_, _06773_);
  nor _39314_ (_06775_, _06774_, _23960_);
  nor _39315_ (_06776_, _06775_, _06772_);
  nor _39316_ (_06777_, _06734_, _24061_);
  nor _39317_ (_06778_, _25931_, _23918_);
  not _39318_ (_06779_, _06778_);
  not _39319_ (_06780_, _06731_);
  nor _39320_ (_06781_, _06780_, _24064_);
  nor _39321_ (_06783_, _06781_, _06779_);
  not _39322_ (_06784_, _06783_);
  nor _39323_ (_06786_, _06784_, _06777_);
  nand _39324_ (_06787_, _06786_, _06776_);
  nor _39325_ (_06788_, _06787_, _06766_);
  nand _39326_ (_06790_, _06788_, _06740_);
  nor _39327_ (_28232_, _06790_, rst);
  nor _39328_ (_28233_[7], _24788_, rst);
  nor _39329_ (_28235_[2], _26403_, rst);
  nand _39330_ (_06793_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  nand _39331_ (_06794_, _05864_, _25099_);
  nand _39332_ (_00748_, _06794_, _06793_);
  nor _39333_ (_06795_, _00430_, _00227_);
  not _39334_ (_06796_, _06795_);
  nor _39335_ (_06797_, _06796_, _24716_);
  nor _39336_ (_06798_, _06795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor _39337_ (_06800_, _06798_, _06797_);
  nor _39338_ (_06801_, _06800_, _00441_);
  nand _39339_ (_06802_, _00441_, _25625_);
  nand _39340_ (_06804_, _06802_, _26487_);
  nor _39341_ (_00821_, _06804_, _06801_);
  nor _39342_ (_28233_[0], _24829_, rst);
  nor _39343_ (_28233_[1], _25098_, rst);
  nor _39344_ (_28233_[2], _28095_, rst);
  nor _39345_ (_28233_[3], _25202_, rst);
  nor _39346_ (_28233_[4], _25038_, rst);
  nor _39347_ (_28233_[5], _24926_, rst);
  nor _39348_ (_28233_[6], _25149_, rst);
  nor _39349_ (_06807_, _00629_, _24073_);
  not _39350_ (_06808_, _06807_);
  nand _39351_ (_06809_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  nand _39352_ (_06810_, _06807_, _24927_);
  nand _39353_ (_00886_, _06810_, _06809_);
  nor _39354_ (_28235_[0], _26407_, rst);
  nor _39355_ (_28235_[1], _26473_, rst);
  nor _39356_ (_06814_, _25322_, _24862_);
  not _39357_ (_06816_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nand _39358_ (_06818_, _24862_, _06816_);
  nand _39359_ (_06820_, _06818_, _26487_);
  nor _39360_ (_28186_[4], _06820_, _06814_);
  nor _39361_ (_06821_, _27724_, _24862_);
  not _39362_ (_06822_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nand _39363_ (_06823_, _24862_, _06822_);
  nand _39364_ (_06825_, _06823_, _26487_);
  nor _39365_ (_28186_[3], _06825_, _06821_);
  nor _39366_ (_06826_, _00954_, _25165_);
  nand _39367_ (_06827_, _06826_, _25099_);
  not _39368_ (_06828_, _06826_);
  nand _39369_ (_06829_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  nand _39370_ (_00907_, _06829_, _06827_);
  not _39371_ (_06830_, _25523_);
  nor _39372_ (_28183_[0], _06830_, rst);
  nor _39373_ (_06833_, _25453_, _24862_);
  not _39374_ (_06834_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nand _39375_ (_06835_, _24862_, _06834_);
  nand _39376_ (_06836_, _06835_, _26487_);
  nor _39377_ (_28186_[0], _06836_, _06833_);
  nor _39378_ (_06837_, _25290_, _24862_);
  not _39379_ (_06838_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nand _39380_ (_06840_, _24862_, _06838_);
  nand _39381_ (_06842_, _06840_, _26487_);
  nor _39382_ (_28186_[2], _06842_, _06837_);
  nor _39383_ (_06843_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _39384_ (_06844_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _28020_);
  nor _39385_ (_06845_, _06844_, _06843_);
  not _39386_ (_06846_, _06845_);
  nor _39387_ (_06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _39388_ (_06848_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _28020_);
  nor _39389_ (_06849_, _06848_, _06847_);
  not _39390_ (_06850_, _06849_);
  nor _39391_ (_06851_, _06850_, _06846_);
  not _39392_ (_06852_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _39393_ (_06853_, _02112_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _39394_ (_06854_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _28020_);
  nor _39395_ (_06855_, _06854_, _06853_);
  nor _39396_ (_06856_, _02182_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _39397_ (_06857_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _28020_);
  nor _39398_ (_06858_, _06857_, _06856_);
  nor _39399_ (_06859_, _06858_, _06855_);
  not _39400_ (_06860_, _06859_);
  nor _39401_ (_06861_, _06860_, _06852_);
  not _39402_ (_06862_, \oc8051_symbolic_cxrom1.regvalid [15]);
  not _39403_ (_06863_, _06855_);
  not _39404_ (_06864_, _06858_);
  nor _39405_ (_06865_, _06864_, _06863_);
  not _39406_ (_06867_, _06865_);
  nor _39407_ (_06868_, _06867_, _06862_);
  nor _39408_ (_06869_, _06868_, _06861_);
  not _39409_ (_06871_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _39410_ (_06872_, _06864_, _06855_);
  not _39411_ (_06873_, _06872_);
  nor _39412_ (_06875_, _06873_, _06871_);
  not _39413_ (_06876_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _39414_ (_06877_, _06858_, _06863_);
  not _39415_ (_06878_, _06877_);
  nor _39416_ (_06879_, _06878_, _06876_);
  nor _39417_ (_06880_, _06879_, _06875_);
  nand _39418_ (_06881_, _06880_, _06869_);
  nand _39419_ (_06882_, _06881_, _06851_);
  not _39420_ (_06883_, _06882_);
  nor _39421_ (_06885_, _06849_, _06846_);
  not _39422_ (_06886_, _06885_);
  not _39423_ (_06888_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _39424_ (_06889_, _06858_, _06888_);
  not _39425_ (_06891_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _39426_ (_06892_, _06864_, _06891_);
  nor _39427_ (_06893_, _06892_, _06889_);
  nor _39428_ (_06894_, _06893_, _06863_);
  not _39429_ (_06895_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _39430_ (_06896_, _06873_, _06895_);
  not _39431_ (_06897_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _39432_ (_06898_, _06860_, _06897_);
  nor _39433_ (_06899_, _06898_, _06896_);
  not _39434_ (_06900_, _06899_);
  nor _39435_ (_06902_, _06900_, _06894_);
  nor _39436_ (_06904_, _06902_, _06886_);
  nor _39437_ (_06905_, _06904_, _06883_);
  nor _39438_ (_06906_, _06849_, _06845_);
  not _39439_ (_06907_, _06906_);
  not _39440_ (_06909_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _39441_ (_06910_, _06860_, _06909_);
  not _39442_ (_06912_, _06910_);
  nand _39443_ (_06913_, _06865_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand _39444_ (_06914_, _06913_, _06912_);
  not _39445_ (_06915_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _39446_ (_06916_, _06873_, _06915_);
  not _39447_ (_06917_, _06916_);
  nand _39448_ (_06919_, _06877_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand _39449_ (_06920_, _06919_, _06917_);
  nor _39450_ (_06922_, _06920_, _06914_);
  nor _39451_ (_06923_, _06922_, _06907_);
  nor _39452_ (_06924_, _06850_, _06845_);
  not _39453_ (_06925_, _06924_);
  nor _39454_ (_06926_, _06864_, \oc8051_symbolic_cxrom1.regvalid [14]);
  not _39455_ (_06928_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand _39456_ (_06929_, _06864_, _06928_);
  nand _39457_ (_06930_, _06929_, _06855_);
  nor _39458_ (_06931_, _06930_, _06926_);
  not _39459_ (_06932_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _39460_ (_06934_, _06873_, _06932_);
  not _39461_ (_06935_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _39462_ (_06936_, _06860_, _06935_);
  nor _39463_ (_06937_, _06936_, _06934_);
  not _39464_ (_06938_, _06937_);
  nor _39465_ (_06939_, _06938_, _06931_);
  nor _39466_ (_06941_, _06939_, _06925_);
  nor _39467_ (_06943_, _06941_, _06923_);
  nand _39468_ (_06944_, _06943_, _06905_);
  nor _39469_ (_06945_, _06846_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor _39470_ (_06947_, _06845_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor _39471_ (_06948_, _06947_, _06945_);
  nand _39472_ (_06950_, _06948_, _06849_);
  nor _39473_ (_06951_, _06846_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor _39474_ (_06952_, _06845_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _39475_ (_06953_, _06952_, _06951_);
  nand _39476_ (_06955_, _06953_, _06850_);
  nand _39477_ (_06957_, _06955_, _06950_);
  nand _39478_ (_06958_, _06957_, _06863_);
  nor _39479_ (_06959_, _06863_, _06850_);
  not _39480_ (_06960_, _06959_);
  nor _39481_ (_06962_, _06846_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor _39482_ (_06964_, _06845_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nor _39483_ (_06966_, _06964_, _06962_);
  not _39484_ (_06967_, _06966_);
  nor _39485_ (_06968_, _06967_, _06960_);
  nor _39486_ (_06969_, _06863_, _06849_);
  not _39487_ (_06970_, _06969_);
  nor _39488_ (_06971_, _06846_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _39489_ (_06972_, _06845_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _39490_ (_06974_, _06972_, _06971_);
  not _39491_ (_06975_, _06974_);
  nor _39492_ (_06976_, _06975_, _06970_);
  nor _39493_ (_06977_, _06976_, _06968_);
  nand _39494_ (_06978_, _06977_, _06958_);
  nand _39495_ (_06979_, _06978_, _06858_);
  nor _39496_ (_06980_, _06846_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor _39497_ (_06981_, _06845_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor _39498_ (_06982_, _06981_, _06980_);
  nand _39499_ (_06983_, _06982_, _06849_);
  nor _39500_ (_06984_, _06846_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _39501_ (_06985_, _06845_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _39502_ (_06986_, _06985_, _06984_);
  nand _39503_ (_06988_, _06986_, _06850_);
  nand _39504_ (_06989_, _06988_, _06983_);
  nand _39505_ (_06990_, _06989_, _06863_);
  nor _39506_ (_06992_, _06846_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _39507_ (_06993_, _06845_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _39508_ (_06994_, _06993_, _06992_);
  nand _39509_ (_06995_, _06994_, _06850_);
  nor _39510_ (_06997_, _06846_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nor _39511_ (_06998_, _06845_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nor _39512_ (_06999_, _06998_, _06997_);
  nand _39513_ (_07000_, _06999_, _06849_);
  nand _39514_ (_07001_, _07000_, _06995_);
  nand _39515_ (_07003_, _07001_, _06855_);
  nand _39516_ (_07004_, _07003_, _06990_);
  nand _39517_ (_07005_, _07004_, _06864_);
  nand _39518_ (_07006_, _07005_, _06979_);
  nand _39519_ (_07007_, _07006_, _06944_);
  not _39520_ (_07009_, _06944_);
  nand _39521_ (_07010_, _07009_, word_in[7]);
  nand _39522_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07010_, _07007_);
  not _39523_ (_07011_, _06851_);
  nor _39524_ (_07012_, _06863_, _07011_);
  nor _39525_ (_07013_, _07012_, _06864_);
  not _39526_ (_07014_, _07012_);
  nor _39527_ (_07015_, _07014_, _06858_);
  nor _39528_ (_07017_, _07015_, _07013_);
  not _39529_ (_07019_, _07017_);
  nor _39530_ (_07020_, _06855_, _06851_);
  nor _39531_ (_07022_, _07020_, _07012_);
  nor _39532_ (_07023_, _07022_, _07019_);
  not _39533_ (_07025_, _07023_);
  nor _39534_ (_07027_, _07025_, _06852_);
  nor _39535_ (_07029_, _07017_, \oc8051_symbolic_cxrom1.regvalid [15]);
  not _39536_ (_07030_, _07022_);
  nor _39537_ (_07032_, _07030_, _06864_);
  nor _39538_ (_07033_, _07030_, _06876_);
  nor _39539_ (_07034_, _07033_, _07032_);
  nor _39540_ (_07036_, _07034_, _07029_);
  nor _39541_ (_07037_, _07022_, _07017_);
  not _39542_ (_07038_, _07037_);
  nor _39543_ (_07039_, _07038_, _06871_);
  nor _39544_ (_07040_, _07039_, _07036_);
  not _39545_ (_07042_, _07040_);
  nor _39546_ (_07044_, _07042_, _07027_);
  nor _39547_ (_07045_, _07044_, _06925_);
  nor _39548_ (_07046_, _07025_, _06897_);
  nor _39549_ (_07048_, _07017_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _39550_ (_07050_, _07030_, _06888_);
  nor _39551_ (_07051_, _07050_, _07032_);
  nor _39552_ (_07053_, _07051_, _07048_);
  nor _39553_ (_07054_, _07038_, _06895_);
  nor _39554_ (_07055_, _07054_, _07053_);
  not _39555_ (_07056_, _07055_);
  nor _39556_ (_07057_, _07056_, _07046_);
  nor _39557_ (_07058_, _07057_, _06907_);
  nor _39558_ (_07059_, _07058_, _07045_);
  nor _39559_ (_07060_, _07025_, _06935_);
  nor _39560_ (_07062_, _07017_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _39561_ (_07063_, _07030_, _06928_);
  nor _39562_ (_07064_, _07063_, _07032_);
  nor _39563_ (_07065_, _07064_, _07062_);
  nor _39564_ (_07066_, _07038_, _06932_);
  nor _39565_ (_07068_, _07066_, _07065_);
  not _39566_ (_07069_, _07068_);
  nor _39567_ (_07071_, _07069_, _07060_);
  nor _39568_ (_07072_, _07071_, _06886_);
  nor _39569_ (_07073_, _07025_, _06909_);
  nor _39570_ (_07075_, _07019_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _39571_ (_07076_, _06864_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _39572_ (_07077_, _07030_, _07076_);
  not _39573_ (_07079_, _07077_);
  nor _39574_ (_07080_, _07079_, _07075_);
  nor _39575_ (_07082_, _07038_, _06915_);
  nor _39576_ (_07083_, _07082_, _07080_);
  not _39577_ (_07084_, _07083_);
  nor _39578_ (_07086_, _07084_, _07073_);
  nor _39579_ (_07088_, _07086_, _07011_);
  nor _39580_ (_07090_, _07088_, _07072_);
  nand _39581_ (_07091_, _07090_, _07059_);
  nor _39582_ (_07093_, _06924_, _06885_);
  nor _39583_ (_07095_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _39584_ (_07096_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor _39585_ (_07097_, _07096_, _07095_);
  nand _39586_ (_07098_, _07097_, _07093_);
  not _39587_ (_07100_, _07093_);
  nor _39588_ (_07101_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor _39589_ (_07102_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor _39590_ (_07104_, _07102_, _07101_);
  nand _39591_ (_07105_, _07104_, _07100_);
  nand _39592_ (_07106_, _07105_, _07098_);
  nand _39593_ (_07107_, _07106_, _07037_);
  nor _39594_ (_07108_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor _39595_ (_07109_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor _39596_ (_07110_, _07109_, _07108_);
  not _39597_ (_07111_, _07110_);
  nor _39598_ (_07112_, _07111_, _07093_);
  nor _39599_ (_07113_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _39600_ (_07114_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _39601_ (_07115_, _07114_, _07113_);
  not _39602_ (_07116_, _07115_);
  nor _39603_ (_07117_, _07116_, _07100_);
  nor _39604_ (_07118_, _07117_, _07112_);
  nor _39605_ (_07119_, _07118_, _07025_);
  nor _39606_ (_07121_, _07030_, _06858_);
  nor _39607_ (_07122_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nor _39608_ (_07123_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nor _39609_ (_07124_, _07123_, _07122_);
  nand _39610_ (_07126_, _07124_, _07100_);
  nor _39611_ (_07127_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _39612_ (_07129_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _39613_ (_07130_, _07129_, _07127_);
  nand _39614_ (_07132_, _07130_, _07093_);
  nand _39615_ (_07134_, _07132_, _07126_);
  nand _39616_ (_07135_, _07134_, _07121_);
  nor _39617_ (_07136_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _39618_ (_07138_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _39619_ (_07139_, _07138_, _07136_);
  nand _39620_ (_07141_, _07139_, _07093_);
  nor _39621_ (_07142_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nor _39622_ (_07144_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor _39623_ (_07145_, _07144_, _07142_);
  nand _39624_ (_07146_, _07145_, _07100_);
  nand _39625_ (_07148_, _07146_, _07141_);
  nand _39626_ (_07150_, _07148_, _07032_);
  nand _39627_ (_07152_, _07150_, _07135_);
  nor _39628_ (_07153_, _07152_, _07119_);
  nand _39629_ (_07155_, _07153_, _07107_);
  nand _39630_ (_07156_, _07155_, _07091_);
  not _39631_ (_07157_, _07091_);
  nand _39632_ (_07159_, _07157_, word_in[15]);
  nand _39633_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07159_, _07156_);
  nor _39634_ (_07160_, _06878_, _06850_);
  nor _39635_ (_07162_, _06959_, _06864_);
  nor _39636_ (_07163_, _07162_, _07160_);
  nor _39637_ (_07164_, _06855_, _06850_);
  nor _39638_ (_07166_, _07164_, _06969_);
  not _39639_ (_07167_, _07166_);
  nor _39640_ (_07168_, _07167_, _07163_);
  not _39641_ (_07169_, _07168_);
  nor _39642_ (_07170_, _07169_, _06932_);
  nor _39643_ (_07171_, _07163_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _39644_ (_07172_, _07166_, _06864_);
  nor _39645_ (_07174_, _07166_, _06928_);
  nor _39646_ (_07175_, _07174_, _07172_);
  nor _39647_ (_07177_, _07175_, _07171_);
  not _39648_ (_07178_, _07163_);
  nor _39649_ (_07179_, _07167_, _07178_);
  not _39650_ (_07181_, _07179_);
  nor _39651_ (_07182_, _07181_, _06935_);
  nor _39652_ (_07183_, _07182_, _07177_);
  not _39653_ (_07184_, _07183_);
  nor _39654_ (_07185_, _07184_, _07170_);
  nor _39655_ (_07186_, _07185_, _06907_);
  nor _39656_ (_07188_, _07181_, _06852_);
  nor _39657_ (_07189_, _07163_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _39658_ (_07190_, _07166_, _06876_);
  nor _39659_ (_07191_, _07190_, _07172_);
  nor _39660_ (_07192_, _07191_, _07189_);
  nor _39661_ (_07193_, _07169_, _06871_);
  nor _39662_ (_07194_, _07193_, _07192_);
  not _39663_ (_07196_, _07194_);
  nor _39664_ (_07197_, _07196_, _07188_);
  nor _39665_ (_07198_, _07197_, _06886_);
  nor _39666_ (_07200_, _07198_, _07186_);
  nor _39667_ (_07201_, _07181_, _06897_);
  nor _39668_ (_07202_, _07163_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _39669_ (_07204_, _07166_, _06888_);
  nor _39670_ (_07205_, _07204_, _07172_);
  nor _39671_ (_07206_, _07205_, _07202_);
  nor _39672_ (_07208_, _07169_, _06895_);
  nor _39673_ (_07209_, _07208_, _07206_);
  not _39674_ (_07210_, _07209_);
  nor _39675_ (_07211_, _07210_, _07201_);
  nor _39676_ (_07212_, _07211_, _07011_);
  nor _39677_ (_07213_, _07181_, _06909_);
  nor _39678_ (_07214_, _07178_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _39679_ (_07215_, _07166_, _07076_);
  not _39680_ (_07216_, _07215_);
  nor _39681_ (_07217_, _07216_, _07214_);
  nor _39682_ (_07218_, _07169_, _06915_);
  nor _39683_ (_07219_, _07218_, _07217_);
  not _39684_ (_07220_, _07219_);
  nor _39685_ (_07221_, _07220_, _07213_);
  nor _39686_ (_07223_, _07221_, _06925_);
  nor _39687_ (_07225_, _07223_, _07212_);
  nand _39688_ (_07226_, _07225_, _07200_);
  not _39689_ (_07227_, _07226_);
  nand _39690_ (_07228_, _07227_, word_in[23]);
  nor _39691_ (_07229_, _06953_, _06850_);
  nor _39692_ (_07230_, _06948_, _06849_);
  nor _39693_ (_07232_, _07230_, _07229_);
  nand _39694_ (_07234_, _07232_, _07166_);
  nor _39695_ (_07235_, _06970_, _06967_);
  not _39696_ (_07236_, _07164_);
  nor _39697_ (_07237_, _06975_, _07236_);
  nor _39698_ (_07238_, _07237_, _07235_);
  nand _39699_ (_07239_, _07238_, _07234_);
  nand _39700_ (_07240_, _07239_, _07178_);
  nor _39701_ (_07241_, _06982_, _06849_);
  nor _39702_ (_07242_, _06986_, _06850_);
  nor _39703_ (_07243_, _07242_, _07241_);
  nand _39704_ (_07244_, _07243_, _07166_);
  nand _39705_ (_07245_, _06994_, _06849_);
  nand _39706_ (_07246_, _06999_, _06850_);
  nand _39707_ (_07247_, _07246_, _07245_);
  nand _39708_ (_07248_, _07247_, _07167_);
  nand _39709_ (_07249_, _07248_, _07244_);
  nand _39710_ (_07250_, _07249_, _07163_);
  nand _39711_ (_07251_, _07250_, _07240_);
  nand _39712_ (_07252_, _07251_, _07226_);
  nand _39713_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07252_, _07228_);
  nor _39714_ (_07254_, _06906_, _06863_);
  not _39715_ (_07255_, _07254_);
  nor _39716_ (_07257_, _07255_, _06864_);
  nor _39717_ (_07258_, _07254_, _06858_);
  nor _39718_ (_07259_, _07258_, _07257_);
  nor _39719_ (_07260_, _07259_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _39720_ (_07262_, _06907_, _06855_);
  nor _39721_ (_07263_, _07262_, _07254_);
  not _39722_ (_07264_, _07263_);
  nor _39723_ (_07265_, _07264_, _06926_);
  not _39724_ (_07266_, _07265_);
  nor _39725_ (_07268_, _07266_, _07260_);
  nor _39726_ (_07269_, _07259_, _06935_);
  not _39727_ (_07271_, _07259_);
  nor _39728_ (_07273_, _07271_, _06932_);
  nor _39729_ (_07274_, _07273_, _07269_);
  nor _39730_ (_07275_, _07274_, _07263_);
  nor _39731_ (_07277_, _07275_, _07268_);
  nor _39732_ (_07279_, _07277_, _07011_);
  nor _39733_ (_07281_, _07259_, _06852_);
  nor _39734_ (_07282_, _07271_, _06871_);
  nor _39735_ (_07283_, _07282_, _07281_);
  nor _39736_ (_07284_, _07283_, _07263_);
  nor _39737_ (_07286_, _07259_, _06876_);
  nor _39738_ (_07287_, _07271_, _06862_);
  nor _39739_ (_07288_, _07287_, _07286_);
  nor _39740_ (_07290_, _07288_, _07264_);
  nor _39741_ (_07291_, _07290_, _07284_);
  nor _39742_ (_07292_, _07291_, _06907_);
  nor _39743_ (_07293_, _07292_, _07279_);
  nor _39744_ (_07294_, _07259_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _39745_ (_07296_, _07264_, _07076_);
  not _39746_ (_07298_, _07296_);
  nor _39747_ (_07299_, _07298_, _07294_);
  nor _39748_ (_07301_, _07259_, _06909_);
  nor _39749_ (_07302_, _07271_, _06915_);
  nor _39750_ (_07303_, _07302_, _07301_);
  nor _39751_ (_07304_, _07303_, _07263_);
  nor _39752_ (_07305_, _07304_, _07299_);
  nor _39753_ (_07306_, _07305_, _06886_);
  nor _39754_ (_07308_, _07259_, _06897_);
  nor _39755_ (_07309_, _07271_, _06895_);
  nor _39756_ (_07310_, _07309_, _07308_);
  nor _39757_ (_07312_, _07310_, _07263_);
  nor _39758_ (_07313_, _07259_, _06888_);
  nor _39759_ (_07315_, _07271_, _06891_);
  nor _39760_ (_07316_, _07315_, _07313_);
  nor _39761_ (_07318_, _07316_, _07264_);
  nor _39762_ (_07320_, _07318_, _07312_);
  nor _39763_ (_07321_, _07320_, _06925_);
  nor _39764_ (_07323_, _07321_, _07306_);
  nand _39765_ (_07324_, _07323_, _07293_);
  nand _39766_ (_07325_, _07145_, _07093_);
  nand _39767_ (_07326_, _07139_, _07100_);
  nand _39768_ (_07327_, _07326_, _07325_);
  nand _39769_ (_07328_, _07327_, _07263_);
  nand _39770_ (_07330_, _07097_, _07100_);
  nand _39771_ (_07331_, _07104_, _07093_);
  nand _39772_ (_07332_, _07331_, _07330_);
  nand _39773_ (_07334_, _07332_, _07264_);
  nand _39774_ (_07336_, _07334_, _07328_);
  nand _39775_ (_07337_, _07336_, _07259_);
  nand _39776_ (_07339_, _07124_, _07093_);
  nand _39777_ (_07340_, _07130_, _07100_);
  nand _39778_ (_07341_, _07340_, _07339_);
  nand _39779_ (_07342_, _07341_, _07263_);
  nand _39780_ (_07344_, _07110_, _07093_);
  nand _39781_ (_07345_, _07115_, _07100_);
  nand _39782_ (_07346_, _07345_, _07344_);
  nand _39783_ (_07348_, _07346_, _07264_);
  nand _39784_ (_07349_, _07348_, _07342_);
  nand _39785_ (_07350_, _07349_, _07271_);
  nand _39786_ (_07351_, _07350_, _07337_);
  nand _39787_ (_07352_, _07351_, _07324_);
  not _39788_ (_07354_, _07324_);
  nand _39789_ (_07355_, _07354_, word_in[31]);
  nand _39790_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _07355_, _07352_);
  not _39791_ (_07357_, _07172_);
  nor _39792_ (_07359_, _07226_, rst);
  not _39793_ (_07361_, _07359_);
  nor _39794_ (_07362_, _07361_, _07357_);
  not _39795_ (_07363_, _07362_);
  nor _39796_ (_07364_, _07363_, _06886_);
  not _39797_ (_07365_, _07364_);
  nor _39798_ (_07366_, _07091_, rst);
  not _39799_ (_07367_, _07366_);
  nor _39800_ (_07368_, _07367_, _07030_);
  nand _39801_ (_07369_, _07368_, _07019_);
  nor _39802_ (_07370_, _07369_, _06925_);
  not _39803_ (_07371_, _07370_);
  not _39804_ (_07372_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor _39805_ (_07373_, _07014_, _06864_);
  not _39806_ (_07374_, _07373_);
  nor _39807_ (_07375_, _06944_, rst);
  not _39808_ (_07376_, _07375_);
  nor _39809_ (_07377_, _07376_, _07374_);
  not _39810_ (_07378_, _07377_);
  nand _39811_ (_07379_, _07378_, _07372_);
  not _39812_ (_07381_, word_in[7]);
  nand _39813_ (_07383_, _07377_, _07381_);
  nand _39814_ (_07385_, _07383_, _07379_);
  nand _39815_ (_07386_, _07385_, _07371_);
  not _39816_ (_07387_, word_in[15]);
  nand _39817_ (_07388_, _07370_, _07387_);
  nand _39818_ (_07389_, _07388_, _07386_);
  nand _39819_ (_07391_, _07389_, _07365_);
  nor _39820_ (_07392_, _07324_, rst);
  not _39821_ (_07393_, _07392_);
  nor _39822_ (_07394_, _07393_, _07271_);
  not _39823_ (_07395_, _07394_);
  nor _39824_ (_07396_, _07395_, _07264_);
  not _39825_ (_07398_, _07396_);
  nor _39826_ (_07399_, _07398_, _06907_);
  nor _39827_ (_07400_, _07228_, rst);
  nor _39828_ (_07402_, _07400_, _07365_);
  nor _39829_ (_07404_, _07402_, _07399_);
  nand _39830_ (_07406_, _07404_, _07391_);
  nor _39831_ (_07408_, _07355_, rst);
  nand _39832_ (_07409_, _07408_, _07399_);
  nand _39833_ (_28173_[7], _07409_, _07406_);
  not _39834_ (_07412_, _07262_);
  nor _39835_ (_07414_, _07412_, _06858_);
  not _39836_ (_07415_, _07257_);
  nand _39837_ (_07417_, _07415_, _06909_);
  nor _39838_ (_07418_, _07417_, _07414_);
  nor _39839_ (_28181_, _07418_, rst);
  nand _39840_ (_07420_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  nand _39841_ (_07421_, _04610_, _24789_);
  nand _39842_ (_01092_, _07421_, _07420_);
  nor _39843_ (_07422_, _07179_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _39844_ (_28135_[1], _07422_, rst);
  nor _39845_ (_07423_, _00122_, _25059_);
  nand _39846_ (_07424_, _07423_, _25150_);
  not _39847_ (_07426_, _07423_);
  nand _39848_ (_07428_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nand _39849_ (_01122_, _07428_, _07424_);
  nor _39850_ (_07431_, _06860_, _06849_);
  not _39851_ (_07432_, _07431_);
  nand _39852_ (_07433_, _07432_, _07374_);
  nor _39853_ (_07434_, _06925_, _06860_);
  not _39854_ (_07435_, _07434_);
  nand _39855_ (_07437_, _07435_, _06935_);
  nor _39856_ (_07439_, _07437_, _07433_);
  nor _39857_ (_28135_[2], _07439_, rst);
  nand _39858_ (_07440_, _07423_, _24927_);
  nand _39859_ (_07441_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nand _39860_ (_01139_, _07441_, _07440_);
  nand _39861_ (_07443_, _04251_, _24830_);
  nand _39862_ (_07444_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  nand _39863_ (_01148_, _07444_, _07443_);
  nor _39864_ (_07445_, _06886_, _06860_);
  not _39865_ (_07447_, _07445_);
  nor _39866_ (_07448_, _06860_, _07011_);
  nor _39867_ (_07449_, _07448_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _39868_ (_07450_, _07449_, _07023_);
  not _39869_ (_07451_, _07450_);
  nand _39870_ (_07452_, _07445_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _39871_ (_07453_, _07452_, _07435_);
  nand _39872_ (_07454_, _07414_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _39873_ (_07456_, _07374_, _06852_);
  not _39874_ (_07457_, _07456_);
  nand _39875_ (_07459_, _07457_, _07454_);
  nor _39876_ (_07460_, _07459_, _07453_);
  nand _39877_ (_07461_, _07460_, _07451_);
  nand _39878_ (_07462_, _07461_, _07181_);
  nand _39879_ (_07463_, _07462_, _07447_);
  nor _39880_ (_07464_, _06925_, _06867_);
  nand _39881_ (_07465_, _07461_, _07464_);
  nor _39882_ (_07466_, _07456_, _07414_);
  nand _39883_ (_07467_, _07466_, _07465_);
  nor _39884_ (_07468_, _07467_, _07463_);
  nor _39885_ (_28135_[3], _07468_, rst);
  not _39886_ (_07469_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand _39887_ (_07470_, _07020_, _06864_);
  nor _39888_ (_07471_, _07470_, _07469_);
  nor _39889_ (_07472_, _06907_, _06878_);
  not _39890_ (_07473_, _07472_);
  nand _39891_ (_07474_, _07258_, _07011_);
  nand _39892_ (_07475_, _07474_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand _39893_ (_07476_, _07475_, _07473_);
  nor _39894_ (_07477_, _07476_, _07471_);
  nor _39895_ (_07478_, _07477_, _06859_);
  not _39896_ (_07480_, _07448_);
  nand _39897_ (_07481_, _07100_, _06859_);
  not _39898_ (_07483_, _07481_);
  nor _39899_ (_07485_, _07432_, _07469_);
  nor _39900_ (_07486_, _07485_, _07483_);
  nand _39901_ (_07487_, _07486_, _07480_);
  nor _39902_ (_07488_, _07487_, _07478_);
  nor _39903_ (_28135_[4], _07488_, rst);
  nand _39904_ (_07490_, _03834_, _28096_);
  nand _39905_ (_07491_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nand _39906_ (_01189_, _07491_, _07490_);
  nand _39907_ (_07493_, _01402_, _24830_);
  nand _39908_ (_07494_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  nand _39909_ (_01220_, _07494_, _07493_);
  nand _39910_ (_07496_, _03139_, _24927_);
  nand _39911_ (_07498_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nand _39912_ (_01223_, _07498_, _07496_);
  nand _39913_ (_07499_, _03139_, _25203_);
  nand _39914_ (_07500_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nand _39915_ (_01225_, _07500_, _07499_);
  nand _39916_ (_07501_, _03442_, _28096_);
  nand _39917_ (_07502_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  nand _39918_ (_01227_, _07502_, _07501_);
  nor _39919_ (_07503_, _06886_, _06878_);
  not _39920_ (_07504_, _07503_);
  nand _39921_ (_07505_, _07504_, _06888_);
  nor _39922_ (_07506_, _07472_, _07448_);
  nand _39923_ (_07507_, _07481_, _07506_);
  not _39924_ (_07508_, _07414_);
  nand _39925_ (_07509_, _07508_, _07374_);
  nor _39926_ (_07510_, _07509_, _07507_);
  nand _39927_ (_07511_, _07510_, _07505_);
  nand _39928_ (_07512_, _07511_, _07473_);
  nand _39929_ (_07513_, _07505_, _07373_);
  nand _39930_ (_07514_, _07262_, _06889_);
  nor _39931_ (_07515_, _07447_, _06888_);
  nor _39932_ (_07517_, _07515_, _07434_);
  nand _39933_ (_07518_, _07517_, _07514_);
  nor _39934_ (_07519_, _07518_, _07448_);
  nand _39935_ (_07521_, _07519_, _07513_);
  nor _39936_ (_07522_, _07521_, _07512_);
  nor _39937_ (_28135_[5], _07522_, rst);
  nand _39938_ (_07525_, _03082_, _24927_);
  nand _39939_ (_07526_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nand _39940_ (_01235_, _07526_, _07525_);
  nand _39941_ (_07528_, _03834_, _25039_);
  nand _39942_ (_07529_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nand _39943_ (_01244_, _07529_, _07528_);
  nor _39944_ (_07530_, _04186_, _01605_);
  nand _39945_ (_07531_, _07530_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _39946_ (_07533_, _07531_, _04182_);
  nor _39947_ (_07534_, _07531_, _04182_);
  nor _39948_ (_07535_, _07534_, _01609_);
  nand _39949_ (_07536_, _07535_, _07533_);
  nor _39950_ (_07537_, _04186_, _01597_);
  nor _39951_ (_07538_, _07537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _39952_ (_07539_, _07537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _39953_ (_07540_, _07539_, _01574_);
  nor _39954_ (_07541_, _07540_, _07538_);
  nor _39955_ (_07542_, _04186_, _01632_);
  nor _39956_ (_07544_, _07542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _39957_ (_07546_, _04187_, _01631_);
  nand _39958_ (_07547_, _07546_, _01615_);
  nor _39959_ (_07548_, _07547_, _07544_);
  nor _39960_ (_07549_, _07548_, _07541_);
  nand _39961_ (_07550_, _07549_, _07536_);
  nand _39962_ (_07551_, _07550_, _01642_);
  nand _39963_ (_07552_, _01644_, _25680_);
  nand _39964_ (_07553_, _07552_, _07551_);
  nor _39965_ (_07554_, _07553_, _01573_);
  nand _39966_ (_07555_, _01573_, _04182_);
  nand _39967_ (_07556_, _07555_, _26487_);
  nor _39968_ (_01268_, _07556_, _07554_);
  nor _39969_ (_07557_, _04175_, _25028_);
  not _39970_ (_07558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  not _39971_ (_07559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _39972_ (_07560_, _01587_, _07559_);
  nand _39973_ (_07561_, _07560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _39974_ (_07562_, _07561_, _07558_);
  not _39975_ (_07563_, _07562_);
  nor _39976_ (_07564_, _07563_, _01589_);
  nor _39977_ (_07565_, _07564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _39978_ (_07566_, _07565_, _01595_);
  nand _39979_ (_07567_, _01614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _39980_ (_07568_, _07567_, _04221_);
  nor _39981_ (_07570_, _07568_, _07566_);
  nor _39982_ (_07571_, _07570_, _01644_);
  nor _39983_ (_07572_, _01642_, _01591_);
  nor _39984_ (_07573_, _07572_, _07571_);
  nand _39985_ (_07574_, _07573_, _04175_);
  nand _39986_ (_07575_, _07574_, _26487_);
  nor _39987_ (_01270_, _07575_, _07557_);
  nand _39988_ (_07576_, _07423_, _25039_);
  nand _39989_ (_07577_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  nand _39990_ (_01273_, _07577_, _07576_);
  not _39991_ (_07578_, _07121_);
  nand _39992_ (_07580_, _07470_, _07578_);
  nor _39993_ (_07581_, _07580_, _06928_);
  nor _39994_ (_07582_, _07470_, _06928_);
  not _39995_ (_07584_, _07582_);
  nor _39996_ (_07585_, _07506_, _06928_);
  nor _39997_ (_07587_, _06925_, _06878_);
  not _39998_ (_07589_, _07587_);
  nand _39999_ (_07591_, _07503_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand _40000_ (_07593_, _07591_, _07589_);
  nor _40001_ (_07595_, _07593_, _07585_);
  nand _40002_ (_07596_, _07595_, _07584_);
  nor _40003_ (_07597_, _07596_, _07581_);
  nor _40004_ (_07598_, _07597_, _07374_);
  nor _40005_ (_07600_, _07013_, _07160_);
  nor _40006_ (_07601_, _07597_, _07600_);
  nor _40007_ (_07602_, _07601_, _07503_);
  nand _40008_ (_07603_, _07584_, _07480_);
  nor _40009_ (_07605_, _07603_, _07472_);
  nand _40010_ (_07606_, _07605_, _07602_);
  nor _40011_ (_07607_, _07606_, _07598_);
  nor _40012_ (_28135_[6], _07607_, rst);
  nand _40013_ (_07609_, _28063_, _24927_);
  nand _40014_ (_07610_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nand _40015_ (_01289_, _07610_, _07609_);
  nand _40016_ (_07612_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  nand _40017_ (_07614_, _04610_, _25099_);
  nand _40018_ (_01311_, _07614_, _07612_);
  nor _40019_ (_07616_, _06864_, _06876_);
  nor _40020_ (_07618_, _07480_, _06876_);
  nor _40021_ (_07619_, _07618_, _07472_);
  not _40022_ (_07620_, _07470_);
  nand _40023_ (_07622_, _07620_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _40024_ (_07624_, _07622_, _07619_);
  nor _40025_ (_07625_, _07624_, _07160_);
  nand _40026_ (_07626_, _07625_, _07504_);
  nor _40027_ (_07627_, _07626_, _07616_);
  nor _40028_ (_28135_[7], _07627_, rst);
  nor _40029_ (_07629_, _05824_, _24821_);
  nand _40030_ (_07630_, _05824_, _01608_);
  nand _40031_ (_07632_, _07630_, _26487_);
  nor _40032_ (_01353_, _07632_, _07629_);
  nor _40033_ (_07633_, _04219_, _01574_);
  nor _40034_ (_07634_, _01597_, _01574_);
  nor _40035_ (_07635_, _07634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _40036_ (_07636_, _07635_, _07633_);
  nand _40037_ (_07637_, _04222_, _01614_);
  nor _40038_ (_07638_, _07637_, _04177_);
  nor _40039_ (_07639_, _07638_, _07636_);
  nor _40040_ (_07641_, _07639_, _01644_);
  nor _40041_ (_07643_, _01642_, _01619_);
  nor _40042_ (_07644_, _07643_, _07641_);
  nor _40043_ (_07645_, _07644_, _01573_);
  nor _40044_ (_07646_, _04175_, _26096_);
  nor _40045_ (_07648_, _07646_, _07645_);
  nor _40046_ (_01356_, _07648_, rst);
  nand _40047_ (_07649_, _03082_, _28096_);
  nand _40048_ (_07650_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand _40049_ (_01359_, _07650_, _07649_);
  nand _40050_ (_07651_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  nand _40051_ (_07652_, _01216_, _25150_);
  nand _40052_ (_01365_, _07652_, _07651_);
  nand _40053_ (_07653_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  nand _40054_ (_07654_, _01216_, _24927_);
  nand _40055_ (_01390_, _07654_, _07653_);
  nand _40056_ (_07655_, _07258_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _40057_ (_07656_, _07262_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _40058_ (_07657_, _07656_, _06864_);
  not _40059_ (_07658_, _07015_);
  nand _40060_ (_07659_, _07504_, _07658_);
  nor _40061_ (_07660_, _07659_, _07657_);
  nand _40062_ (_07661_, _07660_, _07655_);
  nor _40063_ (_07662_, _07661_, _07587_);
  nor _40064_ (_28135_[8], _07662_, rst);
  nor _40065_ (_07663_, _05824_, _25028_);
  not _40066_ (_07664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand _40067_ (_07665_, _05824_, _07664_);
  nand _40068_ (_07666_, _07665_, _26487_);
  nor _40069_ (_01412_, _07666_, _07663_);
  nand _40070_ (_07668_, _03834_, _25203_);
  nand _40071_ (_07669_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nand _40072_ (_01417_, _07669_, _07668_);
  nor _40073_ (_07670_, _28104_, _25057_);
  nand _40074_ (_07672_, _07670_, _24789_);
  not _40075_ (_07674_, _07670_);
  nand _40076_ (_07675_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  nand _40077_ (_01442_, _07675_, _07672_);
  nand _40078_ (_07677_, _03704_, _24830_);
  nand _40079_ (_07679_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nand _40080_ (_01446_, _07679_, _07677_);
  nand _40081_ (_07682_, _03571_, _24927_);
  nand _40082_ (_07683_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  nand _40083_ (_01449_, _07683_, _07682_);
  nand _40084_ (_07685_, _03571_, _25099_);
  nand _40085_ (_07686_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  nand _40086_ (_01451_, _07686_, _07685_);
  nand _40087_ (_07689_, _03561_, _25150_);
  nand _40088_ (_07691_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  nand _40089_ (_01455_, _07691_, _07689_);
  nand _40090_ (_07692_, _03561_, _25099_);
  nand _40091_ (_07693_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nand _40092_ (_01458_, _07693_, _07692_);
  nand _40093_ (_07696_, _03540_, _25150_);
  nand _40094_ (_07698_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nand _40095_ (_01466_, _07698_, _07696_);
  nand _40096_ (_07699_, _03540_, _28096_);
  nand _40097_ (_07700_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nand _40098_ (_01469_, _07700_, _07699_);
  nand _40099_ (_07702_, _01178_, _25039_);
  nand _40100_ (_07704_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand _40101_ (_01472_, _07704_, _07702_);
  nand _40102_ (_07706_, _03520_, _28096_);
  nand _40103_ (_07708_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nand _40104_ (_01478_, _07708_, _07706_);
  nor _40105_ (_07709_, _06886_, _06855_);
  nor _40106_ (_07710_, _07709_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _40107_ (_07711_, _07710_, _06864_);
  nor _40108_ (_07712_, _07507_, _07503_);
  nor _40109_ (_07713_, _07712_, _06895_);
  nor _40110_ (_07714_, _07412_, _06864_);
  not _40111_ (_07716_, _07714_);
  nor _40112_ (_07717_, _07508_, _06895_);
  nor _40113_ (_07718_, _07717_, _07587_);
  nand _40114_ (_07719_, _07718_, _07716_);
  nor _40115_ (_07721_, _07719_, _07713_);
  nand _40116_ (_07722_, _07721_, _07658_);
  nor _40117_ (_07724_, _07722_, _07711_);
  nor _40118_ (_28135_[9], _07724_, rst);
  nand _40119_ (_07725_, _03446_, _24789_);
  nand _40120_ (_07726_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand _40121_ (_01487_, _07726_, _07725_);
  nor _40122_ (_07727_, _04173_, _24920_);
  nor _40123_ (_07728_, _04188_, _01634_);
  nand _40124_ (_07730_, _07728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _40125_ (_07732_, _07730_, _04176_);
  nor _40126_ (_07733_, _07732_, _01616_);
  nor _40127_ (_07734_, _04191_, _01597_);
  not _40128_ (_07736_, _07734_);
  nor _40129_ (_07738_, _07736_, _04176_);
  nor _40130_ (_07739_, _07738_, _04208_);
  nor _40131_ (_07740_, _07739_, _07733_);
  nor _40132_ (_07741_, _07740_, _04177_);
  nand _40133_ (_07742_, _04187_, _01604_);
  nor _40134_ (_07743_, _07742_, _04181_);
  nand _40135_ (_07744_, _07743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _40136_ (_07746_, _07744_, _04177_);
  not _40137_ (_07747_, _01611_);
  nor _40138_ (_07748_, _04194_, _07747_);
  nand _40139_ (_07749_, _07748_, _07746_);
  nand _40140_ (_07750_, _07732_, _01617_);
  nand _40141_ (_07751_, _07738_, _01574_);
  nand _40142_ (_07752_, _07751_, _07750_);
  nand _40143_ (_07753_, _07752_, _04177_);
  nand _40144_ (_07754_, _07753_, _07749_);
  nor _40145_ (_07755_, _07754_, _07741_);
  nand _40146_ (_07756_, _07755_, _04173_);
  nand _40147_ (_07757_, _07756_, _04175_);
  nor _40148_ (_07758_, _07757_, _07727_);
  nor _40149_ (_07760_, _04175_, _04177_);
  nor _40150_ (_07761_, _07760_, _07758_);
  nor _40151_ (_01495_, _07761_, rst);
  nand _40152_ (_07762_, _03446_, _25203_);
  nand _40153_ (_07763_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nand _40154_ (_01505_, _07763_, _07762_);
  nand _40155_ (_07764_, _25160_, _24927_);
  nand _40156_ (_07765_, _25162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand _40157_ (_01510_, _07765_, _07764_);
  nor _40158_ (_07766_, _07166_, _06858_);
  not _40159_ (_07767_, _07766_);
  nor _40160_ (_07768_, _07767_, _06932_);
  nand _40161_ (_07769_, _07432_, _07589_);
  nand _40162_ (_07771_, _07769_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _40163_ (_07773_, _07771_);
  nor _40164_ (_07774_, _07773_, _07768_);
  not _40165_ (_07775_, _07774_);
  nor _40166_ (_07776_, _07775_, _07015_);
  nor _40167_ (_07777_, _07172_, _07464_);
  nand _40168_ (_07778_, _07777_, _07374_);
  nand _40169_ (_07779_, _07714_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _40170_ (_07780_, _07015_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _40171_ (_07781_, _07780_, _07779_);
  nor _40172_ (_07782_, _06925_, _06873_);
  not _40173_ (_07783_, _07782_);
  nor _40174_ (_07785_, _06855_, _06845_);
  nor _40175_ (_07787_, _07785_, _06932_);
  nand _40176_ (_07789_, _07787_, _06858_);
  nand _40177_ (_07790_, _07789_, _07783_);
  nor _40178_ (_07791_, _07790_, _07781_);
  nand _40179_ (_07793_, _07791_, _07774_);
  nand _40180_ (_07794_, _07793_, _07778_);
  nand _40181_ (_07795_, _07794_, _07776_);
  nor _40182_ (_07796_, _06886_, _06873_);
  not _40183_ (_07797_, _07796_);
  nand _40184_ (_07798_, _07797_, _07716_);
  nor _40185_ (_07799_, _07798_, _07795_);
  nor _40186_ (_28135_[10], _07799_, rst);
  nand _40187_ (_07800_, _03139_, _24789_);
  nand _40188_ (_07801_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand _40189_ (_01576_, _07801_, _07800_);
  nand _40190_ (_07802_, _03082_, _24789_);
  nand _40191_ (_07803_, _03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand _40192_ (_01579_, _07803_, _07802_);
  nand _40193_ (_07804_, _03782_, _24789_);
  nand _40194_ (_07805_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  nand _40195_ (_01581_, _07805_, _07804_);
  nand _40196_ (_07806_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  nand _40197_ (_07807_, _04610_, _24830_);
  nand _40198_ (_01583_, _07807_, _07806_);
  nand _40199_ (_07808_, _03782_, _24830_);
  nand _40200_ (_07809_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  nand _40201_ (_01586_, _07809_, _07808_);
  nor _40202_ (_07810_, _28104_, _24999_);
  nand _40203_ (_07811_, _07810_, _25099_);
  not _40204_ (_07812_, _07810_);
  nand _40205_ (_07813_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nand _40206_ (_01596_, _07813_, _07811_);
  not _40207_ (_07814_, _24989_);
  nor _40208_ (_07816_, _07814_, _24069_);
  nand _40209_ (_07818_, _25156_, _07816_);
  nor _40210_ (_07819_, _07818_, _25057_);
  nand _40211_ (_07821_, _07819_, _25203_);
  not _40212_ (_07823_, _07819_);
  nand _40213_ (_07824_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  nand _40214_ (_01600_, _07824_, _07821_);
  nand _40215_ (_07825_, _03520_, _25150_);
  nand _40216_ (_07826_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nand _40217_ (_01610_, _07826_, _07825_);
  nand _40218_ (_07827_, _01398_, _24830_);
  nand _40219_ (_07828_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nand _40220_ (_01623_, _07828_, _07827_);
  nand _40221_ (_07829_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  nand _40222_ (_07830_, _04015_, _25203_);
  nand _40223_ (_01629_, _07830_, _07829_);
  not _40224_ (_07831_, _07032_);
  nor _40225_ (_07832_, _06873_, _07011_);
  nor _40226_ (_07833_, _07832_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _40227_ (_07834_, _07833_, _07831_);
  nor _40228_ (_07835_, _07658_, _06871_);
  nor _40229_ (_07836_, _07835_, _07782_);
  nor _40230_ (_07838_, _07797_, _06871_);
  nor _40231_ (_07839_, _07578_, _06871_);
  nor _40232_ (_07840_, _07839_, _07838_);
  nand _40233_ (_07841_, _07840_, _07836_);
  nor _40234_ (_07843_, _07841_, _07834_);
  nor _40235_ (_07844_, _07843_, _07777_);
  nor _40236_ (_07846_, _07833_, _07374_);
  nor _40237_ (_07848_, _07835_, _07714_);
  nor _40238_ (_07849_, _07481_, _06871_);
  nand _40239_ (_07850_, _07414_, \oc8051_symbolic_cxrom1.regvalid [11]);
  not _40240_ (_07851_, _07839_);
  nand _40241_ (_07852_, _07851_, _07850_);
  nor _40242_ (_07853_, _07852_, _07849_);
  nand _40243_ (_07854_, _07853_, _07848_);
  nor _40244_ (_07855_, _07854_, _07846_);
  nand _40245_ (_07856_, _07855_, _07797_);
  nor _40246_ (_07857_, _07856_, _07844_);
  nor _40247_ (_28135_[11], _07857_, rst);
  nand _40248_ (_07858_, _07423_, _24789_);
  nand _40249_ (_07859_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  nand _40250_ (_01656_, _07859_, _07858_);
  nand _40251_ (_07860_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  nand _40252_ (_07861_, _01216_, _24789_);
  nand _40253_ (_01679_, _07861_, _07860_);
  nand _40254_ (_07862_, _00619_, _23958_);
  nand _40255_ (_07863_, _07862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nand _40256_ (_07864_, _07863_, _00622_);
  not _40257_ (_07865_, _03408_);
  not _40258_ (_07866_, _04721_);
  nand _40259_ (_07867_, _23958_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _40260_ (_07868_, _07867_, _26133_);
  nor _40261_ (_07869_, _07868_, _07866_);
  nor _40262_ (_07870_, _07869_, _07865_);
  nor _40263_ (_07871_, _07870_, _07864_);
  nor _40264_ (_07872_, _00235_, _25627_);
  nand _40265_ (_07873_, _07872_, _25140_);
  nand _40266_ (_07874_, _07873_, _26487_);
  nor _40267_ (_01698_, _07874_, _07871_);
  nand _40268_ (_07875_, _00494_, _26135_);
  nor _40269_ (_07876_, _07875_, _24716_);
  nand _40270_ (_07877_, _07875_, _00543_);
  nand _40271_ (_07878_, _07877_, _00503_);
  nor _40272_ (_07879_, _07878_, _07876_);
  nor _40273_ (_07880_, _00503_, _25625_);
  nor _40274_ (_07881_, _07880_, _07879_);
  nor _40275_ (_01703_, _07881_, rst);
  nor _40276_ (_07882_, _25059_, _25047_);
  nand _40277_ (_07883_, _07882_, _24789_);
  not _40278_ (_07884_, _07882_);
  nand _40279_ (_07885_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  nand _40280_ (_01708_, _07885_, _07883_);
  not _40281_ (_07886_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _40282_ (_07887_, _07415_, _07886_);
  nand _40283_ (_07888_, _06849_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _40284_ (_07889_, _07888_, _06860_);
  nand _40285_ (_07890_, _07445_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand _40286_ (_07891_, _07890_, _07797_);
  nor _40287_ (_07892_, _07891_, _07889_);
  nor _40288_ (_07893_, _06886_, _06867_);
  nor _40289_ (_07894_, _07893_, _07357_);
  nor _40290_ (_07895_, _07262_, _06877_);
  nor _40291_ (_07896_, _07895_, _07886_);
  nor _40292_ (_07897_, _07896_, _07894_);
  nand _40293_ (_07898_, _07897_, _07892_);
  nor _40294_ (_07899_, _07898_, _07887_);
  nor _40295_ (_28135_[12], _07899_, rst);
  nand _40296_ (_07900_, _07882_, _25150_);
  nand _40297_ (_07901_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  nand _40298_ (_01721_, _07901_, _07900_);
  nand _40299_ (_07902_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  nand _40300_ (_07903_, _04601_, _28096_);
  nand _40301_ (_01727_, _07903_, _07902_);
  nand _40302_ (_07904_, _04308_, _24830_);
  nand _40303_ (_07905_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nand _40304_ (_01736_, _07905_, _07904_);
  nand _40305_ (_07906_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  nand _40306_ (_07907_, _04264_, _25039_);
  nand _40307_ (_01744_, _07907_, _07906_);
  nor _40308_ (_07908_, _00631_, _28080_);
  nand _40309_ (_07909_, _07908_, _24789_);
  not _40310_ (_07910_, _07908_);
  nand _40311_ (_07911_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  nand _40312_ (_01755_, _07911_, _07909_);
  nor _40313_ (_07912_, _06849_, _06891_);
  nor _40314_ (_07913_, _07912_, _07164_);
  nor _40315_ (_07914_, _07913_, _06859_);
  nor _40316_ (_07915_, _07914_, _06865_);
  nor _40317_ (_07916_, _07915_, _07257_);
  nand _40318_ (_07917_, _06959_, _06892_);
  nand _40319_ (_07918_, _06864_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _40320_ (_07919_, _07918_, _06969_);
  nor _40321_ (_07920_, _07919_, _07893_);
  nand _40322_ (_07921_, _07920_, _07917_);
  nor _40323_ (_07922_, _07921_, _07916_);
  nor _40324_ (_28135_[13], _07922_, rst);
  nand _40325_ (_07923_, _01153_, _28096_);
  nand _40326_ (_07924_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nand _40327_ (_01784_, _07924_, _07923_);
  nand _40328_ (_07925_, _07882_, _24927_);
  nand _40329_ (_07926_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  nand _40330_ (_01798_, _07926_, _07925_);
  nand _40331_ (_07927_, _03704_, _25099_);
  nand _40332_ (_07928_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  nand _40333_ (_01802_, _07928_, _07927_);
  nand _40334_ (_07929_, _03561_, _28096_);
  nand _40335_ (_07930_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nand _40336_ (_01805_, _07930_, _07929_);
  nand _40337_ (_07931_, _01178_, _24927_);
  nand _40338_ (_07932_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand _40339_ (_01807_, _07932_, _07931_);
  nand _40340_ (_07933_, _07810_, _24830_);
  nand _40341_ (_07934_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  nand _40342_ (_01817_, _07934_, _07933_);
  nand _40343_ (_07935_, _07819_, _24830_);
  nand _40344_ (_07936_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  nand _40345_ (_01821_, _07936_, _07935_);
  not _40346_ (_07937_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nand _40347_ (_07938_, _06865_, _07011_);
  nand _40348_ (_07939_, _07938_, _07937_);
  nor _40349_ (_07940_, _07939_, _07832_);
  nor _40350_ (_28135_[14], _07940_, rst);
  nor _40351_ (_07941_, _00267_, _25627_);
  not _40352_ (_07942_, _07941_);
  nor _40353_ (_07943_, _07942_, _24782_);
  not _40354_ (_07944_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _40355_ (_07945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _05826_);
  nor _40356_ (_07946_, _07664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _40357_ (_07947_, _07946_, _07945_);
  nor _40358_ (_07948_, _00139_, _25627_);
  nor _40359_ (_07949_, _07948_, _07947_);
  nor _40360_ (_07950_, _07949_, _07944_);
  not _40361_ (_07951_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  not _40362_ (_07952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not _40363_ (_07953_, t1_i);
  nand _40364_ (_07954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _07953_);
  nand _40365_ (_07955_, _07954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nor _40366_ (_07956_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _01603_);
  not _40367_ (_07957_, _07956_);
  nor _40368_ (_07958_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nor _40369_ (_07959_, _07958_, _07957_);
  nand _40370_ (_07960_, _07959_, _07955_);
  not _40371_ (_07961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _40372_ (_07962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand _40373_ (_07963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _40374_ (_07964_, _07963_, _07962_);
  not _40375_ (_07965_, _07964_);
  nor _40376_ (_07966_, _07965_, _07961_);
  not _40377_ (_07967_, _07966_);
  nor _40378_ (_07968_, _07967_, _07960_);
  not _40379_ (_07969_, _07968_);
  nor _40380_ (_07970_, _07969_, _07952_);
  not _40381_ (_07971_, _07970_);
  nor _40382_ (_07972_, _07971_, _07951_);
  nor _40383_ (_07973_, _07972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _40384_ (_07974_, _07965_, _07960_);
  not _40385_ (_07975_, _07974_);
  nor _40386_ (_07976_, _07975_, _07961_);
  not _40387_ (_07977_, _07976_);
  nor _40388_ (_07978_, _07952_, _07944_);
  nand _40389_ (_07979_, _07978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _40390_ (_07980_, _07979_, _07977_);
  nor _40391_ (_07981_, _07980_, _07973_);
  nand _40392_ (_07982_, _07981_, _07949_);
  not _40393_ (_07983_, _07948_);
  not _40394_ (_07984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not _40395_ (_07985_, _07972_);
  nor _40396_ (_07986_, _07985_, _07944_);
  nand _40397_ (_07987_, _07986_, _07945_);
  nor _40398_ (_07988_, _07987_, _07984_);
  nand _40399_ (_07989_, _07988_, _07983_);
  nand _40400_ (_07990_, _07989_, _07982_);
  nor _40401_ (_07991_, _07990_, _07950_);
  nand _40402_ (_07992_, _07942_, _07991_);
  nand _40403_ (_07993_, _07992_, _26487_);
  nor _40404_ (_01847_, _07993_, _07943_);
  nor _40405_ (_07994_, _01604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nand _40406_ (_07995_, _01611_, _26487_);
  nor _40407_ (_07996_, _07995_, _07994_);
  nand _40408_ (_07997_, _07996_, _04173_);
  not _40409_ (_07998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _40410_ (_07999_, _04232_, _07998_);
  not _40411_ (_08000_, _07999_);
  nand _40412_ (_08001_, _08000_, _01604_);
  nand _40413_ (_08002_, _08001_, _04175_);
  nor _40414_ (_01872_, _08002_, _07997_);
  nand _40415_ (_08003_, _24927_, _24852_);
  nand _40416_ (_08004_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nand _40417_ (_01876_, _08004_, _08003_);
  nand _40418_ (_08005_, _07423_, _28096_);
  nand _40419_ (_08006_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  nand _40420_ (_01886_, _08006_, _08005_);
  nor _40421_ (_08007_, _03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _40422_ (_01891_, _08007_, _04336_);
  nand _40423_ (_08008_, _07423_, _25099_);
  nand _40424_ (_08009_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nand _40425_ (_01897_, _08009_, _08008_);
  nor _40426_ (_08010_, _06865_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _40427_ (_28135_[15], _08010_, rst);
  nor _40428_ (_08011_, _07393_, _07264_);
  nor _40429_ (_08012_, _08011_, _07394_);
  not _40430_ (_08013_, _08012_);
  nor _40431_ (_08014_, _08013_, _06886_);
  nand _40432_ (_08015_, _08014_, _07392_);
  not _40433_ (_08016_, _08015_);
  not _40434_ (_08017_, _07464_);
  nor _40435_ (_08018_, _07361_, _08017_);
  nor _40436_ (_08019_, _07367_, _07374_);
  not _40437_ (_08020_, _08019_);
  nor _40438_ (_08021_, _07376_, _07508_);
  nor _40439_ (_08022_, _08021_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  not _40440_ (_08023_, _08021_);
  nor _40441_ (_08024_, _08023_, word_in[0]);
  nor _40442_ (_08025_, _08024_, _08022_);
  nand _40443_ (_08026_, _08025_, _08020_);
  not _40444_ (_08027_, word_in[8]);
  nor _40445_ (_08028_, _07367_, _08027_);
  nand _40446_ (_08029_, _08028_, _08019_);
  nand _40447_ (_08030_, _08029_, _08026_);
  nor _40448_ (_08031_, _08030_, _08018_);
  not _40449_ (_08032_, _08018_);
  nor _40450_ (_08033_, _08032_, word_in[16]);
  nor _40451_ (_08034_, _08033_, _08031_);
  nor _40452_ (_08035_, _08034_, _08016_);
  nor _40453_ (_08036_, _08015_, word_in[24]);
  nor _40454_ (_28169_[0], _08036_, _08035_);
  nand _40455_ (_08037_, _07354_, word_in[25]);
  nor _40456_ (_08038_, _08037_, rst);
  nand _40457_ (_08039_, _08038_, _08014_);
  not _40458_ (_08040_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nand _40459_ (_08041_, _08023_, _08040_);
  not _40460_ (_08042_, word_in[1]);
  nand _40461_ (_08043_, _08021_, _08042_);
  nand _40462_ (_08044_, _08043_, _08041_);
  nand _40463_ (_08045_, _08044_, _08020_);
  not _40464_ (_08046_, word_in[9]);
  nand _40465_ (_08047_, _08019_, _08046_);
  nand _40466_ (_08048_, _08047_, _08045_);
  nand _40467_ (_08049_, _08048_, _08032_);
  nor _40468_ (_08050_, _08032_, word_in[17]);
  nor _40469_ (_08051_, _08050_, _08016_);
  nand _40470_ (_08052_, _08051_, _08049_);
  nand _40471_ (_28169_[1], _08052_, _08039_);
  nand _40472_ (_08053_, _07354_, word_in[26]);
  nor _40473_ (_08054_, _08053_, rst);
  nand _40474_ (_08055_, _08054_, _08014_);
  not _40475_ (_08056_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand _40476_ (_08058_, _08023_, _08056_);
  not _40477_ (_08059_, word_in[2]);
  nand _40478_ (_08061_, _08021_, _08059_);
  nand _40479_ (_08062_, _08061_, _08058_);
  nand _40480_ (_08063_, _08062_, _08020_);
  not _40481_ (_08064_, word_in[10]);
  nand _40482_ (_08065_, _08019_, _08064_);
  nand _40483_ (_08066_, _08065_, _08063_);
  nand _40484_ (_08067_, _08066_, _08032_);
  nor _40485_ (_08068_, _08032_, word_in[18]);
  nor _40486_ (_08069_, _08068_, _08016_);
  nand _40487_ (_08070_, _08069_, _08067_);
  nand _40488_ (_28169_[2], _08070_, _08055_);
  nor _40489_ (_08071_, _08021_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _40490_ (_08072_, _08023_, word_in[3]);
  nor _40491_ (_08073_, _08072_, _08071_);
  nor _40492_ (_08075_, _08073_, _08019_);
  nor _40493_ (_08076_, _08020_, word_in[11]);
  nor _40494_ (_08077_, _08076_, _08075_);
  nor _40495_ (_08078_, _08077_, _08018_);
  nor _40496_ (_08079_, _08032_, word_in[19]);
  nor _40497_ (_08080_, _08079_, _08078_);
  nor _40498_ (_08081_, _08080_, _08016_);
  nor _40499_ (_08082_, _08015_, word_in[27]);
  nor _40500_ (_28169_[3], _08082_, _08081_);
  nand _40501_ (_08083_, _07354_, word_in[28]);
  nor _40502_ (_08084_, _08083_, rst);
  nand _40503_ (_08085_, _08084_, _08014_);
  not _40504_ (_08086_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nand _40505_ (_08087_, _08023_, _08086_);
  not _40506_ (_08088_, word_in[4]);
  nand _40507_ (_08089_, _08021_, _08088_);
  nand _40508_ (_08090_, _08089_, _08087_);
  nand _40509_ (_08091_, _08090_, _08020_);
  not _40510_ (_08092_, word_in[12]);
  nand _40511_ (_08094_, _08019_, _08092_);
  nand _40512_ (_08095_, _08094_, _08091_);
  nand _40513_ (_08096_, _08095_, _08032_);
  nor _40514_ (_08097_, _08032_, word_in[20]);
  nor _40515_ (_08099_, _08097_, _08016_);
  nand _40516_ (_08100_, _08099_, _08096_);
  nand _40517_ (_28169_[4], _08100_, _08085_);
  nand _40518_ (_08101_, _07354_, word_in[29]);
  nor _40519_ (_08102_, _08101_, rst);
  nand _40520_ (_08103_, _08102_, _08014_);
  not _40521_ (_08104_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nand _40522_ (_08105_, _08023_, _08104_);
  not _40523_ (_08106_, word_in[5]);
  nand _40524_ (_08107_, _08021_, _08106_);
  nand _40525_ (_08108_, _08107_, _08105_);
  nand _40526_ (_08109_, _08108_, _08020_);
  not _40527_ (_08110_, word_in[13]);
  nand _40528_ (_08111_, _08019_, _08110_);
  nand _40529_ (_08112_, _08111_, _08109_);
  nand _40530_ (_08113_, _08112_, _08032_);
  nor _40531_ (_08114_, _08032_, word_in[21]);
  nor _40532_ (_08115_, _08114_, _08016_);
  nand _40533_ (_08116_, _08115_, _08113_);
  nand _40534_ (_28169_[5], _08116_, _08103_);
  nor _40535_ (_08117_, _08021_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _40536_ (_08118_, _08023_, word_in[6]);
  nor _40537_ (_08119_, _08118_, _08117_);
  nor _40538_ (_08120_, _08119_, _08019_);
  nor _40539_ (_08121_, _08020_, word_in[14]);
  nor _40540_ (_08122_, _08121_, _08120_);
  nor _40541_ (_08123_, _08122_, _08018_);
  nor _40542_ (_08124_, _08032_, word_in[22]);
  nor _40543_ (_08125_, _08124_, _08123_);
  nor _40544_ (_08126_, _08125_, _08016_);
  nor _40545_ (_08127_, _08015_, word_in[30]);
  nor _40546_ (_28169_[6], _08127_, _08126_);
  nand _40547_ (_08128_, _08014_, _07408_);
  not _40548_ (_08129_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _40549_ (_08130_, _08023_, _08129_);
  nand _40550_ (_08131_, _08021_, _07381_);
  nand _40551_ (_08132_, _08131_, _08130_);
  nand _40552_ (_08133_, _08132_, _08020_);
  nand _40553_ (_08134_, _08019_, _07387_);
  nand _40554_ (_08135_, _08134_, _08133_);
  nand _40555_ (_08136_, _08135_, _08032_);
  nor _40556_ (_08137_, _08032_, word_in[23]);
  nor _40557_ (_08138_, _08137_, _08016_);
  nand _40558_ (_08139_, _08138_, _08136_);
  nand _40559_ (_28169_[7], _08139_, _08128_);
  nor _40560_ (_08141_, _25049_, _24884_);
  not _40561_ (_08142_, _08141_);
  nor _40562_ (_08144_, _08142_, _24795_);
  not _40563_ (_08146_, _08144_);
  nand _40564_ (_08147_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  nand _40565_ (_08148_, _08144_, _25203_);
  nand _40566_ (_02121_, _08148_, _08147_);
  nor _40567_ (_08149_, _08142_, _24978_);
  not _40568_ (_08150_, _08149_);
  nand _40569_ (_08151_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  nand _40570_ (_08152_, _08149_, _24789_);
  nand _40571_ (_02126_, _08152_, _08151_);
  nor _40572_ (_08153_, _08142_, _24999_);
  not _40573_ (_08154_, _08153_);
  nand _40574_ (_08156_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  nand _40575_ (_08157_, _08153_, _25099_);
  nand _40576_ (_02140_, _08157_, _08156_);
  nor _40577_ (_08158_, _08142_, _25057_);
  not _40578_ (_08159_, _08158_);
  nand _40579_ (_08160_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nand _40580_ (_08161_, _08158_, _28096_);
  nand _40581_ (_02144_, _08161_, _08160_);
  nor _40582_ (_08163_, _08142_, _28080_);
  not _40583_ (_08164_, _08163_);
  nand _40584_ (_08165_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  nand _40585_ (_08166_, _08163_, _25203_);
  nand _40586_ (_02148_, _08166_, _08165_);
  nor _40587_ (_08167_, _08142_, _25047_);
  not _40588_ (_08168_, _08167_);
  nand _40589_ (_08170_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nand _40590_ (_08171_, _08167_, _25099_);
  nand _40591_ (_02157_, _08171_, _08170_);
  nor _40592_ (_08172_, _07393_, _06925_);
  nand _40593_ (_08173_, _08172_, _08012_);
  nor _40594_ (_08174_, _07361_, _07011_);
  not _40595_ (_08175_, _08174_);
  nor _40596_ (_08176_, _08175_, _07181_);
  not _40597_ (_08177_, _08176_);
  nor _40598_ (_08178_, _07367_, _06907_);
  not _40599_ (_08179_, _08178_);
  nor _40600_ (_08180_, _08179_, _07025_);
  not _40601_ (_08181_, _08180_);
  not _40602_ (_08182_, word_in[0]);
  nor _40603_ (_08183_, _07376_, _08182_);
  nand _40604_ (_08184_, _08183_, _07445_);
  nor _40605_ (_08185_, _07376_, _07447_);
  not _40606_ (_08186_, _08185_);
  nand _40607_ (_08187_, _08186_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _40608_ (_08188_, _08187_, _08184_);
  nand _40609_ (_08189_, _08188_, _08181_);
  nand _40610_ (_08190_, _08180_, word_in[8]);
  nand _40611_ (_08191_, _08190_, _08189_);
  nand _40612_ (_08192_, _08191_, _08177_);
  nand _40613_ (_08193_, _08176_, word_in[16]);
  nand _40614_ (_08194_, _08193_, _08192_);
  nand _40615_ (_08195_, _08194_, _08173_);
  not _40616_ (_08196_, _08173_);
  nand _40617_ (_08197_, _08196_, word_in[24]);
  nand _40618_ (_28174_[0], _08197_, _08195_);
  not _40619_ (_08198_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _40620_ (_08199_, _08185_, _08198_);
  nor _40621_ (_08200_, _07376_, _08042_);
  not _40622_ (_08201_, _08200_);
  nor _40623_ (_08202_, _08201_, _07447_);
  nor _40624_ (_08203_, _08202_, _08199_);
  nor _40625_ (_08204_, _08203_, _08180_);
  nor _40626_ (_08205_, _08181_, _08046_);
  nor _40627_ (_08206_, _08205_, _08204_);
  nor _40628_ (_08207_, _08206_, _08176_);
  nand _40629_ (_08208_, _08176_, word_in[17]);
  nand _40630_ (_08209_, _08208_, _08173_);
  nor _40631_ (_08210_, _08209_, _08207_);
  nor _40632_ (_08211_, _08173_, _08038_);
  nor _40633_ (_28174_[1], _08211_, _08210_);
  nor _40634_ (_08212_, _08142_, _00954_);
  not _40635_ (_08213_, _08212_);
  nand _40636_ (_08214_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  nand _40637_ (_08215_, _08212_, _25203_);
  nand _40638_ (_02171_, _08215_, _08214_);
  not _40639_ (_08216_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _40640_ (_08217_, _08185_, _08216_);
  nor _40641_ (_08218_, _07376_, _08059_);
  not _40642_ (_08219_, _08218_);
  nor _40643_ (_08220_, _08219_, _07447_);
  nor _40644_ (_08221_, _08220_, _08217_);
  nor _40645_ (_08222_, _08221_, _08180_);
  nor _40646_ (_08223_, _08181_, _08064_);
  nor _40647_ (_08224_, _08223_, _08222_);
  nor _40648_ (_08225_, _08224_, _08176_);
  nand _40649_ (_08226_, _08176_, word_in[18]);
  nand _40650_ (_08227_, _08226_, _08173_);
  nor _40651_ (_08228_, _08227_, _08225_);
  nor _40652_ (_08229_, _08173_, _08054_);
  nor _40653_ (_28174_[2], _08229_, _08228_);
  nor _40654_ (_08230_, _08142_, _00393_);
  not _40655_ (_08231_, _08230_);
  nand _40656_ (_08232_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nand _40657_ (_08233_, _08230_, _25150_);
  nand _40658_ (_02175_, _08233_, _08232_);
  nand _40659_ (_08234_, _07354_, word_in[27]);
  nor _40660_ (_08235_, _08234_, rst);
  nand _40661_ (_08236_, _08196_, _08235_);
  not _40662_ (_08237_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _40663_ (_08238_, _08185_, _08237_);
  nand _40664_ (_08239_, _07375_, word_in[3]);
  nor _40665_ (_08240_, _08239_, _07447_);
  nor _40666_ (_08241_, _08240_, _08238_);
  nor _40667_ (_08242_, _08241_, _08180_);
  not _40668_ (_08243_, word_in[11]);
  nor _40669_ (_08244_, _08181_, _08243_);
  nor _40670_ (_08245_, _08244_, _08242_);
  nand _40671_ (_08246_, _08245_, _08177_);
  nand _40672_ (_08247_, _07227_, word_in[19]);
  nor _40673_ (_08248_, _08247_, rst);
  nor _40674_ (_08249_, _08177_, _08248_);
  nor _40675_ (_08250_, _08249_, _08196_);
  nand _40676_ (_08251_, _08250_, _08246_);
  nand _40677_ (_28174_[3], _08251_, _08236_);
  nand _40678_ (_08252_, _08196_, _08084_);
  nand _40679_ (_08253_, _08186_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _40680_ (_08254_, _07376_, _08088_);
  nand _40681_ (_08255_, _08254_, _07445_);
  nand _40682_ (_08256_, _08255_, _08253_);
  nand _40683_ (_08257_, _08256_, _08181_);
  nand _40684_ (_08258_, _08180_, word_in[12]);
  nand _40685_ (_08259_, _08258_, _08257_);
  nand _40686_ (_08260_, _08259_, _08177_);
  nand _40687_ (_08261_, _08176_, word_in[20]);
  nand _40688_ (_08262_, _08261_, _08260_);
  nand _40689_ (_08263_, _08262_, _08173_);
  nand _40690_ (_28174_[4], _08263_, _08252_);
  nor _40691_ (_08264_, _08142_, _24882_);
  not _40692_ (_08265_, _08264_);
  nand _40693_ (_08266_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  nand _40694_ (_08267_, _08264_, _25039_);
  nand _40695_ (_02180_, _08267_, _08266_);
  not _40696_ (_08269_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _40697_ (_08270_, _08185_, _08269_);
  nand _40698_ (_08271_, _07375_, word_in[5]);
  nor _40699_ (_08272_, _08271_, _07447_);
  nor _40700_ (_08273_, _08272_, _08270_);
  nor _40701_ (_08274_, _08273_, _08180_);
  nor _40702_ (_08275_, _08181_, _08110_);
  nor _40703_ (_08276_, _08275_, _08274_);
  nor _40704_ (_08277_, _08276_, _08176_);
  nand _40705_ (_08278_, _08176_, word_in[21]);
  nand _40706_ (_08279_, _08278_, _08173_);
  nor _40707_ (_08280_, _08279_, _08277_);
  nor _40708_ (_08281_, _08173_, _08102_);
  nor _40709_ (_28174_[5], _08281_, _08280_);
  nand _40710_ (_08282_, _07354_, word_in[30]);
  nor _40711_ (_08283_, _08282_, rst);
  nand _40712_ (_08284_, _08196_, _08283_);
  not _40713_ (_08285_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _40714_ (_08286_, _08185_, _08285_);
  nand _40715_ (_08287_, _07375_, word_in[6]);
  nor _40716_ (_08289_, _08287_, _07447_);
  nor _40717_ (_08290_, _08289_, _08286_);
  nor _40718_ (_08291_, _08290_, _08180_);
  not _40719_ (_08293_, word_in[14]);
  nor _40720_ (_08294_, _08181_, _08293_);
  nor _40721_ (_08295_, _08294_, _08291_);
  nand _40722_ (_08296_, _08295_, _08177_);
  nand _40723_ (_08297_, _07227_, word_in[22]);
  nor _40724_ (_08298_, _08297_, rst);
  nor _40725_ (_08299_, _08177_, _08298_);
  nor _40726_ (_08300_, _08299_, _08196_);
  nand _40727_ (_08301_, _08300_, _08296_);
  nand _40728_ (_28174_[6], _08301_, _08284_);
  nand _40729_ (_08302_, _08196_, _07408_);
  not _40730_ (_08304_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _40731_ (_08305_, _08185_, _08304_);
  nor _40732_ (_08306_, _07376_, _07381_);
  not _40733_ (_08307_, _08306_);
  nor _40734_ (_08308_, _08307_, _07447_);
  nor _40735_ (_08309_, _08308_, _08305_);
  nor _40736_ (_08310_, _08309_, _08180_);
  nor _40737_ (_08311_, _08181_, _07387_);
  nor _40738_ (_08312_, _08311_, _08310_);
  nand _40739_ (_08313_, _08312_, _08177_);
  nor _40740_ (_08314_, _08177_, _07400_);
  nor _40741_ (_08315_, _08314_, _08196_);
  nand _40742_ (_08317_, _08315_, _08313_);
  nand _40743_ (_28174_[7], _08317_, _08302_);
  nor _40744_ (_08319_, _08142_, _00114_);
  not _40745_ (_08320_, _08319_);
  nand _40746_ (_08321_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  nand _40747_ (_08323_, _08319_, _24927_);
  nand _40748_ (_02193_, _08323_, _08321_);
  nor _40749_ (_08324_, _00926_, _25051_);
  not _40750_ (_08325_, _08324_);
  nand _40751_ (_08326_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  nand _40752_ (_08327_, _08324_, _25150_);
  nand _40753_ (_02198_, _08327_, _08326_);
  nor _40754_ (_08329_, _25051_, _24059_);
  not _40755_ (_08331_, _08329_);
  nand _40756_ (_08332_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  nand _40757_ (_08333_, _08329_, _24830_);
  nand _40758_ (_02209_, _08333_, _08332_);
  nor _40759_ (_08334_, _25051_, _24999_);
  not _40760_ (_08336_, _08334_);
  nand _40761_ (_08337_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nand _40762_ (_08338_, _08334_, _25203_);
  nand _40763_ (_02223_, _08338_, _08337_);
  nor _40764_ (_08339_, _25057_, _25051_);
  not _40765_ (_08340_, _08339_);
  nand _40766_ (_08341_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  nand _40767_ (_08342_, _08339_, _25039_);
  nand _40768_ (_02227_, _08342_, _08341_);
  nor _40769_ (_08343_, _00393_, _25051_);
  not _40770_ (_08344_, _08343_);
  nand _40771_ (_08345_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  nand _40772_ (_08346_, _08343_, _24927_);
  nand _40773_ (_02237_, _08346_, _08345_);
  nand _40774_ (_08347_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  nand _40775_ (_08348_, _04021_, _24789_);
  nand _40776_ (_02247_, _08348_, _08347_);
  nand _40777_ (_08349_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  nand _40778_ (_08351_, _04021_, _25099_);
  nand _40779_ (_02250_, _08351_, _08349_);
  nand _40780_ (_08352_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  nand _40781_ (_08353_, _03867_, _25203_);
  nand _40782_ (_02253_, _08353_, _08352_);
  nor _40783_ (_08354_, _00122_, _28057_);
  nand _40784_ (_08355_, _08354_, _24789_);
  not _40785_ (_08356_, _08354_);
  nand _40786_ (_08357_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  nand _40787_ (_02256_, _08357_, _08355_);
  nand _40788_ (_08358_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nand _40789_ (_08359_, _04601_, _24830_);
  nand _40790_ (_02260_, _08359_, _08358_);
  nor _40791_ (_08360_, _07393_, _07011_);
  nand _40792_ (_08361_, _08360_, _08012_);
  nor _40793_ (_08362_, _07361_, _06907_);
  not _40794_ (_08363_, _08362_);
  nor _40795_ (_08365_, _08363_, _07181_);
  not _40796_ (_08366_, _08365_);
  nor _40797_ (_08367_, _07367_, _06886_);
  not _40798_ (_08368_, _08367_);
  nor _40799_ (_08369_, _08368_, _07025_);
  not _40800_ (_08370_, _08369_);
  nand _40801_ (_08371_, _08183_, _07434_);
  nor _40802_ (_08373_, _07376_, _07435_);
  not _40803_ (_08374_, _08373_);
  nand _40804_ (_08375_, _08374_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand _40805_ (_08376_, _08375_, _08371_);
  nand _40806_ (_08378_, _08376_, _08370_);
  nand _40807_ (_08379_, _08369_, word_in[8]);
  nand _40808_ (_08380_, _08379_, _08378_);
  nand _40809_ (_08381_, _08380_, _08366_);
  nand _40810_ (_08382_, _08365_, word_in[16]);
  nand _40811_ (_08383_, _08382_, _08381_);
  nand _40812_ (_08384_, _08383_, _08361_);
  not _40813_ (_08385_, _08361_);
  nand _40814_ (_08386_, _08385_, word_in[24]);
  nand _40815_ (_28152_, _08386_, _08384_);
  nor _40816_ (_08387_, _25165_, _25057_);
  nand _40817_ (_08389_, _08387_, _24927_);
  not _40818_ (_08390_, _08387_);
  nand _40819_ (_08391_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  nand _40820_ (_02275_, _08391_, _08389_);
  not _40821_ (_08393_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _40822_ (_08394_, _08373_, _08393_);
  nor _40823_ (_08395_, _08201_, _07435_);
  nor _40824_ (_08396_, _08395_, _08394_);
  nor _40825_ (_08397_, _08396_, _08369_);
  nor _40826_ (_08398_, _08370_, _08046_);
  nor _40827_ (_08399_, _08398_, _08397_);
  nand _40828_ (_08400_, _08399_, _08366_);
  nand _40829_ (_08401_, _07227_, word_in[17]);
  nor _40830_ (_08402_, _08401_, rst);
  nor _40831_ (_08403_, _08366_, _08402_);
  nor _40832_ (_08404_, _08403_, _08385_);
  nand _40833_ (_08405_, _08404_, _08400_);
  nand _40834_ (_08406_, _08385_, _08038_);
  nand _40835_ (_28153_, _08406_, _08405_);
  not _40836_ (_08407_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _40837_ (_08408_, _08373_, _08407_);
  nor _40838_ (_08409_, _08219_, _07435_);
  nor _40839_ (_08410_, _08409_, _08408_);
  nor _40840_ (_08411_, _08410_, _08369_);
  nor _40841_ (_08412_, _08370_, _08064_);
  nor _40842_ (_08413_, _08412_, _08411_);
  nor _40843_ (_08414_, _08413_, _08365_);
  nand _40844_ (_08415_, _08365_, word_in[18]);
  nand _40845_ (_08416_, _08415_, _08361_);
  nor _40846_ (_08417_, _08416_, _08414_);
  nor _40847_ (_08418_, _08361_, _08054_);
  nor _40848_ (_28154_, _08418_, _08417_);
  not _40849_ (_08419_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _40850_ (_08420_, _08373_, _08419_);
  nor _40851_ (_08421_, _08239_, _07435_);
  nor _40852_ (_08422_, _08421_, _08420_);
  nor _40853_ (_08423_, _08422_, _08369_);
  nor _40854_ (_08424_, _08370_, _08243_);
  nor _40855_ (_08425_, _08424_, _08423_);
  nor _40856_ (_08426_, _08425_, _08365_);
  nand _40857_ (_08427_, _08365_, word_in[19]);
  nand _40858_ (_08428_, _08427_, _08361_);
  nor _40859_ (_08429_, _08428_, _08426_);
  nor _40860_ (_08431_, _08361_, _08235_);
  nor _40861_ (_28155_, _08431_, _08429_);
  nand _40862_ (_08433_, _08354_, _25150_);
  nand _40863_ (_08434_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  nand _40864_ (_02284_, _08434_, _08433_);
  nand _40865_ (_08435_, _08374_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nand _40866_ (_08436_, _08254_, _07434_);
  nand _40867_ (_08437_, _08436_, _08435_);
  nand _40868_ (_08438_, _08437_, _08370_);
  nand _40869_ (_08439_, _08369_, word_in[12]);
  nand _40870_ (_08440_, _08439_, _08438_);
  nand _40871_ (_08441_, _08440_, _08366_);
  nand _40872_ (_08442_, _08365_, word_in[20]);
  nand _40873_ (_08443_, _08442_, _08441_);
  nand _40874_ (_08444_, _08443_, _08361_);
  nand _40875_ (_08445_, _08385_, word_in[28]);
  nand _40876_ (_28156_, _08445_, _08444_);
  not _40877_ (_08447_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _40878_ (_08448_, _08373_, _08447_);
  nor _40879_ (_08449_, _08271_, _07435_);
  nor _40880_ (_08450_, _08449_, _08448_);
  nor _40881_ (_08451_, _08450_, _08369_);
  nor _40882_ (_08452_, _08370_, _08110_);
  nor _40883_ (_08453_, _08452_, _08451_);
  nor _40884_ (_08454_, _08453_, _08365_);
  nand _40885_ (_08455_, _08365_, word_in[21]);
  nand _40886_ (_08456_, _08455_, _08361_);
  nor _40887_ (_08457_, _08456_, _08454_);
  nor _40888_ (_08458_, _08361_, _08102_);
  nor _40889_ (_28157_, _08458_, _08457_);
  not _40890_ (_08459_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _40891_ (_08460_, _08373_, _08459_);
  nor _40892_ (_08461_, _08287_, _07435_);
  nor _40893_ (_08462_, _08461_, _08460_);
  nor _40894_ (_08463_, _08462_, _08369_);
  nor _40895_ (_08464_, _08370_, _08293_);
  nor _40896_ (_08465_, _08464_, _08463_);
  nand _40897_ (_08466_, _08465_, _08366_);
  nor _40898_ (_08467_, _08366_, _08298_);
  nor _40899_ (_08468_, _08467_, _08385_);
  nand _40900_ (_08469_, _08468_, _08466_);
  nand _40901_ (_08470_, _08385_, _08283_);
  nand _40902_ (_28158_, _08470_, _08469_);
  nand _40903_ (_08471_, _08374_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _40904_ (_08472_, _08306_, _07434_);
  nand _40905_ (_08473_, _08472_, _08471_);
  nor _40906_ (_08474_, _08473_, _08369_);
  nand _40907_ (_08475_, _08369_, _07387_);
  nand _40908_ (_08476_, _08475_, _08366_);
  nor _40909_ (_08477_, _08476_, _08474_);
  nand _40910_ (_08478_, _08365_, _07400_);
  nand _40911_ (_08479_, _08478_, _08361_);
  nor _40912_ (_08480_, _08479_, _08477_);
  nor _40913_ (_08481_, _08361_, _07408_);
  nor _40914_ (_28159_, _08481_, _08480_);
  nand _40915_ (_08482_, _07810_, _28096_);
  nand _40916_ (_08483_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  nand _40917_ (_02298_, _08483_, _08482_);
  nand _40918_ (_08485_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  nand _40919_ (_08486_, _04264_, _25203_);
  nand _40920_ (_02306_, _08486_, _08485_);
  nand _40921_ (_08487_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  nand _40922_ (_08489_, _04264_, _24830_);
  nand _40923_ (_02310_, _08489_, _08487_);
  nand _40924_ (_08490_, _03850_, _25150_);
  nand _40925_ (_08491_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  nand _40926_ (_02315_, _08491_, _08490_);
  nor _40927_ (_08492_, _08142_, _00122_);
  not _40928_ (_08494_, _08492_);
  nand _40929_ (_08496_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  nand _40930_ (_08498_, _08492_, _25150_);
  nand _40931_ (_02340_, _08498_, _08496_);
  nand _40932_ (_08499_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  nand _40933_ (_08500_, _08230_, _25099_);
  nand _40934_ (_02345_, _08500_, _08499_);
  nor _40935_ (_08501_, _08142_, _00629_);
  not _40936_ (_08502_, _08501_);
  nand _40937_ (_08503_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nand _40938_ (_08504_, _08501_, _25039_);
  nand _40939_ (_02349_, _08504_, _08503_);
  nor _40940_ (_08505_, _07367_, _06925_);
  not _40941_ (_08506_, _08505_);
  nor _40942_ (_08508_, _08506_, _07025_);
  nand _40943_ (_08509_, _08183_, _07448_);
  nor _40944_ (_08510_, _07376_, _07480_);
  not _40945_ (_08511_, _08510_);
  nand _40946_ (_08512_, _08511_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _40947_ (_08513_, _08512_, _08509_);
  nor _40948_ (_08515_, _08513_, _08508_);
  nor _40949_ (_08516_, _07361_, _06886_);
  not _40950_ (_08517_, _08516_);
  nor _40951_ (_08518_, _08517_, _07181_);
  not _40952_ (_08519_, _08518_);
  nand _40953_ (_08520_, _08508_, _08027_);
  nand _40954_ (_08521_, _08520_, _08519_);
  nor _40955_ (_08522_, _08521_, _08515_);
  nor _40956_ (_08524_, _08013_, _06907_);
  nand _40957_ (_08525_, _08524_, _07392_);
  nand _40958_ (_08526_, _08518_, word_in[16]);
  nand _40959_ (_08527_, _08526_, _08525_);
  nor _40960_ (_08528_, _08527_, _08522_);
  nor _40961_ (_08529_, _08525_, word_in[24]);
  nor _40962_ (_28175_[0], _08529_, _08528_);
  nand _40963_ (_08531_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  nand _40964_ (_08532_, _08329_, _24789_);
  nand _40965_ (_02359_, _08532_, _08531_);
  not _40966_ (_08533_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _40967_ (_08534_, _08510_, _08533_);
  nor _40968_ (_08536_, _08201_, _07480_);
  nor _40969_ (_08537_, _08536_, _08534_);
  nor _40970_ (_08538_, _08537_, _08508_);
  not _40971_ (_08540_, _08508_);
  nor _40972_ (_08541_, _08540_, _08046_);
  nor _40973_ (_08543_, _08541_, _08538_);
  nor _40974_ (_08544_, _08543_, _08518_);
  nand _40975_ (_08545_, _08518_, word_in[17]);
  nand _40976_ (_08546_, _08545_, _08525_);
  nor _40977_ (_08547_, _08546_, _08544_);
  nor _40978_ (_08548_, _08525_, word_in[25]);
  nor _40979_ (_28175_[1], _08548_, _08547_);
  nor _40980_ (_08549_, _25051_, _24978_);
  not _40981_ (_08551_, _08549_);
  nand _40982_ (_08552_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  nand _40983_ (_08554_, _08549_, _28096_);
  nand _40984_ (_02363_, _08554_, _08552_);
  nand _40985_ (_08556_, _08524_, _08054_);
  nand _40986_ (_08557_, _08510_, word_in[2]);
  nand _40987_ (_08558_, _08511_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _40988_ (_08560_, _08558_, _08557_);
  nand _40989_ (_08561_, _08560_, _08540_);
  nand _40990_ (_08562_, _08508_, word_in[10]);
  nand _40991_ (_08563_, _08562_, _08561_);
  nand _40992_ (_08564_, _08563_, _08519_);
  nand _40993_ (_08565_, _08518_, word_in[18]);
  nand _40994_ (_08566_, _08565_, _08564_);
  nand _40995_ (_08567_, _08566_, _08525_);
  nand _40996_ (_28175_[2], _08567_, _08556_);
  nand _40997_ (_08568_, _08524_, _08235_);
  nand _40998_ (_08569_, _08510_, word_in[3]);
  nand _40999_ (_08570_, _08511_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nand _41000_ (_08571_, _08570_, _08569_);
  nand _41001_ (_08572_, _08571_, _08540_);
  nand _41002_ (_08573_, _08508_, word_in[11]);
  nand _41003_ (_08574_, _08573_, _08572_);
  nand _41004_ (_08575_, _08574_, _08519_);
  nand _41005_ (_08576_, _08518_, word_in[19]);
  nand _41006_ (_08577_, _08576_, _08575_);
  nand _41007_ (_08579_, _08577_, _08525_);
  nand _41008_ (_28175_[3], _08579_, _08568_);
  nand _41009_ (_08580_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nand _41010_ (_08581_, _04015_, _28096_);
  nand _41011_ (_02368_, _08581_, _08580_);
  nand _41012_ (_08583_, _08524_, _08084_);
  nand _41013_ (_08584_, _08511_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand _41014_ (_08585_, _08254_, _07448_);
  nand _41015_ (_08587_, _08585_, _08584_);
  nand _41016_ (_08588_, _08587_, _08540_);
  nand _41017_ (_08590_, _08508_, word_in[12]);
  nand _41018_ (_08592_, _08590_, _08588_);
  nand _41019_ (_08593_, _08592_, _08519_);
  nand _41020_ (_08594_, _08518_, word_in[20]);
  nand _41021_ (_08595_, _08594_, _08593_);
  nand _41022_ (_08596_, _08595_, _08525_);
  nand _41023_ (_28175_[4], _08596_, _08583_);
  nand _41024_ (_08597_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nand _41025_ (_08599_, _04610_, _25039_);
  nand _41026_ (_02371_, _08599_, _08597_);
  nand _41027_ (_08602_, _08524_, _08102_);
  nor _41028_ (_08603_, _08511_, _08106_);
  not _41029_ (_08604_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _41030_ (_08605_, _08510_, _08604_);
  nor _41031_ (_08606_, _08605_, _08603_);
  nor _41032_ (_08607_, _08606_, _08508_);
  nor _41033_ (_08608_, _08540_, _08110_);
  nor _41034_ (_08609_, _08608_, _08607_);
  nand _41035_ (_08610_, _08609_, _08519_);
  not _41036_ (_08611_, _08525_);
  nand _41037_ (_08612_, _07227_, word_in[21]);
  nor _41038_ (_08613_, _08612_, rst);
  nor _41039_ (_08614_, _08519_, _08613_);
  nor _41040_ (_08615_, _08614_, _08611_);
  nand _41041_ (_08616_, _08615_, _08610_);
  nand _41042_ (_28160_, _08616_, _08602_);
  nand _41043_ (_08617_, _08524_, _08283_);
  not _41044_ (_08618_, word_in[6]);
  nor _41045_ (_08619_, _08511_, _08618_);
  not _41046_ (_08620_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _41047_ (_08622_, _08510_, _08620_);
  nor _41048_ (_08623_, _08622_, _08619_);
  nor _41049_ (_08624_, _08623_, _08508_);
  nor _41050_ (_08625_, _08540_, _08293_);
  nor _41051_ (_08627_, _08625_, _08624_);
  nand _41052_ (_08629_, _08627_, _08519_);
  nor _41053_ (_08630_, _08519_, _08298_);
  nor _41054_ (_08631_, _08630_, _08611_);
  nand _41055_ (_08633_, _08631_, _08629_);
  nand _41056_ (_28175_[6], _08633_, _08617_);
  not _41057_ (_08635_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor _41058_ (_08636_, _08510_, _08635_);
  nor _41059_ (_08637_, _08307_, _07480_);
  nor _41060_ (_08638_, _08637_, _08636_);
  nor _41061_ (_08639_, _08638_, _08508_);
  nor _41062_ (_08640_, _08540_, _07387_);
  nor _41063_ (_08641_, _08640_, _08639_);
  nor _41064_ (_08642_, _08641_, _08518_);
  nand _41065_ (_08643_, _08518_, _07400_);
  nand _41066_ (_08644_, _08643_, _08525_);
  nor _41067_ (_08645_, _08644_, _08642_);
  nor _41068_ (_08647_, _08525_, word_in[31]);
  nor _41069_ (_28175_[7], _08647_, _08645_);
  nand _41070_ (_08649_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nand _41071_ (_08650_, _04021_, _25150_);
  nand _41072_ (_02391_, _08650_, _08649_);
  nand _41073_ (_08651_, _28105_, _25099_);
  nand _41074_ (_08652_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  nand _41075_ (_02395_, _08652_, _08651_);
  nor _41076_ (_08653_, _28104_, _24978_);
  nand _41077_ (_08654_, _08653_, _24789_);
  not _41078_ (_08655_, _08653_);
  nand _41079_ (_08656_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  nand _41080_ (_02400_, _08656_, _08654_);
  nand _41081_ (_08658_, _07810_, _25150_);
  nand _41082_ (_08659_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  nand _41083_ (_02405_, _08659_, _08658_);
  nand _41084_ (_08660_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  nand _41085_ (_08661_, _04264_, _24789_);
  nand _41086_ (_02418_, _08661_, _08660_);
  nand _41087_ (_08663_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  nand _41088_ (_08665_, _01216_, _25039_);
  nand _41089_ (_02423_, _08665_, _08663_);
  nand _41090_ (_08666_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  nand _41091_ (_08667_, _08144_, _25039_);
  nand _41092_ (_02427_, _08667_, _08666_);
  nand _41093_ (_08668_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  nand _41094_ (_08669_, _08153_, _28096_);
  nand _41095_ (_02430_, _08669_, _08668_);
  nand _41096_ (_08670_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  nand _41097_ (_08671_, _08212_, _25039_);
  nand _41098_ (_02440_, _08671_, _08670_);
  nand _41099_ (_08672_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  nand _41100_ (_08673_, _08339_, _24927_);
  nand _41101_ (_02449_, _08673_, _08672_);
  nand _41102_ (_08674_, _08011_, _07271_);
  nor _41103_ (_08676_, _08674_, _06886_);
  nor _41104_ (_08677_, _07767_, _07361_);
  not _41105_ (_08678_, _08677_);
  nor _41106_ (_08679_, _08678_, _06925_);
  not _41107_ (_08680_, _08679_);
  nor _41108_ (_08681_, _07367_, _07480_);
  nor _41109_ (_08682_, _07376_, _07473_);
  not _41110_ (_08683_, _08682_);
  nand _41111_ (_08684_, _08683_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand _41112_ (_08685_, _08183_, _07472_);
  nand _41113_ (_08686_, _08685_, _08684_);
  nor _41114_ (_08687_, _08686_, _08681_);
  not _41115_ (_08688_, _08681_);
  nor _41116_ (_08690_, _08688_, word_in[8]);
  nor _41117_ (_08691_, _08690_, _08687_);
  nand _41118_ (_08692_, _08691_, _08680_);
  nand _41119_ (_08693_, _07227_, word_in[16]);
  nor _41120_ (_08694_, _08693_, rst);
  nand _41121_ (_08695_, _08679_, _08694_);
  nand _41122_ (_08696_, _08695_, _08692_);
  nor _41123_ (_08697_, _08696_, _08676_);
  nand _41124_ (_08698_, _07354_, word_in[24]);
  nor _41125_ (_08699_, _08698_, rst);
  not _41126_ (_08700_, _08676_);
  nor _41127_ (_08702_, _08700_, _08699_);
  nor _41128_ (_28176_[0], _08702_, _08697_);
  nand _41129_ (_08705_, _08683_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nand _41130_ (_08707_, _08200_, _07472_);
  nand _41131_ (_08708_, _08707_, _08705_);
  nand _41132_ (_08709_, _08708_, _08688_);
  nand _41133_ (_08710_, _08681_, word_in[9]);
  nand _41134_ (_08711_, _08710_, _08709_);
  nand _41135_ (_08712_, _08711_, _08680_);
  nand _41136_ (_08713_, _08679_, _08402_);
  nand _41137_ (_08714_, _08713_, _08712_);
  nand _41138_ (_08715_, _08714_, _08700_);
  nand _41139_ (_08716_, _08676_, _08038_);
  nand _41140_ (_28176_[1], _08716_, _08715_);
  nand _41141_ (_08717_, _07227_, word_in[18]);
  nor _41142_ (_08719_, _08717_, rst);
  nand _41143_ (_08720_, _08679_, _08719_);
  nand _41144_ (_08721_, _08682_, word_in[2]);
  nand _41145_ (_08723_, _08683_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand _41146_ (_08725_, _08723_, _08721_);
  nand _41147_ (_08727_, _08725_, _08688_);
  nand _41148_ (_08728_, _08681_, word_in[10]);
  nand _41149_ (_08729_, _08728_, _08727_);
  nand _41150_ (_08730_, _08729_, _08680_);
  nand _41151_ (_08731_, _08730_, _08720_);
  nand _41152_ (_08732_, _08731_, _08700_);
  nand _41153_ (_08733_, _08676_, _08054_);
  nand _41154_ (_28176_[2], _08733_, _08732_);
  nand _41155_ (_08735_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  nand _41156_ (_08736_, _25099_, _25052_);
  nand _41157_ (_02466_, _08736_, _08735_);
  not _41158_ (_08737_, word_in[3]);
  nor _41159_ (_08738_, _08683_, _08737_);
  not _41160_ (_08739_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _41161_ (_08740_, _08682_, _08739_);
  nor _41162_ (_08741_, _08740_, _08738_);
  nor _41163_ (_08742_, _08741_, _08681_);
  nor _41164_ (_08744_, _08688_, _08243_);
  nor _41165_ (_08745_, _08744_, _08742_);
  nor _41166_ (_08746_, _08745_, _08679_);
  nand _41167_ (_08747_, _08679_, _08248_);
  nand _41168_ (_08749_, _08747_, _08700_);
  nor _41169_ (_08750_, _08749_, _08746_);
  nor _41170_ (_08751_, _08700_, _08235_);
  nor _41171_ (_28176_[3], _08751_, _08750_);
  nand _41172_ (_08753_, _08683_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nand _41173_ (_08754_, _08254_, _07472_);
  nand _41174_ (_08756_, _08754_, _08753_);
  nor _41175_ (_08757_, _08756_, _08681_);
  nor _41176_ (_08758_, _08688_, word_in[12]);
  nor _41177_ (_08759_, _08758_, _08757_);
  nor _41178_ (_08760_, _08759_, _08679_);
  nand _41179_ (_08761_, _07227_, word_in[20]);
  nor _41180_ (_08763_, _08761_, rst);
  nor _41181_ (_08764_, _08680_, _08763_);
  nor _41182_ (_08765_, _08764_, _08760_);
  nor _41183_ (_08766_, _08765_, _08676_);
  nor _41184_ (_08767_, _08700_, _08084_);
  nor _41185_ (_28176_[4], _08767_, _08766_);
  nor _41186_ (_08768_, _08683_, _08106_);
  not _41187_ (_08769_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _41188_ (_08770_, _08682_, _08769_);
  nor _41189_ (_08771_, _08770_, _08768_);
  nor _41190_ (_08772_, _08771_, _08681_);
  nor _41191_ (_08773_, _08688_, _08110_);
  nor _41192_ (_08774_, _08773_, _08772_);
  nor _41193_ (_08775_, _08774_, _08679_);
  nand _41194_ (_08776_, _08679_, _08613_);
  nand _41195_ (_08777_, _08776_, _08700_);
  nor _41196_ (_08778_, _08777_, _08775_);
  nor _41197_ (_08779_, _08700_, _08102_);
  nor _41198_ (_28176_[5], _08779_, _08778_);
  nor _41199_ (_08780_, _08683_, _08618_);
  not _41200_ (_08781_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _41201_ (_08782_, _08682_, _08781_);
  nor _41202_ (_08783_, _08782_, _08780_);
  nor _41203_ (_08784_, _08783_, _08681_);
  nor _41204_ (_08785_, _08688_, _08293_);
  nor _41205_ (_08786_, _08785_, _08784_);
  nor _41206_ (_08787_, _08786_, _08679_);
  nand _41207_ (_08788_, _08679_, _08298_);
  nand _41208_ (_08789_, _08788_, _08700_);
  nor _41209_ (_08790_, _08789_, _08787_);
  nor _41210_ (_08791_, _08700_, _08283_);
  nor _41211_ (_28176_[6], _08791_, _08790_);
  nand _41212_ (_08792_, _08679_, _07400_);
  nand _41213_ (_08793_, _08683_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _41214_ (_08794_, _08306_, _07472_);
  nand _41215_ (_08795_, _08794_, _08793_);
  nand _41216_ (_08796_, _08795_, _08688_);
  nand _41217_ (_08797_, _08681_, word_in[15]);
  nand _41218_ (_08799_, _08797_, _08796_);
  nand _41219_ (_08800_, _08799_, _08680_);
  nand _41220_ (_08801_, _08800_, _08792_);
  nand _41221_ (_08802_, _08801_, _08700_);
  nand _41222_ (_08803_, _08676_, _07408_);
  nand _41223_ (_28176_[7], _08803_, _08802_);
  nand _41224_ (_08804_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  nand _41225_ (_08805_, _04610_, _24927_);
  nand _41226_ (_02483_, _08805_, _08804_);
  nor _41227_ (_08806_, _00926_, _28104_);
  nand _41228_ (_08807_, _08806_, _24830_);
  not _41229_ (_08808_, _08806_);
  nand _41230_ (_08809_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  nand _41231_ (_02489_, _08809_, _08807_);
  nand _41232_ (_08811_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  nand _41233_ (_08812_, _08212_, _24927_);
  nand _41234_ (_02496_, _08812_, _08811_);
  nor _41235_ (_08813_, _08678_, _07011_);
  nor _41236_ (_08814_, _08179_, _07578_);
  not _41237_ (_08815_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _41238_ (_08816_, _07376_, _07504_);
  nor _41239_ (_08817_, _08816_, _08815_);
  not _41240_ (_08818_, _08816_);
  nor _41241_ (_08819_, _08818_, _08182_);
  nor _41242_ (_08820_, _08819_, _08817_);
  nor _41243_ (_08821_, _08820_, _08814_);
  not _41244_ (_08822_, _08814_);
  nor _41245_ (_08824_, _08822_, _08027_);
  nor _41246_ (_08825_, _08824_, _08821_);
  nor _41247_ (_08827_, _08825_, _08813_);
  nor _41248_ (_08828_, _08674_, _06925_);
  not _41249_ (_08829_, _08828_);
  nand _41250_ (_08831_, _08813_, _08694_);
  nand _41251_ (_08833_, _08831_, _08829_);
  nor _41252_ (_08834_, _08833_, _08827_);
  nor _41253_ (_08835_, _08829_, _08699_);
  nor _41254_ (_28177_[0], _08835_, _08834_);
  nor _41255_ (_08836_, _08818_, _08042_);
  not _41256_ (_08837_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _41257_ (_08838_, _08816_, _08837_);
  nor _41258_ (_08839_, _08838_, _08836_);
  nor _41259_ (_08840_, _08839_, _08814_);
  nor _41260_ (_08841_, _08822_, _08046_);
  nor _41261_ (_08842_, _08841_, _08840_);
  nor _41262_ (_08843_, _08842_, _08813_);
  nand _41263_ (_08844_, _08813_, _08402_);
  nand _41264_ (_08845_, _08844_, _08829_);
  nor _41265_ (_08847_, _08845_, _08843_);
  nor _41266_ (_08848_, _08829_, _08038_);
  nor _41267_ (_28177_[1], _08848_, _08847_);
  nor _41268_ (_08849_, _08816_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _41269_ (_08851_, _08818_, word_in[2]);
  nor _41270_ (_08852_, _08851_, _08849_);
  nor _41271_ (_08853_, _08852_, _08814_);
  nor _41272_ (_08854_, _08822_, word_in[10]);
  nor _41273_ (_08856_, _08854_, _08853_);
  nor _41274_ (_08857_, _08856_, _08813_);
  not _41275_ (_08858_, _08813_);
  nor _41276_ (_08859_, _08858_, _08719_);
  nor _41277_ (_08860_, _08859_, _08857_);
  nor _41278_ (_08861_, _08860_, _08828_);
  nor _41279_ (_08862_, _08829_, _08054_);
  nor _41280_ (_28177_[2], _08862_, _08861_);
  nor _41281_ (_08863_, _08818_, _08737_);
  not _41282_ (_08864_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _41283_ (_08865_, _08816_, _08864_);
  nor _41284_ (_08866_, _08865_, _08863_);
  nor _41285_ (_08868_, _08866_, _08814_);
  nor _41286_ (_08870_, _08822_, _08243_);
  nor _41287_ (_08872_, _08870_, _08868_);
  nor _41288_ (_08873_, _08872_, _08813_);
  nand _41289_ (_08874_, _08813_, _08248_);
  nand _41290_ (_08875_, _08874_, _08829_);
  nor _41291_ (_08876_, _08875_, _08873_);
  nor _41292_ (_08877_, _08829_, _08235_);
  nor _41293_ (_28177_[3], _08877_, _08876_);
  not _41294_ (_08878_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _41295_ (_08879_, _08816_, _08878_);
  nor _41296_ (_08880_, _08818_, _08088_);
  nor _41297_ (_08881_, _08880_, _08879_);
  nor _41298_ (_08882_, _08881_, _08814_);
  nor _41299_ (_08883_, _08822_, _08092_);
  nor _41300_ (_08884_, _08883_, _08882_);
  nor _41301_ (_08885_, _08884_, _08813_);
  nand _41302_ (_08887_, _08813_, _08763_);
  nand _41303_ (_08889_, _08887_, _08829_);
  nor _41304_ (_08891_, _08889_, _08885_);
  nor _41305_ (_08892_, _08829_, _08084_);
  nor _41306_ (_28177_[4], _08892_, _08891_);
  nand _41307_ (_08894_, _08814_, _08110_);
  nor _41308_ (_08896_, _08816_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _41309_ (_08898_, _08818_, word_in[5]);
  nor _41310_ (_08900_, _08898_, _08896_);
  nor _41311_ (_08901_, _08900_, _08814_);
  nor _41312_ (_08902_, _08901_, _08813_);
  nand _41313_ (_08903_, _08902_, _08894_);
  nand _41314_ (_08905_, _08813_, _08613_);
  nand _41315_ (_08906_, _08905_, _08903_);
  nor _41316_ (_08907_, _08906_, _08828_);
  nor _41317_ (_08908_, _08829_, _08102_);
  nor _41318_ (_28177_[5], _08908_, _08907_);
  nand _41319_ (_08909_, _08814_, _08293_);
  nand _41320_ (_08910_, _08818_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nand _41321_ (_08911_, _08816_, word_in[6]);
  nand _41322_ (_08912_, _08911_, _08910_);
  nor _41323_ (_08913_, _08912_, _08814_);
  nor _41324_ (_08914_, _08913_, _08813_);
  nand _41325_ (_08915_, _08914_, _08909_);
  nand _41326_ (_08916_, _08813_, _08298_);
  nand _41327_ (_08917_, _08916_, _08915_);
  nand _41328_ (_08918_, _08917_, _08829_);
  nand _41329_ (_08919_, _08828_, _08283_);
  nand _41330_ (_28177_[6], _08919_, _08918_);
  nand _41331_ (_08920_, _08813_, _07400_);
  nand _41332_ (_08921_, _08814_, _07387_);
  nand _41333_ (_08922_, _08816_, word_in[7]);
  nand _41334_ (_08924_, _08818_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _41335_ (_08925_, _08924_, _08922_);
  nor _41336_ (_08927_, _08925_, _08814_);
  nor _41337_ (_08929_, _08927_, _08813_);
  nand _41338_ (_08931_, _08929_, _08921_);
  nand _41339_ (_08933_, _08931_, _08920_);
  nand _41340_ (_08934_, _08933_, _08829_);
  nand _41341_ (_08935_, _08828_, _07408_);
  nand _41342_ (_28177_[7], _08935_, _08934_);
  nor _41343_ (_08936_, _08678_, _06907_);
  nor _41344_ (_08937_, _08368_, _07578_);
  not _41345_ (_08938_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _41346_ (_08940_, _07376_, _07589_);
  nor _41347_ (_08942_, _08940_, _08938_);
  not _41348_ (_08943_, _08940_);
  nor _41349_ (_08945_, _08943_, _08182_);
  nor _41350_ (_08946_, _08945_, _08942_);
  nor _41351_ (_08947_, _08946_, _08937_);
  not _41352_ (_08949_, _08937_);
  nor _41353_ (_08951_, _08949_, _08027_);
  nor _41354_ (_08953_, _08951_, _08947_);
  nor _41355_ (_08954_, _08953_, _08936_);
  nor _41356_ (_08955_, _08674_, _07011_);
  not _41357_ (_08956_, _08955_);
  nand _41358_ (_08958_, _08936_, _08694_);
  nand _41359_ (_08959_, _08958_, _08956_);
  nor _41360_ (_08960_, _08959_, _08954_);
  nor _41361_ (_08961_, _08956_, _08699_);
  nor _41362_ (_28178_[0], _08961_, _08960_);
  not _41363_ (_08964_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _41364_ (_08966_, _08940_, _08964_);
  nor _41365_ (_08967_, _08943_, _08042_);
  nor _41366_ (_08968_, _08967_, _08966_);
  nor _41367_ (_08970_, _08968_, _08937_);
  nor _41368_ (_08972_, _08949_, _08046_);
  nor _41369_ (_08973_, _08972_, _08970_);
  nor _41370_ (_08974_, _08973_, _08936_);
  nand _41371_ (_08975_, _08936_, _08402_);
  nand _41372_ (_08977_, _08975_, _08956_);
  nor _41373_ (_08979_, _08977_, _08974_);
  nor _41374_ (_08981_, _08956_, _08038_);
  nor _41375_ (_28178_[1], _08981_, _08979_);
  not _41376_ (_08982_, _08936_);
  not _41377_ (_08983_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand _41378_ (_08984_, _08943_, _08983_);
  nand _41379_ (_08985_, _08940_, _08059_);
  nand _41380_ (_08987_, _08985_, _08984_);
  nand _41381_ (_08988_, _08987_, _08949_);
  nand _41382_ (_08989_, _08937_, _08064_);
  nand _41383_ (_08990_, _08989_, _08988_);
  nand _41384_ (_08991_, _08990_, _08982_);
  nor _41385_ (_08992_, _08982_, _08719_);
  nor _41386_ (_08993_, _08992_, _08955_);
  nand _41387_ (_08994_, _08993_, _08991_);
  nand _41388_ (_08995_, _08955_, _08054_);
  nand _41389_ (_28178_[2], _08995_, _08994_);
  not _41390_ (_08996_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _41391_ (_08997_, _08940_, _08996_);
  nor _41392_ (_08998_, _08943_, _08737_);
  nor _41393_ (_08999_, _08998_, _08997_);
  nor _41394_ (_09000_, _08999_, _08937_);
  nor _41395_ (_09001_, _08949_, _08243_);
  nor _41396_ (_09002_, _09001_, _09000_);
  nor _41397_ (_09003_, _09002_, _08936_);
  nand _41398_ (_09004_, _08936_, _08248_);
  nand _41399_ (_09005_, _09004_, _08956_);
  nor _41400_ (_09006_, _09005_, _09003_);
  nor _41401_ (_09007_, _08956_, _08235_);
  nor _41402_ (_28178_[3], _09007_, _09006_);
  not _41403_ (_09008_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _41404_ (_09010_, _08940_, _09008_);
  nor _41405_ (_09012_, _08943_, _08088_);
  nor _41406_ (_09013_, _09012_, _09010_);
  nor _41407_ (_09015_, _09013_, _08937_);
  nor _41408_ (_09017_, _08949_, _08092_);
  nor _41409_ (_09018_, _09017_, _09015_);
  nor _41410_ (_09019_, _09018_, _08936_);
  nand _41411_ (_09021_, _08936_, _08763_);
  nand _41412_ (_09022_, _09021_, _08956_);
  nor _41413_ (_09023_, _09022_, _09019_);
  nor _41414_ (_09025_, _08956_, _08084_);
  nor _41415_ (_28178_[4], _09025_, _09023_);
  not _41416_ (_09027_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nand _41417_ (_09028_, _08943_, _09027_);
  nand _41418_ (_09029_, _08940_, _08106_);
  nand _41419_ (_09030_, _09029_, _09028_);
  nand _41420_ (_09031_, _09030_, _08949_);
  nand _41421_ (_09032_, _08937_, _08110_);
  nand _41422_ (_09033_, _09032_, _09031_);
  nand _41423_ (_09034_, _09033_, _08982_);
  nor _41424_ (_09035_, _08982_, _08613_);
  nor _41425_ (_09036_, _09035_, _08955_);
  nand _41426_ (_09037_, _09036_, _09034_);
  nand _41427_ (_09038_, _08955_, _08102_);
  nand _41428_ (_28178_[5], _09038_, _09037_);
  nand _41429_ (_09040_, _08936_, _08298_);
  nand _41430_ (_09041_, _08937_, _08293_);
  nand _41431_ (_09042_, _08943_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nand _41432_ (_09043_, _08940_, word_in[6]);
  nand _41433_ (_09044_, _09043_, _09042_);
  nor _41434_ (_09045_, _09044_, _08937_);
  nor _41435_ (_09046_, _09045_, _08936_);
  nand _41436_ (_09047_, _09046_, _09041_);
  nand _41437_ (_09048_, _09047_, _09040_);
  nand _41438_ (_09049_, _09048_, _08956_);
  nand _41439_ (_09051_, _08955_, _08283_);
  nand _41440_ (_28178_[6], _09051_, _09049_);
  not _41441_ (_09052_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nor _41442_ (_09053_, _08940_, _09052_);
  nor _41443_ (_09054_, _08943_, _07381_);
  nor _41444_ (_09055_, _09054_, _09053_);
  nor _41445_ (_09056_, _09055_, _08937_);
  nor _41446_ (_09057_, _08949_, _07387_);
  nor _41447_ (_09058_, _09057_, _09056_);
  nor _41448_ (_09059_, _09058_, _08936_);
  nand _41449_ (_09061_, _08936_, _07400_);
  nand _41450_ (_09063_, _09061_, _08956_);
  nor _41451_ (_09064_, _09063_, _09059_);
  nor _41452_ (_09065_, _08956_, _07408_);
  nor _41453_ (_28178_[7], _09065_, _09064_);
  nor _41454_ (_09067_, _08674_, _06907_);
  not _41455_ (_09069_, _09067_);
  nor _41456_ (_09070_, _08506_, _07578_);
  nand _41457_ (_09071_, _09070_, _08027_);
  nor _41458_ (_09073_, _08678_, _06886_);
  nor _41459_ (_09074_, _07376_, _07658_);
  nand _41460_ (_09075_, _09074_, word_in[0]);
  not _41461_ (_09076_, _09074_);
  nand _41462_ (_09078_, _09076_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand _41463_ (_09079_, _09078_, _09075_);
  nor _41464_ (_09080_, _09079_, _09070_);
  nor _41465_ (_09082_, _09080_, _09073_);
  nand _41466_ (_09083_, _09082_, _09071_);
  nand _41467_ (_09084_, _09073_, _08694_);
  nand _41468_ (_09085_, _09084_, _09083_);
  nand _41469_ (_09086_, _09085_, _09069_);
  nand _41470_ (_09087_, _09067_, _08699_);
  nand _41471_ (_28179_[0], _09087_, _09086_);
  nand _41472_ (_09088_, _09070_, _08046_);
  nand _41473_ (_09090_, _09074_, word_in[1]);
  nand _41474_ (_09091_, _09076_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nand _41475_ (_09092_, _09091_, _09090_);
  nor _41476_ (_09093_, _09092_, _09070_);
  nor _41477_ (_09094_, _09093_, _09073_);
  nand _41478_ (_09096_, _09094_, _09088_);
  nand _41479_ (_09097_, _09073_, _08402_);
  nand _41480_ (_09098_, _09097_, _09096_);
  nand _41481_ (_09099_, _09098_, _09069_);
  nand _41482_ (_09100_, _09067_, _08038_);
  nand _41483_ (_28179_[1], _09100_, _09099_);
  nor _41484_ (_09101_, _09074_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _41485_ (_09102_, _09076_, word_in[2]);
  nor _41486_ (_09103_, _09102_, _09101_);
  nor _41487_ (_09104_, _09103_, _09070_);
  not _41488_ (_09105_, _09070_);
  nor _41489_ (_09107_, _09105_, word_in[10]);
  nor _41490_ (_09109_, _09107_, _09104_);
  nor _41491_ (_09111_, _09109_, _09073_);
  not _41492_ (_09113_, _09073_);
  nor _41493_ (_09115_, _09113_, _08719_);
  nor _41494_ (_09116_, _09115_, _09111_);
  nor _41495_ (_09117_, _09116_, _09067_);
  nor _41496_ (_09118_, _09069_, _08054_);
  nor _41497_ (_28179_[2], _09118_, _09117_);
  nor _41498_ (_09119_, _09074_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _41499_ (_09120_, _09076_, word_in[3]);
  nor _41500_ (_09121_, _09120_, _09119_);
  nor _41501_ (_09122_, _09121_, _09070_);
  nor _41502_ (_09123_, _09105_, word_in[11]);
  nor _41503_ (_09124_, _09123_, _09122_);
  nor _41504_ (_09125_, _09124_, _09073_);
  nor _41505_ (_09126_, _09113_, _08248_);
  nor _41506_ (_09127_, _09126_, _09125_);
  nor _41507_ (_09128_, _09127_, _09067_);
  nor _41508_ (_09129_, _09069_, _08235_);
  nor _41509_ (_28179_[3], _09129_, _09128_);
  nand _41510_ (_09130_, _09073_, _08763_);
  nand _41511_ (_09131_, _09070_, _08092_);
  nand _41512_ (_09132_, _09074_, word_in[4]);
  nand _41513_ (_09133_, _09076_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand _41514_ (_09134_, _09133_, _09132_);
  nor _41515_ (_09135_, _09134_, _09070_);
  nor _41516_ (_09136_, _09135_, _09073_);
  nand _41517_ (_09137_, _09136_, _09131_);
  nand _41518_ (_09138_, _09137_, _09130_);
  nand _41519_ (_09139_, _09138_, _09069_);
  nand _41520_ (_09140_, _09067_, _08084_);
  nand _41521_ (_28179_[4], _09140_, _09139_);
  nand _41522_ (_09142_, _08387_, _25150_);
  nand _41523_ (_09143_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nand _41524_ (_02634_, _09143_, _09142_);
  nand _41525_ (_09144_, _09070_, _08110_);
  nand _41526_ (_09145_, _09074_, word_in[5]);
  nand _41527_ (_09146_, _09076_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nand _41528_ (_09147_, _09146_, _09145_);
  nor _41529_ (_09148_, _09147_, _09070_);
  nor _41530_ (_09149_, _09148_, _09073_);
  nand _41531_ (_09150_, _09149_, _09144_);
  nand _41532_ (_09151_, _09073_, _08613_);
  nand _41533_ (_09152_, _09151_, _09150_);
  nand _41534_ (_09153_, _09152_, _09069_);
  nand _41535_ (_09154_, _09067_, _08102_);
  nand _41536_ (_28179_[5], _09154_, _09153_);
  nand _41537_ (_09156_, _09070_, _08293_);
  nand _41538_ (_09157_, _09074_, word_in[6]);
  nand _41539_ (_09158_, _09076_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nand _41540_ (_09160_, _09158_, _09157_);
  nor _41541_ (_09161_, _09160_, _09070_);
  nor _41542_ (_09162_, _09161_, _09073_);
  nand _41543_ (_09163_, _09162_, _09156_);
  nand _41544_ (_09164_, _09073_, _08298_);
  nand _41545_ (_09165_, _09164_, _09163_);
  nand _41546_ (_09166_, _09165_, _09069_);
  nand _41547_ (_09167_, _09067_, _08283_);
  nand _41548_ (_28179_[6], _09167_, _09166_);
  nand _41549_ (_09168_, _09073_, _07400_);
  nand _41550_ (_09170_, _09070_, _07387_);
  nand _41551_ (_09171_, _09074_, word_in[7]);
  nand _41552_ (_09172_, _09076_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _41553_ (_09173_, _09172_, _09171_);
  nor _41554_ (_09174_, _09173_, _09070_);
  nor _41555_ (_09175_, _09174_, _09073_);
  nand _41556_ (_09176_, _09175_, _09170_);
  nand _41557_ (_09177_, _09176_, _09168_);
  nand _41558_ (_09178_, _09177_, _09069_);
  nand _41559_ (_09179_, _09067_, _07408_);
  nand _41560_ (_28179_[7], _09179_, _09178_);
  nor _41561_ (_09180_, _07395_, _07263_);
  not _41562_ (_09181_, _09180_);
  nor _41563_ (_09182_, _09181_, _06886_);
  not _41564_ (_09184_, _09182_);
  nor _41565_ (_09185_, _07367_, _07658_);
  not _41566_ (_09186_, _09185_);
  nor _41567_ (_09187_, _07716_, _07376_);
  nand _41568_ (_09188_, _09187_, word_in[0]);
  not _41569_ (_09189_, _09187_);
  nand _41570_ (_09190_, _09189_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nand _41571_ (_09191_, _09190_, _09188_);
  nand _41572_ (_09192_, _09191_, _09186_);
  nand _41573_ (_09193_, _09185_, word_in[8]);
  nand _41574_ (_09194_, _09193_, _09192_);
  nor _41575_ (_09195_, _07361_, _07589_);
  not _41576_ (_09196_, _09195_);
  nand _41577_ (_09197_, _09196_, _09194_);
  nand _41578_ (_09198_, _09195_, word_in[16]);
  nand _41579_ (_09199_, _09198_, _09197_);
  nand _41580_ (_09200_, _09199_, _09184_);
  nand _41581_ (_09201_, _09182_, _08699_);
  nand _41582_ (_28161_, _09201_, _09200_);
  nand _41583_ (_09202_, _09187_, word_in[1]);
  nand _41584_ (_09203_, _09189_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nand _41585_ (_09204_, _09203_, _09202_);
  nand _41586_ (_09205_, _09204_, _09186_);
  nand _41587_ (_09206_, _09185_, word_in[9]);
  nand _41588_ (_09207_, _09206_, _09205_);
  nand _41589_ (_09208_, _09207_, _09196_);
  nand _41590_ (_09209_, _09195_, word_in[17]);
  nand _41591_ (_09210_, _09209_, _09208_);
  nand _41592_ (_09211_, _09210_, _09184_);
  nand _41593_ (_09212_, _09182_, _08038_);
  nand _41594_ (_28162_, _09212_, _09211_);
  nand _41595_ (_09213_, _07359_, _06925_);
  nor _41596_ (_09214_, _07361_, _07169_);
  nand _41597_ (_09215_, _09214_, _09213_);
  nor _41598_ (_09216_, _09187_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _41599_ (_09217_, _09189_, word_in[2]);
  nor _41600_ (_09218_, _09217_, _09216_);
  nor _41601_ (_09219_, _09218_, _09185_);
  nor _41602_ (_09220_, _09186_, word_in[10]);
  nor _41603_ (_09221_, _09220_, _09219_);
  nand _41604_ (_09222_, _09221_, _09215_);
  not _41605_ (_09223_, _09214_);
  nor _41606_ (_09224_, _09223_, _06925_);
  nand _41607_ (_09225_, _09224_, word_in[18]);
  nand _41608_ (_09226_, _09225_, _09222_);
  nor _41609_ (_09227_, _09226_, _09182_);
  nor _41610_ (_09228_, _09184_, _08054_);
  nor _41611_ (_28163_, _09228_, _09227_);
  nand _41612_ (_09229_, _09187_, word_in[3]);
  nand _41613_ (_09230_, _09189_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nand _41614_ (_09231_, _09230_, _09229_);
  nand _41615_ (_09232_, _09231_, _09186_);
  nand _41616_ (_09233_, _09185_, word_in[11]);
  nand _41617_ (_09234_, _09233_, _09232_);
  nand _41618_ (_09235_, _09234_, _09196_);
  nand _41619_ (_09236_, _09195_, word_in[19]);
  nand _41620_ (_09237_, _09236_, _09235_);
  nand _41621_ (_09238_, _09237_, _09184_);
  nand _41622_ (_09240_, _09182_, _08235_);
  nand _41623_ (_28164_, _09240_, _09238_);
  nand _41624_ (_09241_, _09187_, word_in[4]);
  nand _41625_ (_09242_, _09189_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nand _41626_ (_09243_, _09242_, _09241_);
  nand _41627_ (_09244_, _09243_, _09186_);
  nand _41628_ (_09245_, _09185_, word_in[12]);
  nand _41629_ (_09246_, _09245_, _09244_);
  nand _41630_ (_09247_, _09246_, _09196_);
  nand _41631_ (_09248_, _09195_, word_in[20]);
  nand _41632_ (_09249_, _09248_, _09247_);
  nand _41633_ (_09250_, _09249_, _09184_);
  nand _41634_ (_09251_, _09182_, _08084_);
  nand _41635_ (_28165_, _09251_, _09250_);
  nor _41636_ (_09253_, _09187_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _41637_ (_09254_, _09189_, word_in[5]);
  nor _41638_ (_09255_, _09254_, _09253_);
  nor _41639_ (_09256_, _09255_, _09185_);
  nor _41640_ (_09257_, _09186_, word_in[13]);
  nor _41641_ (_09258_, _09257_, _09256_);
  nand _41642_ (_09259_, _09258_, _09215_);
  nand _41643_ (_09260_, _09224_, word_in[21]);
  nand _41644_ (_09262_, _09260_, _09259_);
  nor _41645_ (_09264_, _09262_, _09182_);
  nor _41646_ (_09265_, _09184_, _08102_);
  nor _41647_ (_28166_, _09265_, _09264_);
  nor _41648_ (_09267_, _09187_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _41649_ (_09268_, _09189_, word_in[6]);
  nor _41650_ (_09269_, _09268_, _09267_);
  nor _41651_ (_09270_, _09269_, _09185_);
  nor _41652_ (_09271_, _09186_, word_in[14]);
  nor _41653_ (_09272_, _09271_, _09270_);
  nor _41654_ (_09273_, _09272_, _09195_);
  nor _41655_ (_09274_, _09196_, word_in[22]);
  nor _41656_ (_09275_, _09274_, _09273_);
  nand _41657_ (_09276_, _09275_, _09184_);
  nand _41658_ (_09278_, _09182_, _08283_);
  nand _41659_ (_28167_, _09278_, _09276_);
  nand _41660_ (_09279_, _09187_, word_in[7]);
  nand _41661_ (_09280_, _09189_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _41662_ (_09281_, _09280_, _09279_);
  nand _41663_ (_09282_, _09281_, _09186_);
  nand _41664_ (_09283_, _09185_, word_in[15]);
  nand _41665_ (_09284_, _09283_, _09282_);
  nand _41666_ (_09285_, _09284_, _09196_);
  nand _41667_ (_09286_, _09224_, word_in[23]);
  nand _41668_ (_09287_, _09286_, _09285_);
  nand _41669_ (_09288_, _09287_, _09184_);
  nand _41670_ (_09289_, _09182_, _07408_);
  nand _41671_ (_28168_, _09289_, _09288_);
  nand _41672_ (_09290_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  nand _41673_ (_09291_, _25052_, _24830_);
  nand _41674_ (_02744_, _09291_, _09290_);
  nand _41675_ (_09292_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  nand _41676_ (_09293_, _01216_, _24830_);
  nand _41677_ (_02751_, _09293_, _09292_);
  nor _41678_ (_09294_, _08175_, _07169_);
  not _41679_ (_09295_, _09294_);
  nor _41680_ (_09296_, _08179_, _07038_);
  nor _41681_ (_09297_, _07797_, _07376_);
  not _41682_ (_09298_, _09297_);
  nor _41683_ (_09299_, _09298_, _08182_);
  not _41684_ (_09300_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _41685_ (_09301_, _09297_, _09300_);
  nor _41686_ (_09302_, _09301_, _09299_);
  nor _41687_ (_09303_, _09302_, _09296_);
  not _41688_ (_09304_, _09296_);
  nor _41689_ (_09306_, _09304_, _08027_);
  nor _41690_ (_09307_, _09306_, _09303_);
  nand _41691_ (_09308_, _09307_, _09295_);
  nor _41692_ (_09309_, _09181_, _06925_);
  nor _41693_ (_09310_, _09295_, _08694_);
  nor _41694_ (_09311_, _09310_, _09309_);
  nand _41695_ (_09312_, _09311_, _09308_);
  nand _41696_ (_09313_, _09309_, _08699_);
  nand _41697_ (_28180_[0], _09313_, _09312_);
  nor _41698_ (_09314_, _04173_, _25028_);
  nand _41699_ (_09315_, _04193_, _04176_);
  nand _41700_ (_09317_, _09315_, _07744_);
  nor _41701_ (_09318_, _09317_, _07747_);
  nor _41702_ (_09319_, _04188_, _01587_);
  not _41703_ (_09320_, _09319_);
  nor _41704_ (_09321_, _09320_, _01594_);
  nand _41705_ (_09322_, _09321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _41706_ (_09323_, _09322_, _04176_);
  nand _41707_ (_09324_, _09323_, _07739_);
  nor _41708_ (_09325_, _04191_, _01625_);
  nand _41709_ (_09326_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _41710_ (_09327_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _41711_ (_09328_, _09327_, _01616_);
  nand _41712_ (_09329_, _09328_, _09326_);
  nand _41713_ (_09330_, _09329_, _09324_);
  nor _41714_ (_09331_, _09330_, _09318_);
  nand _41715_ (_09332_, _09331_, _04173_);
  nand _41716_ (_09333_, _09332_, _04175_);
  nor _41717_ (_09334_, _09333_, _09314_);
  nor _41718_ (_09335_, _04175_, _04176_);
  nor _41719_ (_09336_, _09335_, _09334_);
  nor _41720_ (_02759_, _09336_, rst);
  nor _41721_ (_09337_, _09297_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _41722_ (_09338_, _09298_, word_in[1]);
  nor _41723_ (_09339_, _09338_, _09337_);
  nor _41724_ (_09340_, _09339_, _09296_);
  nor _41725_ (_09341_, _09304_, word_in[9]);
  nor _41726_ (_09342_, _09341_, _09340_);
  nor _41727_ (_09343_, _09342_, _09294_);
  nor _41728_ (_09344_, _09295_, _08402_);
  nor _41729_ (_09345_, _09344_, _09343_);
  nor _41730_ (_09347_, _09345_, _09309_);
  not _41731_ (_09348_, _09309_);
  nor _41732_ (_09349_, _09348_, _08038_);
  nor _41733_ (_28180_[1], _09349_, _09347_);
  nand _41734_ (_09351_, _09294_, _08719_);
  nand _41735_ (_09352_, _09297_, word_in[2]);
  nand _41736_ (_09353_, _09298_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand _41737_ (_09354_, _09353_, _09352_);
  nand _41738_ (_09355_, _09354_, _09304_);
  nand _41739_ (_09356_, _09296_, word_in[10]);
  nand _41740_ (_09357_, _09356_, _09355_);
  nand _41741_ (_09358_, _09357_, _09295_);
  nand _41742_ (_09359_, _09358_, _09351_);
  nand _41743_ (_09361_, _09359_, _09348_);
  nand _41744_ (_09362_, _09309_, _08054_);
  nand _41745_ (_28180_[2], _09362_, _09361_);
  nand _41746_ (_09363_, _01217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  nand _41747_ (_09364_, _01216_, _25203_);
  nand _41748_ (_02763_, _09364_, _09363_);
  not _41749_ (_09365_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nand _41750_ (_09366_, _09298_, _09365_);
  nand _41751_ (_09367_, _09297_, _08737_);
  nand _41752_ (_09368_, _09367_, _09366_);
  nand _41753_ (_09369_, _09368_, _09304_);
  nand _41754_ (_09370_, _09296_, _08243_);
  nand _41755_ (_09371_, _09370_, _09369_);
  nand _41756_ (_09372_, _09371_, _09295_);
  nor _41757_ (_09373_, _09295_, _08248_);
  nor _41758_ (_09374_, _09373_, _09309_);
  nand _41759_ (_09375_, _09374_, _09372_);
  nand _41760_ (_09376_, _09309_, _08235_);
  nand _41761_ (_28180_[3], _09376_, _09375_);
  nand _41762_ (_09377_, _09294_, _08763_);
  nand _41763_ (_09378_, _09298_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nand _41764_ (_09379_, _09297_, _08254_);
  nand _41765_ (_09380_, _09379_, _09378_);
  nand _41766_ (_09381_, _09380_, _09304_);
  nand _41767_ (_09382_, _09296_, word_in[12]);
  nand _41768_ (_09383_, _09382_, _09381_);
  nand _41769_ (_09384_, _09383_, _09295_);
  nand _41770_ (_09385_, _09384_, _09377_);
  nand _41771_ (_09386_, _09385_, _09348_);
  nand _41772_ (_09387_, _09309_, _08084_);
  nand _41773_ (_28180_[4], _09387_, _09386_);
  nand _41774_ (_09388_, _09294_, _08613_);
  nand _41775_ (_09389_, _09297_, word_in[5]);
  nand _41776_ (_09390_, _09298_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nand _41777_ (_09391_, _09390_, _09389_);
  nand _41778_ (_09392_, _09391_, _09304_);
  nand _41779_ (_09393_, _09296_, word_in[13]);
  nand _41780_ (_09394_, _09393_, _09392_);
  nand _41781_ (_09395_, _09394_, _09295_);
  nand _41782_ (_09396_, _09395_, _09388_);
  nand _41783_ (_09397_, _09396_, _09348_);
  nand _41784_ (_09398_, _09309_, _08102_);
  nand _41785_ (_28180_[5], _09398_, _09397_);
  nand _41786_ (_09399_, _09294_, _08298_);
  nand _41787_ (_09400_, _09297_, word_in[6]);
  nand _41788_ (_09401_, _09298_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nand _41789_ (_09402_, _09401_, _09400_);
  nand _41790_ (_09403_, _09402_, _09304_);
  nand _41791_ (_09404_, _09296_, word_in[14]);
  nand _41792_ (_09405_, _09404_, _09403_);
  nand _41793_ (_09406_, _09405_, _09295_);
  nand _41794_ (_09407_, _09406_, _09399_);
  nand _41795_ (_09408_, _09407_, _09348_);
  nand _41796_ (_09409_, _09309_, _08283_);
  nand _41797_ (_28180_[6], _09409_, _09408_);
  nand _41798_ (_09410_, _09297_, word_in[7]);
  nand _41799_ (_09411_, _09298_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _41800_ (_09412_, _09411_, _09410_);
  nor _41801_ (_09414_, _09412_, _09296_);
  nand _41802_ (_09415_, _09296_, _07387_);
  nand _41803_ (_09416_, _09415_, _09295_);
  nor _41804_ (_09417_, _09416_, _09414_);
  nand _41805_ (_09418_, _09294_, _07400_);
  nand _41806_ (_09420_, _09418_, _09348_);
  nor _41807_ (_09421_, _09420_, _09417_);
  nor _41808_ (_09422_, _09348_, _07408_);
  nor _41809_ (_28180_[7], _09422_, _09421_);
  nand _41810_ (_09423_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nand _41811_ (_09424_, _25052_, _25039_);
  nand _41812_ (_02774_, _09424_, _09423_);
  nand _41813_ (_09425_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  nand _41814_ (_09426_, _28096_, _25052_);
  nand _41815_ (_02780_, _09426_, _09425_);
  nand _41816_ (_09427_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  nand _41817_ (_09429_, _04264_, _28096_);
  nand _41818_ (_02801_, _09429_, _09427_);
  nand _41819_ (_09430_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  nand _41820_ (_09431_, _04264_, _25150_);
  nand _41821_ (_02805_, _09431_, _09430_);
  nand _41822_ (_09432_, _04265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  nand _41823_ (_09433_, _04264_, _24927_);
  nand _41824_ (_02812_, _09433_, _09432_);
  nor _41825_ (_09434_, _07395_, _07014_);
  not _41826_ (_09435_, _09434_);
  nor _41827_ (_09436_, _08363_, _07169_);
  nand _41828_ (_09437_, _09436_, _08694_);
  not _41829_ (_09438_, _09436_);
  nor _41830_ (_09439_, _08368_, _07038_);
  not _41831_ (_09440_, _09439_);
  nor _41832_ (_09441_, _07783_, _07376_);
  not _41833_ (_09442_, _09441_);
  nand _41834_ (_09443_, _09442_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nand _41835_ (_09444_, _09441_, _08183_);
  nand _41836_ (_09445_, _09444_, _09443_);
  nand _41837_ (_09446_, _09445_, _09440_);
  nand _41838_ (_09447_, _09439_, word_in[8]);
  nand _41839_ (_09448_, _09447_, _09446_);
  nand _41840_ (_09449_, _09448_, _09438_);
  nand _41841_ (_09450_, _09449_, _09437_);
  nand _41842_ (_09451_, _09450_, _09435_);
  nand _41843_ (_09452_, _09434_, word_in[24]);
  nand _41844_ (_28170_[0], _09452_, _09451_);
  nand _41845_ (_09453_, _07810_, _24927_);
  nand _41846_ (_09454_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  nand _41847_ (_02827_, _09454_, _09453_);
  nand _41848_ (_09455_, _09439_, _08046_);
  nand _41849_ (_09456_, _09442_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand _41850_ (_09458_, _09441_, _08200_);
  nand _41851_ (_09459_, _09458_, _09456_);
  nor _41852_ (_09460_, _09459_, _09439_);
  nor _41853_ (_09461_, _09460_, _09436_);
  nand _41854_ (_09462_, _09461_, _09455_);
  nand _41855_ (_09463_, _09436_, _08402_);
  nand _41856_ (_09464_, _09463_, _09462_);
  nand _41857_ (_09465_, _09464_, _09435_);
  nand _41858_ (_09466_, _09434_, word_in[25]);
  nand _41859_ (_28170_[1], _09466_, _09465_);
  nand _41860_ (_09467_, _09436_, _08719_);
  nand _41861_ (_09468_, _09442_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand _41862_ (_09469_, _09441_, _08218_);
  nand _41863_ (_09470_, _09469_, _09468_);
  nand _41864_ (_09472_, _09470_, _09440_);
  nand _41865_ (_09473_, _09439_, word_in[10]);
  nand _41866_ (_09475_, _09473_, _09472_);
  nand _41867_ (_09476_, _09475_, _09438_);
  nand _41868_ (_09477_, _09476_, _09467_);
  nand _41869_ (_09478_, _09477_, _09435_);
  nand _41870_ (_09480_, _09434_, word_in[26]);
  nand _41871_ (_28170_[2], _09480_, _09478_);
  nor _41872_ (_09481_, _09441_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _41873_ (_09482_, _09442_, word_in[3]);
  nor _41874_ (_09483_, _09482_, _09481_);
  nor _41875_ (_09484_, _09483_, _09439_);
  nand _41876_ (_09485_, _09439_, _08243_);
  nand _41877_ (_09486_, _09485_, _09438_);
  nor _41878_ (_09487_, _09486_, _09484_);
  nand _41879_ (_09488_, _09436_, _08248_);
  nand _41880_ (_09489_, _09488_, _09435_);
  nor _41881_ (_09490_, _09489_, _09487_);
  nor _41882_ (_09491_, _09435_, word_in[27]);
  nor _41883_ (_28170_[3], _09491_, _09490_);
  nand _41884_ (_09492_, _09436_, _08763_);
  nand _41885_ (_09493_, _09442_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nand _41886_ (_09494_, _09441_, _08254_);
  nand _41887_ (_09495_, _09494_, _09493_);
  nand _41888_ (_09496_, _09495_, _09440_);
  nand _41889_ (_09497_, _09439_, word_in[12]);
  nand _41890_ (_09498_, _09497_, _09496_);
  nand _41891_ (_09499_, _09498_, _09438_);
  nand _41892_ (_09500_, _09499_, _09492_);
  nand _41893_ (_09501_, _09500_, _09435_);
  nand _41894_ (_09503_, _09434_, word_in[28]);
  nand _41895_ (_28170_[4], _09503_, _09501_);
  nand _41896_ (_09504_, _08653_, _28096_);
  nand _41897_ (_09505_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nand _41898_ (_02834_, _09505_, _09504_);
  nor _41899_ (_09506_, _09442_, _08106_);
  not _41900_ (_09507_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _41901_ (_09508_, _09441_, _09507_);
  nor _41902_ (_09509_, _09508_, _09506_);
  nor _41903_ (_09510_, _09509_, _09439_);
  nor _41904_ (_09511_, _09440_, _08110_);
  nor _41905_ (_09512_, _09511_, _09510_);
  nor _41906_ (_09513_, _09512_, _09436_);
  nand _41907_ (_09514_, _09436_, _08613_);
  nand _41908_ (_09515_, _09514_, _09435_);
  nor _41909_ (_09516_, _09515_, _09513_);
  nor _41910_ (_09517_, _09435_, _08102_);
  nor _41911_ (_28170_[5], _09517_, _09516_);
  nand _41912_ (_09518_, _09436_, _08298_);
  nand _41913_ (_09519_, _09441_, word_in[6]);
  nand _41914_ (_09520_, _09442_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nand _41915_ (_09521_, _09520_, _09519_);
  nand _41916_ (_09522_, _09521_, _09440_);
  nand _41917_ (_09523_, _09439_, word_in[14]);
  nand _41918_ (_09524_, _09523_, _09522_);
  nand _41919_ (_09525_, _09524_, _09438_);
  nand _41920_ (_09526_, _09525_, _09518_);
  nand _41921_ (_09527_, _09526_, _09435_);
  nand _41922_ (_09528_, _09434_, word_in[30]);
  nand _41923_ (_28170_[6], _09528_, _09527_);
  nand _41924_ (_09530_, _09442_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _41925_ (_09531_, _09441_, _08306_);
  nand _41926_ (_09532_, _09531_, _09530_);
  nor _41927_ (_09533_, _09532_, _09439_);
  nand _41928_ (_09534_, _09439_, _07387_);
  nand _41929_ (_09535_, _09534_, _09438_);
  nor _41930_ (_09536_, _09535_, _09533_);
  nand _41931_ (_09537_, _09436_, _07400_);
  nand _41932_ (_09538_, _09537_, _09435_);
  nor _41933_ (_09539_, _09538_, _09536_);
  nor _41934_ (_09540_, _09435_, _07408_);
  nor _41935_ (_28170_[7], _09540_, _09539_);
  nand _41936_ (_09541_, _08653_, _25150_);
  nand _41937_ (_09542_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  nand _41938_ (_02848_, _09542_, _09541_);
  nand _41939_ (_09543_, _08653_, _25039_);
  nand _41940_ (_09545_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  nand _41941_ (_02855_, _09545_, _09543_);
  nor _41942_ (_09547_, _28104_, _24059_);
  nand _41943_ (_09548_, _09547_, _28096_);
  not _41944_ (_09549_, _09547_);
  nand _41945_ (_09550_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  nand _41946_ (_02869_, _09550_, _09548_);
  nand _41947_ (_09551_, _28105_, _24830_);
  nand _41948_ (_09552_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  nand _41949_ (_02874_, _09552_, _09551_);
  nand _41950_ (_09553_, _09547_, _24789_);
  nand _41951_ (_09554_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  nand _41952_ (_02877_, _09554_, _09553_);
  nand _41953_ (_09555_, _28105_, _25039_);
  nand _41954_ (_09556_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nand _41955_ (_02885_, _09556_, _09555_);
  nand _41956_ (_09557_, _28105_, _25203_);
  nand _41957_ (_09558_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  nand _41958_ (_02890_, _09558_, _09557_);
  nor _41959_ (_09559_, _07716_, _07393_);
  not _41960_ (_09560_, _09559_);
  nor _41961_ (_09561_, _08517_, _07169_);
  nand _41962_ (_09562_, _09561_, _08694_);
  not _41963_ (_09563_, _09561_);
  nor _41964_ (_09564_, _08506_, _07038_);
  not _41965_ (_09565_, _09564_);
  not _41966_ (_09566_, _07832_);
  nor _41967_ (_09567_, _09566_, _07376_);
  not _41968_ (_09568_, _09567_);
  nand _41969_ (_09569_, _09568_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nand _41970_ (_09570_, _09567_, _08183_);
  nand _41971_ (_09571_, _09570_, _09569_);
  nand _41972_ (_09572_, _09571_, _09565_);
  nand _41973_ (_09573_, _09564_, word_in[8]);
  nand _41974_ (_09574_, _09573_, _09572_);
  nand _41975_ (_09575_, _09574_, _09563_);
  nand _41976_ (_09576_, _09575_, _09562_);
  nand _41977_ (_09577_, _09576_, _09560_);
  nand _41978_ (_09579_, _09559_, word_in[24]);
  nand _41979_ (_28136_, _09579_, _09577_);
  nand _41980_ (_09580_, _28105_, _25150_);
  nand _41981_ (_09581_, _28107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  nand _41982_ (_02898_, _09581_, _09580_);
  nand _41983_ (_09582_, _09564_, _08046_);
  nand _41984_ (_09583_, _09568_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nand _41985_ (_09584_, _09567_, _08200_);
  nand _41986_ (_09585_, _09584_, _09583_);
  nor _41987_ (_09586_, _09585_, _09564_);
  nor _41988_ (_09587_, _09586_, _09561_);
  nand _41989_ (_09588_, _09587_, _09582_);
  nand _41990_ (_09589_, _09561_, _08402_);
  nand _41991_ (_09590_, _09589_, _09588_);
  nand _41992_ (_09591_, _09590_, _09560_);
  nand _41993_ (_09592_, _09559_, word_in[25]);
  nand _41994_ (_28137_, _09592_, _09591_);
  nand _41995_ (_09593_, _09561_, _08719_);
  nand _41996_ (_09594_, _09567_, word_in[2]);
  nand _41997_ (_09595_, _09568_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nand _41998_ (_09596_, _09595_, _09594_);
  nand _41999_ (_09597_, _09596_, _09565_);
  nand _42000_ (_09598_, _09564_, word_in[10]);
  nand _42001_ (_09599_, _09598_, _09597_);
  nand _42002_ (_09600_, _09599_, _09563_);
  nand _42003_ (_09601_, _09600_, _09593_);
  nand _42004_ (_09602_, _09601_, _09560_);
  nand _42005_ (_09603_, _09559_, word_in[26]);
  nand _42006_ (_28138_, _09603_, _09602_);
  nand _42007_ (_09604_, _08806_, _25039_);
  nand _42008_ (_09605_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  nand _42009_ (_02903_, _09605_, _09604_);
  nand _42010_ (_09606_, _09561_, _08248_);
  nand _42011_ (_09607_, _09567_, word_in[3]);
  nand _42012_ (_09608_, _09568_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nand _42013_ (_09609_, _09608_, _09607_);
  nand _42014_ (_09610_, _09609_, _09565_);
  nand _42015_ (_09611_, _09564_, word_in[11]);
  nand _42016_ (_09612_, _09611_, _09610_);
  nand _42017_ (_09613_, _09612_, _09563_);
  nand _42018_ (_09614_, _09613_, _09606_);
  nand _42019_ (_09615_, _09614_, _09560_);
  nand _42020_ (_09616_, _09559_, word_in[27]);
  nand _42021_ (_28139_, _09616_, _09615_);
  nand _42022_ (_09617_, _09564_, _08092_);
  nand _42023_ (_09618_, _09568_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nand _42024_ (_09619_, _09567_, _08254_);
  nand _42025_ (_09620_, _09619_, _09618_);
  nor _42026_ (_09622_, _09620_, _09564_);
  nor _42027_ (_09623_, _09622_, _09561_);
  nand _42028_ (_09624_, _09623_, _09617_);
  nand _42029_ (_09625_, _09561_, _08763_);
  nand _42030_ (_09626_, _09625_, _09624_);
  nand _42031_ (_09627_, _09626_, _09560_);
  nand _42032_ (_09628_, _09559_, word_in[28]);
  nand _42033_ (_28140_, _09628_, _09627_);
  nand _42034_ (_09629_, _09561_, _08613_);
  nand _42035_ (_09630_, _09567_, word_in[5]);
  nand _42036_ (_09631_, _09568_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nand _42037_ (_09632_, _09631_, _09630_);
  nand _42038_ (_09633_, _09632_, _09565_);
  nand _42039_ (_09634_, _09564_, word_in[13]);
  nand _42040_ (_09635_, _09634_, _09633_);
  nand _42041_ (_09637_, _09635_, _09563_);
  nand _42042_ (_09639_, _09637_, _09629_);
  nand _42043_ (_09640_, _09639_, _09560_);
  nand _42044_ (_09642_, _09559_, word_in[29]);
  nand _42045_ (_28141_, _09642_, _09640_);
  not _42046_ (_09644_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nand _42047_ (_09645_, _09568_, _09644_);
  nand _42048_ (_09647_, _09567_, _08618_);
  nand _42049_ (_09649_, _09647_, _09645_);
  nand _42050_ (_09652_, _09649_, _09565_);
  nand _42051_ (_09653_, _09564_, _08293_);
  nand _42052_ (_09654_, _09653_, _09652_);
  nand _42053_ (_09655_, _09654_, _09563_);
  nor _42054_ (_09656_, _09563_, _08298_);
  nor _42055_ (_09657_, _09656_, _09559_);
  nand _42056_ (_09658_, _09657_, _09655_);
  nand _42057_ (_09659_, _09559_, word_in[30]);
  nand _42058_ (_28142_, _09659_, _09658_);
  nand _42059_ (_09660_, _09564_, _07387_);
  nand _42060_ (_09661_, _09568_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _42061_ (_09662_, _09567_, _08306_);
  nand _42062_ (_09663_, _09662_, _09661_);
  nor _42063_ (_09664_, _09663_, _09564_);
  nor _42064_ (_09665_, _09664_, _09561_);
  nand _42065_ (_09666_, _09665_, _09660_);
  nand _42066_ (_09668_, _09561_, _07400_);
  nand _42067_ (_09669_, _09668_, _09666_);
  nand _42068_ (_09670_, _09669_, _09560_);
  nand _42069_ (_09671_, _09559_, word_in[31]);
  nand _42070_ (_28143_, _09671_, _09670_);
  nand _42071_ (_09672_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nand _42072_ (_09673_, _04601_, _25039_);
  nand _42073_ (_02925_, _09673_, _09672_);
  nand _42074_ (_09674_, _03442_, _25039_);
  nand _42075_ (_09675_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nand _42076_ (_02944_, _09675_, _09674_);
  nand _42077_ (_09676_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nand _42078_ (_09677_, _04021_, _25039_);
  nand _42079_ (_02958_, _09677_, _09676_);
  nor _42080_ (_09678_, _07398_, _06886_);
  not _42081_ (_09679_, _09678_);
  nor _42082_ (_09680_, _07363_, _06925_);
  nand _42083_ (_09681_, _09680_, word_in[16]);
  not _42084_ (_09682_, _09680_);
  nor _42085_ (_09684_, _09566_, _07367_);
  not _42086_ (_09685_, _09684_);
  nor _42087_ (_09686_, _06907_, _06867_);
  nand _42088_ (_09687_, _09686_, _07375_);
  not _42089_ (_09688_, _09687_);
  nand _42090_ (_09689_, _09688_, word_in[0]);
  nand _42091_ (_09690_, _09687_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nand _42092_ (_09692_, _09690_, _09689_);
  nand _42093_ (_09694_, _09692_, _09685_);
  nand _42094_ (_09696_, _09684_, _08028_);
  nand _42095_ (_09697_, _09696_, _09694_);
  nand _42096_ (_09698_, _09697_, _09682_);
  nand _42097_ (_09699_, _09698_, _09681_);
  nand _42098_ (_09700_, _09699_, _09679_);
  nand _42099_ (_09701_, _09678_, word_in[24]);
  nand _42100_ (_28171_[0], _09701_, _09700_);
  nand _42101_ (_09703_, _09688_, word_in[1]);
  nand _42102_ (_09704_, _09687_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nand _42103_ (_09705_, _09704_, _09703_);
  nand _42104_ (_09706_, _09705_, _09685_);
  nor _42105_ (_09708_, _07367_, _08046_);
  nand _42106_ (_09709_, _09684_, _09708_);
  nand _42107_ (_09710_, _09709_, _09706_);
  nand _42108_ (_09711_, _09710_, _09682_);
  nand _42109_ (_09712_, _09680_, word_in[17]);
  nand _42110_ (_09713_, _09712_, _09711_);
  nand _42111_ (_09715_, _09713_, _09679_);
  nand _42112_ (_09716_, _09678_, word_in[25]);
  nand _42113_ (_28171_[1], _09716_, _09715_);
  nor _42114_ (_09717_, _09688_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _42115_ (_09718_, _09687_, word_in[2]);
  nor _42116_ (_09719_, _09718_, _09717_);
  nor _42117_ (_09720_, _09719_, _09684_);
  nor _42118_ (_09721_, _07367_, _08064_);
  nor _42119_ (_09722_, _09685_, _09721_);
  nor _42120_ (_09723_, _09722_, _09720_);
  nor _42121_ (_09724_, _09723_, _09680_);
  nor _42122_ (_09726_, _09682_, word_in[18]);
  nor _42123_ (_09727_, _09726_, _09724_);
  nor _42124_ (_09729_, _09727_, _09678_);
  nor _42125_ (_09730_, _09679_, word_in[26]);
  nor _42126_ (_28171_[2], _09730_, _09729_);
  nor _42127_ (_09731_, _09688_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _42128_ (_09733_, _09687_, word_in[3]);
  nor _42129_ (_09734_, _09733_, _09731_);
  nor _42130_ (_09735_, _09734_, _09684_);
  nor _42131_ (_09736_, _07367_, _08243_);
  nor _42132_ (_09737_, _09685_, _09736_);
  nor _42133_ (_09738_, _09737_, _09735_);
  nor _42134_ (_09739_, _09738_, _09680_);
  nor _42135_ (_09740_, _09682_, word_in[19]);
  nor _42136_ (_09741_, _09740_, _09739_);
  nor _42137_ (_09743_, _09741_, _09678_);
  nor _42138_ (_09744_, _09679_, word_in[27]);
  nor _42139_ (_28171_[3], _09744_, _09743_);
  nand _42140_ (_09745_, _09688_, word_in[4]);
  nand _42141_ (_09746_, _09687_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand _42142_ (_09747_, _09746_, _09745_);
  nand _42143_ (_09748_, _09747_, _09685_);
  nor _42144_ (_09749_, _07367_, _08092_);
  nand _42145_ (_09750_, _09684_, _09749_);
  nand _42146_ (_09751_, _09750_, _09748_);
  nand _42147_ (_09752_, _09751_, _09682_);
  nand _42148_ (_09753_, _09680_, word_in[20]);
  nand _42149_ (_09754_, _09753_, _09752_);
  nand _42150_ (_09755_, _09754_, _09679_);
  nand _42151_ (_09756_, _09678_, word_in[28]);
  nand _42152_ (_28171_[4], _09756_, _09755_);
  nand _42153_ (_09757_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nand _42154_ (_09758_, _04610_, _25203_);
  nand _42155_ (_02970_, _09758_, _09757_);
  nand _42156_ (_09760_, _09688_, word_in[5]);
  nand _42157_ (_09761_, _09687_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nand _42158_ (_09762_, _09761_, _09760_);
  nand _42159_ (_09763_, _09762_, _09685_);
  nor _42160_ (_09764_, _07367_, _08110_);
  nand _42161_ (_09765_, _09684_, _09764_);
  nand _42162_ (_09766_, _09765_, _09763_);
  nand _42163_ (_09767_, _09766_, _09682_);
  nand _42164_ (_09768_, _09680_, word_in[21]);
  nand _42165_ (_09769_, _09768_, _09767_);
  nand _42166_ (_09771_, _09769_, _09679_);
  nand _42167_ (_09772_, _09678_, word_in[29]);
  nand _42168_ (_28171_[5], _09772_, _09771_);
  nor _42169_ (_09773_, _09688_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _42170_ (_09775_, _09687_, word_in[6]);
  nor _42171_ (_09776_, _09775_, _09773_);
  nor _42172_ (_09778_, _09776_, _09684_);
  nor _42173_ (_09779_, _07367_, _08293_);
  nor _42174_ (_09780_, _09685_, _09779_);
  nor _42175_ (_09782_, _09780_, _09778_);
  nor _42176_ (_09783_, _09782_, _09680_);
  nor _42177_ (_09784_, _09682_, word_in[22]);
  nor _42178_ (_09785_, _09784_, _09783_);
  nand _42179_ (_09786_, _09785_, _09679_);
  nand _42180_ (_09787_, _09678_, _08283_);
  nand _42181_ (_28171_[6], _09787_, _09786_);
  not _42182_ (_09788_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _42183_ (_09789_, _09688_, _09788_);
  nor _42184_ (_09790_, _09687_, _07381_);
  nor _42185_ (_09792_, _09790_, _09789_);
  nand _42186_ (_09793_, _09792_, _09685_);
  nor _42187_ (_09794_, _07367_, _07387_);
  nor _42188_ (_09795_, _09685_, _09794_);
  nor _42189_ (_09796_, _09795_, _09680_);
  nand _42190_ (_09797_, _09796_, _09793_);
  nand _42191_ (_09798_, _09680_, _07400_);
  nand _42192_ (_09799_, _09798_, _09797_);
  nand _42193_ (_09800_, _09799_, _09679_);
  nand _42194_ (_09802_, _09678_, word_in[31]);
  nand _42195_ (_28171_[7], _09802_, _09800_);
  nand _42196_ (_09803_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  nand _42197_ (_09804_, _04021_, _24927_);
  nand _42198_ (_02978_, _09804_, _09803_);
  nand _42199_ (_09807_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nand _42200_ (_09808_, _28074_, _25039_);
  nand _42201_ (_02983_, _09808_, _09807_);
  nand _42202_ (_09810_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  nand _42203_ (_09811_, _28096_, _28074_);
  nand _42204_ (_02989_, _09811_, _09810_);
  nand _42205_ (_09812_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nand _42206_ (_09813_, _04015_, _25099_);
  nand _42207_ (_02998_, _09813_, _09812_);
  nand _42208_ (_09815_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  nand _42209_ (_09816_, _28074_, _24789_);
  nand _42210_ (_03002_, _09816_, _09815_);
  nand _42211_ (_09818_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nand _42212_ (_09819_, _04015_, _24789_);
  nand _42213_ (_03007_, _09819_, _09818_);
  nand _42214_ (_09821_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  nand _42215_ (_09822_, _04015_, _25039_);
  nand _42216_ (_03010_, _09822_, _09821_);
  nor _42217_ (_09823_, _07398_, _06925_);
  not _42218_ (_09824_, _09823_);
  nor _42219_ (_09825_, _08175_, _07357_);
  nand _42220_ (_09826_, _09825_, word_in[16]);
  not _42221_ (_09827_, _09825_);
  nor _42222_ (_09828_, _07369_, _06907_);
  not _42223_ (_09830_, _09828_);
  nand _42224_ (_09832_, _07893_, _07375_);
  not _42225_ (_09833_, _09832_);
  nand _42226_ (_09834_, _09833_, word_in[0]);
  nand _42227_ (_09835_, _09832_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nand _42228_ (_09836_, _09835_, _09834_);
  nand _42229_ (_09837_, _09836_, _09830_);
  nand _42230_ (_09839_, _09828_, _08028_);
  nand _42231_ (_09840_, _09839_, _09837_);
  nand _42232_ (_09841_, _09840_, _09827_);
  nand _42233_ (_09842_, _09841_, _09826_);
  nand _42234_ (_09843_, _09842_, _09824_);
  nand _42235_ (_09844_, _09823_, _08699_);
  nand _42236_ (_28172_[0], _09844_, _09843_);
  nand _42237_ (_09845_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nand _42238_ (_09846_, _08334_, _24830_);
  nand _42239_ (_03027_, _09846_, _09845_);
  nand _42240_ (_09847_, _09833_, word_in[1]);
  nand _42241_ (_09848_, _09832_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nand _42242_ (_09850_, _09848_, _09847_);
  nand _42243_ (_09851_, _09850_, _09830_);
  nand _42244_ (_09852_, _09828_, _09708_);
  nand _42245_ (_09853_, _09852_, _09851_);
  nand _42246_ (_09854_, _09853_, _09827_);
  nand _42247_ (_09856_, _09825_, word_in[17]);
  nand _42248_ (_09857_, _09856_, _09854_);
  nand _42249_ (_09858_, _09857_, _09824_);
  nand _42250_ (_09859_, _09823_, _08038_);
  nand _42251_ (_28172_[1], _09859_, _09858_);
  nor _42252_ (_09860_, _09833_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _42253_ (_09862_, _09832_, word_in[2]);
  nor _42254_ (_09863_, _09862_, _09860_);
  nor _42255_ (_09865_, _09863_, _09828_);
  nor _42256_ (_09866_, _09830_, _09721_);
  nor _42257_ (_09867_, _09866_, _09865_);
  nor _42258_ (_09868_, _09867_, _09825_);
  nor _42259_ (_09869_, _09827_, word_in[18]);
  nor _42260_ (_09870_, _09869_, _09868_);
  nor _42261_ (_09871_, _09870_, _09823_);
  nor _42262_ (_09872_, _09824_, _08054_);
  nor _42263_ (_28172_[2], _09872_, _09871_);
  nand _42264_ (_09873_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nand _42265_ (_09874_, _08549_, _25099_);
  nand _42266_ (_03030_, _09874_, _09873_);
  nand _42267_ (_09875_, _09833_, word_in[3]);
  nand _42268_ (_09877_, _09832_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nand _42269_ (_09878_, _09877_, _09875_);
  nand _42270_ (_09879_, _09878_, _09830_);
  nand _42271_ (_09880_, _09828_, _09736_);
  nand _42272_ (_09881_, _09880_, _09879_);
  nand _42273_ (_09882_, _09881_, _09827_);
  nand _42274_ (_09883_, _09825_, word_in[19]);
  nand _42275_ (_09884_, _09883_, _09882_);
  nand _42276_ (_09885_, _09884_, _09824_);
  nand _42277_ (_09886_, _09823_, _08235_);
  nand _42278_ (_28172_[3], _09886_, _09885_);
  nor _42279_ (_09888_, _09833_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _42280_ (_09890_, _09832_, word_in[4]);
  nor _42281_ (_09891_, _09890_, _09888_);
  nor _42282_ (_09892_, _09891_, _09828_);
  nor _42283_ (_09893_, _09830_, _09749_);
  nor _42284_ (_09894_, _09893_, _09892_);
  nor _42285_ (_09895_, _09894_, _09825_);
  nor _42286_ (_09896_, _09827_, word_in[20]);
  nor _42287_ (_09897_, _09896_, _09895_);
  nor _42288_ (_09899_, _09897_, _09823_);
  nor _42289_ (_09901_, _09824_, _08084_);
  nor _42290_ (_28172_[4], _09901_, _09899_);
  nand _42291_ (_09903_, _09833_, word_in[5]);
  nand _42292_ (_09904_, _09832_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nand _42293_ (_09905_, _09904_, _09903_);
  nand _42294_ (_09906_, _09905_, _09830_);
  nand _42295_ (_09907_, _09828_, _09764_);
  nand _42296_ (_09908_, _09907_, _09906_);
  nand _42297_ (_09909_, _09908_, _09827_);
  nand _42298_ (_09910_, _09825_, word_in[21]);
  nand _42299_ (_09912_, _09910_, _09909_);
  nand _42300_ (_09914_, _09912_, _09824_);
  nand _42301_ (_09915_, _09823_, _08102_);
  nand _42302_ (_28172_[5], _09915_, _09914_);
  nor _42303_ (_09916_, _09833_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _42304_ (_09917_, _09832_, word_in[6]);
  nor _42305_ (_09918_, _09917_, _09916_);
  nor _42306_ (_09919_, _09918_, _09828_);
  nor _42307_ (_09920_, _09830_, _09779_);
  nor _42308_ (_09921_, _09920_, _09919_);
  nor _42309_ (_09922_, _09921_, _09825_);
  nor _42310_ (_09923_, _09827_, word_in[22]);
  nor _42311_ (_09924_, _09923_, _09922_);
  nor _42312_ (_09925_, _09924_, _09823_);
  nor _42313_ (_09927_, _09824_, _08283_);
  nor _42314_ (_28172_[6], _09927_, _09925_);
  nor _42315_ (_09928_, _09833_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _42316_ (_09929_, _09832_, word_in[7]);
  nor _42317_ (_09930_, _09929_, _09928_);
  nor _42318_ (_09931_, _09930_, _09828_);
  nor _42319_ (_09932_, _09830_, _09794_);
  nor _42320_ (_09933_, _09932_, _09931_);
  nor _42321_ (_09934_, _09933_, _09825_);
  nor _42322_ (_09936_, _09827_, word_in[23]);
  nor _42323_ (_09937_, _09936_, _09934_);
  nor _42324_ (_09938_, _09937_, _09823_);
  nor _42325_ (_09939_, _09824_, _07408_);
  nor _42326_ (_28172_[7], _09939_, _09938_);
  nand _42327_ (_09940_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  nand _42328_ (_09941_, _08549_, _25150_);
  nand _42329_ (_03042_, _09941_, _09940_);
  nand _42330_ (_09942_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nand _42331_ (_09943_, _08329_, _25150_);
  nand _42332_ (_03046_, _09943_, _09942_);
  nor _42333_ (_09944_, _28057_, _24978_);
  nand _42334_ (_09945_, _09944_, _25150_);
  not _42335_ (_09946_, _09944_);
  nand _42336_ (_09947_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nand _42337_ (_03071_, _09947_, _09945_);
  nand _42338_ (_09949_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nand _42339_ (_09950_, _08319_, _25099_);
  nand _42340_ (_03078_, _09950_, _09949_);
  nor _42341_ (_09951_, _07398_, _07011_);
  not _42342_ (_09952_, _09951_);
  nor _42343_ (_09953_, _08363_, _07357_);
  not _42344_ (_09954_, _09953_);
  nor _42345_ (_09955_, _07369_, _06886_);
  not _42346_ (_09956_, _09955_);
  nor _42347_ (_09957_, _07376_, _08017_);
  nand _42348_ (_09958_, _09957_, word_in[0]);
  not _42349_ (_09959_, _09957_);
  nand _42350_ (_09960_, _09959_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nand _42351_ (_09961_, _09960_, _09958_);
  nand _42352_ (_09962_, _09961_, _09956_);
  nand _42353_ (_09963_, _09955_, _08028_);
  nand _42354_ (_09964_, _09963_, _09962_);
  nand _42355_ (_09966_, _09964_, _09954_);
  nand _42356_ (_09968_, _09953_, word_in[16]);
  nand _42357_ (_09969_, _09968_, _09966_);
  nand _42358_ (_09970_, _09969_, _09952_);
  nand _42359_ (_09971_, _09951_, _08699_);
  nand _42360_ (_28144_, _09971_, _09970_);
  nand _42361_ (_09973_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  nand _42362_ (_09974_, _08501_, _25203_);
  nand _42363_ (_03084_, _09974_, _09973_);
  nor _42364_ (_09975_, _09957_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _42365_ (_09976_, _09959_, word_in[1]);
  nor _42366_ (_09977_, _09976_, _09975_);
  nor _42367_ (_09978_, _09977_, _09955_);
  nor _42368_ (_09979_, _09956_, _09708_);
  nor _42369_ (_09981_, _09979_, _09978_);
  nor _42370_ (_09982_, _09981_, _09953_);
  nor _42371_ (_09983_, _09954_, word_in[17]);
  nor _42372_ (_09984_, _09983_, _09982_);
  nor _42373_ (_09985_, _09984_, _09951_);
  nor _42374_ (_09986_, _09952_, _08038_);
  nor _42375_ (_28145_, _09986_, _09985_);
  nand _42376_ (_09987_, _09957_, word_in[2]);
  nand _42377_ (_09988_, _09959_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand _42378_ (_09989_, _09988_, _09987_);
  nand _42379_ (_09990_, _09989_, _09956_);
  nand _42380_ (_09991_, _09955_, _09721_);
  nand _42381_ (_09993_, _09991_, _09990_);
  nand _42382_ (_09994_, _09993_, _09954_);
  nand _42383_ (_09996_, _09953_, word_in[18]);
  nand _42384_ (_09998_, _09996_, _09994_);
  nand _42385_ (_10000_, _09998_, _09952_);
  nand _42386_ (_10001_, _09951_, _08054_);
  nand _42387_ (_28146_, _10001_, _10000_);
  nand _42388_ (_10003_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nand _42389_ (_10004_, _08501_, _24830_);
  nand _42390_ (_03087_, _10004_, _10003_);
  nand _42391_ (_10006_, _09957_, word_in[3]);
  nand _42392_ (_10008_, _09959_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nand _42393_ (_10009_, _10008_, _10006_);
  nand _42394_ (_10011_, _10009_, _09956_);
  nand _42395_ (_10012_, _09955_, _09736_);
  nand _42396_ (_10013_, _10012_, _10011_);
  nand _42397_ (_10014_, _10013_, _09954_);
  nand _42398_ (_10015_, _09953_, word_in[19]);
  nand _42399_ (_10016_, _10015_, _10014_);
  nand _42400_ (_10017_, _10016_, _09952_);
  nand _42401_ (_10019_, _09951_, _08235_);
  nand _42402_ (_28147_, _10019_, _10017_);
  nor _42403_ (_10021_, _09957_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _42404_ (_10022_, _09959_, word_in[4]);
  nor _42405_ (_10023_, _10022_, _10021_);
  nor _42406_ (_10024_, _10023_, _09955_);
  nor _42407_ (_10025_, _09956_, _09749_);
  nor _42408_ (_10026_, _10025_, _10024_);
  nor _42409_ (_10028_, _10026_, _09953_);
  nor _42410_ (_10029_, _09954_, word_in[20]);
  nor _42411_ (_10030_, _10029_, _10028_);
  nor _42412_ (_10031_, _10030_, _09951_);
  nor _42413_ (_10032_, _09952_, _08084_);
  nor _42414_ (_28148_, _10032_, _10031_);
  nand _42415_ (_10033_, _09953_, word_in[21]);
  nand _42416_ (_10034_, _09957_, word_in[5]);
  nand _42417_ (_10035_, _09959_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nand _42418_ (_10036_, _10035_, _10034_);
  nand _42419_ (_10037_, _10036_, _09956_);
  nand _42420_ (_10038_, _09955_, _09764_);
  nand _42421_ (_10040_, _10038_, _10037_);
  nand _42422_ (_10041_, _10040_, _09954_);
  nand _42423_ (_10042_, _10041_, _10033_);
  nand _42424_ (_10043_, _10042_, _09952_);
  nand _42425_ (_10044_, _09951_, _08102_);
  nand _42426_ (_28149_, _10044_, _10043_);
  nand _42427_ (_10045_, _09957_, word_in[6]);
  nand _42428_ (_10046_, _09959_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nand _42429_ (_10047_, _10046_, _10045_);
  nand _42430_ (_10049_, _10047_, _09956_);
  nand _42431_ (_10050_, _09955_, _09779_);
  nand _42432_ (_10051_, _10050_, _10049_);
  nand _42433_ (_10053_, _10051_, _09954_);
  nand _42434_ (_10054_, _09953_, word_in[22]);
  nand _42435_ (_10055_, _10054_, _10053_);
  nand _42436_ (_10057_, _10055_, _09952_);
  nand _42437_ (_10058_, _09951_, _08283_);
  nand _42438_ (_28150_, _10058_, _10057_);
  nor _42439_ (_10059_, _09957_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nor _42440_ (_10060_, _09959_, word_in[7]);
  nor _42441_ (_10062_, _10060_, _10059_);
  nor _42442_ (_10063_, _10062_, _09955_);
  nor _42443_ (_10064_, _09956_, _09794_);
  nor _42444_ (_10066_, _10064_, _10063_);
  nor _42445_ (_10067_, _10066_, _09953_);
  nor _42446_ (_10068_, _09954_, word_in[23]);
  nor _42447_ (_10069_, _10068_, _10067_);
  nor _42448_ (_10070_, _10069_, _09951_);
  nor _42449_ (_10071_, _09952_, _07408_);
  nor _42450_ (_28151_, _10071_, _10070_);
  nand _42451_ (_10073_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  nand _42452_ (_10074_, _08264_, _24830_);
  nand _42453_ (_03096_, _10074_, _10073_);
  nand _42454_ (_10075_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  nand _42455_ (_10076_, _08230_, _24830_);
  nand _42456_ (_03102_, _10076_, _10075_);
  nand _42457_ (_10077_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nand _42458_ (_10078_, _08230_, _25039_);
  nand _42459_ (_03118_, _10078_, _10077_);
  nand _42460_ (_10081_, _01402_, _24789_);
  nand _42461_ (_10082_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nand _42462_ (_03121_, _10082_, _10081_);
  nor _42463_ (_10084_, _08142_, _00415_);
  not _42464_ (_10085_, _10084_);
  nand _42465_ (_10087_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  nand _42466_ (_10089_, _10084_, _25203_);
  nand _42467_ (_03129_, _10089_, _10087_);
  nand _42468_ (_10090_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nand _42469_ (_10091_, _10084_, _24830_);
  nand _42470_ (_03133_, _10091_, _10090_);
  nor _42471_ (_10092_, _07377_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _42472_ (_10093_, _07378_, word_in[0]);
  nor _42473_ (_10095_, _10093_, _10092_);
  nor _42474_ (_10096_, _10095_, _07370_);
  nor _42475_ (_10097_, _07371_, word_in[8]);
  nor _42476_ (_10098_, _10097_, _10096_);
  nor _42477_ (_10100_, _10098_, _07364_);
  nor _42478_ (_10102_, _07365_, word_in[16]);
  nor _42479_ (_10104_, _10102_, _10100_);
  nor _42480_ (_10105_, _10104_, _07399_);
  not _42481_ (_10107_, _07399_);
  nor _42482_ (_10108_, _08699_, _10107_);
  nor _42483_ (_28173_[0], _10108_, _10105_);
  nor _42484_ (_10110_, _07377_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _42485_ (_10111_, _07378_, word_in[1]);
  nor _42486_ (_10113_, _10111_, _10110_);
  nor _42487_ (_10114_, _10113_, _07370_);
  nor _42488_ (_10115_, _07371_, word_in[9]);
  nor _42489_ (_10117_, _10115_, _10114_);
  nor _42490_ (_10119_, _10117_, _07364_);
  nor _42491_ (_10120_, _07365_, word_in[17]);
  nor _42492_ (_10121_, _10120_, _10119_);
  nor _42493_ (_10122_, _10121_, _07399_);
  nor _42494_ (_10123_, _08038_, _10107_);
  nor _42495_ (_28173_[1], _10123_, _10122_);
  nor _42496_ (_10124_, _07377_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _42497_ (_10125_, _07378_, word_in[2]);
  nor _42498_ (_10126_, _10125_, _10124_);
  nor _42499_ (_10127_, _10126_, _07370_);
  nor _42500_ (_10129_, _07371_, word_in[10]);
  nor _42501_ (_10131_, _10129_, _10127_);
  nor _42502_ (_10133_, _10131_, _07364_);
  nor _42503_ (_10135_, _07365_, word_in[18]);
  nor _42504_ (_10137_, _10135_, _10133_);
  nor _42505_ (_10138_, _10137_, _07399_);
  nor _42506_ (_10140_, _08054_, _10107_);
  nor _42507_ (_28173_[2], _10140_, _10138_);
  nand _42508_ (_10142_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  nand _42509_ (_10144_, _08167_, _24789_);
  nand _42510_ (_03143_, _10144_, _10142_);
  nand _42511_ (_10147_, _07377_, word_in[3]);
  nand _42512_ (_10148_, _07378_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nand _42513_ (_10149_, _10148_, _10147_);
  nand _42514_ (_10150_, _10149_, _07371_);
  nand _42515_ (_10152_, _07370_, word_in[11]);
  nand _42516_ (_10154_, _10152_, _10150_);
  nand _42517_ (_10156_, _10154_, _07365_);
  nand _42518_ (_10157_, _07364_, word_in[19]);
  nand _42519_ (_10158_, _10157_, _10156_);
  nand _42520_ (_10160_, _10158_, _10107_);
  nand _42521_ (_10161_, _08235_, _07399_);
  nand _42522_ (_28173_[3], _10161_, _10160_);
  nand _42523_ (_10162_, _07364_, word_in[20]);
  nand _42524_ (_10163_, _07377_, word_in[4]);
  nand _42525_ (_10165_, _07378_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand _42526_ (_10166_, _10165_, _10163_);
  nand _42527_ (_10167_, _10166_, _07371_);
  nand _42528_ (_10168_, _07370_, word_in[12]);
  nand _42529_ (_10169_, _10168_, _10167_);
  nand _42530_ (_10170_, _10169_, _07365_);
  nand _42531_ (_10171_, _10170_, _10162_);
  nand _42532_ (_10173_, _10171_, _10107_);
  nand _42533_ (_10174_, _08084_, _07399_);
  nand _42534_ (_28173_[4], _10174_, _10173_);
  nand _42535_ (_10175_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nand _42536_ (_10176_, _08167_, _25039_);
  nand _42537_ (_03144_, _10176_, _10175_);
  nand _42538_ (_10177_, _07364_, word_in[21]);
  nand _42539_ (_10178_, _07377_, word_in[5]);
  nand _42540_ (_10179_, _07378_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nand _42541_ (_10180_, _10179_, _10178_);
  nand _42542_ (_10181_, _10180_, _07371_);
  nand _42543_ (_10182_, _07370_, word_in[13]);
  nand _42544_ (_10183_, _10182_, _10181_);
  nand _42545_ (_10184_, _10183_, _07365_);
  nand _42546_ (_10185_, _10184_, _10177_);
  nand _42547_ (_10186_, _10185_, _10107_);
  nand _42548_ (_10187_, _08102_, _07399_);
  nand _42549_ (_28173_[5], _10187_, _10186_);
  nand _42550_ (_10188_, _07364_, word_in[22]);
  nand _42551_ (_10189_, _07377_, word_in[6]);
  nand _42552_ (_10190_, _07378_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nand _42553_ (_10191_, _10190_, _10189_);
  nand _42554_ (_10192_, _10191_, _07371_);
  nand _42555_ (_10193_, _07370_, word_in[14]);
  nand _42556_ (_10195_, _10193_, _10192_);
  nand _42557_ (_10196_, _10195_, _07365_);
  nand _42558_ (_10197_, _10196_, _10188_);
  nand _42559_ (_10198_, _10197_, _10107_);
  nand _42560_ (_10200_, _08283_, _07399_);
  nand _42561_ (_28173_[6], _10200_, _10198_);
  nand _42562_ (_10201_, _04624_, _25099_);
  nand _42563_ (_10202_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  nand _42564_ (_03159_, _10202_, _10201_);
  nand _42565_ (_10204_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  nand _42566_ (_10205_, _08492_, _24927_);
  nand _42567_ (_03161_, _10205_, _10204_);
  nand _42568_ (_10206_, _04624_, _24830_);
  nand _42569_ (_10207_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nand _42570_ (_03167_, _10207_, _10206_);
  nand _42571_ (_10209_, _01182_, _25203_);
  nand _42572_ (_10211_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nand _42573_ (_03196_, _10211_, _10209_);
  nand _42574_ (_10212_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nand _42575_ (_10213_, _08492_, _28096_);
  nand _42576_ (_03202_, _10213_, _10212_);
  nor _42577_ (_10214_, _08142_, _28073_);
  not _42578_ (_10215_, _10214_);
  nand _42579_ (_10216_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  nand _42580_ (_10217_, _10214_, _24927_);
  nand _42581_ (_03212_, _10217_, _10216_);
  nand _42582_ (_10218_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  nand _42583_ (_10220_, _06807_, _24789_);
  nand _42584_ (_03219_, _10220_, _10218_);
  nor _42585_ (_10222_, _24984_, _24795_);
  nand _42586_ (_10223_, _10222_, _25039_);
  not _42587_ (_10224_, _10222_);
  nand _42588_ (_10225_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  nand _42589_ (_03241_, _10225_, _10223_);
  nor _42590_ (_10226_, _28073_, _25159_);
  nand _42591_ (_10228_, _10226_, _25150_);
  not _42592_ (_10230_, _10226_);
  nand _42593_ (_10232_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nand _42594_ (_03245_, _10232_, _10228_);
  nand _42595_ (_10233_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nand _42596_ (_10234_, _06807_, _25150_);
  nand _42597_ (_03247_, _10234_, _10233_);
  nand _42598_ (_10235_, _07009_, word_in[0]);
  nor _42599_ (_10237_, _06846_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _42600_ (_10238_, _06845_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor _42601_ (_10240_, _10238_, _10237_);
  nand _42602_ (_10241_, _10240_, _06849_);
  nor _42603_ (_10242_, _06846_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _42604_ (_10243_, _06845_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _42605_ (_10244_, _10243_, _10242_);
  nand _42606_ (_10245_, _10244_, _06850_);
  nand _42607_ (_10246_, _10245_, _10241_);
  nand _42608_ (_10247_, _10246_, _06863_);
  nor _42609_ (_10248_, _06846_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _42610_ (_10249_, _06845_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _42611_ (_10250_, _10249_, _10248_);
  nand _42612_ (_10251_, _10250_, _06969_);
  nand _42613_ (_10252_, _10251_, _10247_);
  nand _42614_ (_10253_, _10252_, _06858_);
  nor _42615_ (_10254_, _06960_, _06864_);
  not _42616_ (_10255_, _10254_);
  nor _42617_ (_10256_, _06846_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _42618_ (_10257_, _06845_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _42619_ (_10258_, _10257_, _10256_);
  not _42620_ (_10259_, _10258_);
  nor _42621_ (_10260_, _10259_, _10255_);
  nor _42622_ (_10262_, _06846_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _42623_ (_10263_, _06845_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _42624_ (_10264_, _10263_, _10262_);
  not _42625_ (_10265_, _10264_);
  nor _42626_ (_10266_, _10265_, _06850_);
  nor _42627_ (_10267_, _06846_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _42628_ (_10268_, _06845_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _42629_ (_10270_, _10268_, _10267_);
  not _42630_ (_10272_, _10270_);
  nor _42631_ (_10273_, _10272_, _06849_);
  nor _42632_ (_10274_, _10273_, _10266_);
  nor _42633_ (_10275_, _10274_, _06855_);
  nor _42634_ (_10276_, _06846_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _42635_ (_10277_, _06845_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _42636_ (_10278_, _10277_, _10276_);
  nand _42637_ (_10280_, _10278_, _06959_);
  nor _42638_ (_10281_, _06846_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _42639_ (_10282_, _06845_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _42640_ (_10283_, _10282_, _10281_);
  nand _42641_ (_10284_, _10283_, _06969_);
  nand _42642_ (_10285_, _10284_, _10280_);
  nor _42643_ (_10286_, _10285_, _10275_);
  nor _42644_ (_10287_, _10286_, _06858_);
  nor _42645_ (_10288_, _10287_, _10260_);
  nand _42646_ (_10289_, _10288_, _10253_);
  nand _42647_ (_10290_, _10289_, _06944_);
  nand _42648_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _10290_, _10235_);
  nand _42649_ (_10291_, _07009_, word_in[1]);
  nor _42650_ (_10292_, _06846_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _42651_ (_10293_, _06845_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _42652_ (_10294_, _10293_, _10292_);
  nor _42653_ (_10296_, _10294_, _06849_);
  nor _42654_ (_10297_, _06846_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _42655_ (_10298_, _06845_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _42656_ (_10299_, _10298_, _10297_);
  nor _42657_ (_10300_, _10299_, _06850_);
  nor _42658_ (_10302_, _10300_, _10296_);
  nand _42659_ (_10303_, _10302_, _06863_);
  nor _42660_ (_10305_, _06846_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _42661_ (_10306_, _06845_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _42662_ (_10308_, _10306_, _10305_);
  nand _42663_ (_10309_, _10308_, _06969_);
  nand _42664_ (_10311_, _10309_, _10303_);
  nand _42665_ (_10312_, _10311_, _06858_);
  not _42666_ (_10313_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nand _42667_ (_10314_, _06845_, _10313_);
  not _42668_ (_10315_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nand _42669_ (_10316_, _06846_, _10315_);
  nand _42670_ (_10317_, _10316_, _10314_);
  nor _42671_ (_10318_, _10317_, _10255_);
  nand _42672_ (_10319_, _06845_, _08198_);
  nand _42673_ (_10320_, _06846_, _08040_);
  nand _42674_ (_10322_, _10320_, _10319_);
  nand _42675_ (_10324_, _10322_, _06850_);
  nand _42676_ (_10325_, _06845_, _08533_);
  nand _42677_ (_10326_, _06846_, _08393_);
  nand _42678_ (_10327_, _10326_, _10325_);
  nand _42679_ (_10328_, _10327_, _06849_);
  nand _42680_ (_10329_, _10328_, _10324_);
  nor _42681_ (_10330_, _10329_, _06855_);
  nor _42682_ (_10331_, _06846_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _42683_ (_10332_, _06845_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _42684_ (_10333_, _10332_, _10331_);
  nand _42685_ (_10334_, _10333_, _06969_);
  nor _42686_ (_10335_, _06846_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _42687_ (_10336_, _06845_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _42688_ (_10337_, _10336_, _10335_);
  nand _42689_ (_10338_, _10337_, _06959_);
  nand _42690_ (_10339_, _10338_, _10334_);
  nor _42691_ (_10341_, _10339_, _10330_);
  nor _42692_ (_10343_, _10341_, _06858_);
  nor _42693_ (_10345_, _10343_, _10318_);
  nand _42694_ (_10346_, _10345_, _10312_);
  nand _42695_ (_10348_, _10346_, _06944_);
  nand _42696_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _10348_, _10291_);
  nand _42697_ (_10350_, _07009_, word_in[2]);
  nor _42698_ (_10351_, _06846_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _42699_ (_10352_, _06845_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _42700_ (_10353_, _10352_, _10351_);
  nor _42701_ (_10354_, _10353_, _06849_);
  nor _42702_ (_10355_, _06846_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _42703_ (_10356_, _06845_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _42704_ (_10357_, _10356_, _10355_);
  nor _42705_ (_10359_, _10357_, _06850_);
  nor _42706_ (_10360_, _10359_, _10354_);
  nand _42707_ (_10362_, _10360_, _06863_);
  nor _42708_ (_10363_, _06846_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _42709_ (_10365_, _06845_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _42710_ (_10366_, _10365_, _10363_);
  nand _42711_ (_10368_, _10366_, _06969_);
  nand _42712_ (_10369_, _10368_, _10362_);
  nand _42713_ (_10370_, _10369_, _06858_);
  not _42714_ (_10372_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nand _42715_ (_10374_, _06845_, _10372_);
  not _42716_ (_10375_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand _42717_ (_10376_, _06846_, _10375_);
  nand _42718_ (_10377_, _10376_, _10374_);
  nor _42719_ (_10378_, _10377_, _10255_);
  nand _42720_ (_10380_, _06845_, _08216_);
  nand _42721_ (_10381_, _06846_, _08056_);
  nand _42722_ (_10382_, _10381_, _10380_);
  nand _42723_ (_10383_, _10382_, _06850_);
  not _42724_ (_10384_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _42725_ (_10386_, _06845_, _10384_);
  nand _42726_ (_10387_, _06846_, _08407_);
  nand _42727_ (_10388_, _10387_, _10386_);
  nand _42728_ (_10389_, _10388_, _06849_);
  nand _42729_ (_10390_, _10389_, _10383_);
  nor _42730_ (_10391_, _10390_, _06855_);
  nor _42731_ (_10392_, _06846_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _42732_ (_10394_, _06845_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _42733_ (_10395_, _10394_, _10392_);
  nand _42734_ (_10396_, _10395_, _06969_);
  nor _42735_ (_10397_, _06846_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _42736_ (_10398_, _06845_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _42737_ (_10400_, _10398_, _10397_);
  nand _42738_ (_10402_, _10400_, _06959_);
  nand _42739_ (_10404_, _10402_, _10396_);
  nor _42740_ (_10406_, _10404_, _10391_);
  nor _42741_ (_10408_, _10406_, _06858_);
  nor _42742_ (_10409_, _10408_, _10378_);
  nand _42743_ (_10410_, _10409_, _10370_);
  nand _42744_ (_10411_, _10410_, _06944_);
  nand _42745_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _10411_, _10350_);
  nand _42746_ (_10412_, _07009_, word_in[3]);
  nor _42747_ (_10414_, _06846_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _42748_ (_10415_, _06845_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _42749_ (_10416_, _10415_, _10414_);
  nor _42750_ (_10417_, _10416_, _06849_);
  nor _42751_ (_10418_, _06846_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _42752_ (_10420_, _06845_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _42753_ (_10421_, _10420_, _10418_);
  nor _42754_ (_10422_, _10421_, _06850_);
  nor _42755_ (_10423_, _10422_, _10417_);
  nand _42756_ (_10424_, _10423_, _06863_);
  nor _42757_ (_10425_, _06846_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _42758_ (_10426_, _06845_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _42759_ (_10427_, _10426_, _10425_);
  nand _42760_ (_10428_, _10427_, _06969_);
  nand _42761_ (_10429_, _10428_, _10424_);
  nand _42762_ (_10430_, _10429_, _06858_);
  not _42763_ (_10431_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nand _42764_ (_10432_, _06845_, _10431_);
  not _42765_ (_10433_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nand _42766_ (_10434_, _06846_, _10433_);
  nand _42767_ (_10435_, _10434_, _10432_);
  nor _42768_ (_10436_, _10435_, _10255_);
  nand _42769_ (_10437_, _06845_, _08237_);
  not _42770_ (_10438_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nand _42771_ (_10439_, _06846_, _10438_);
  nand _42772_ (_10440_, _10439_, _10437_);
  nand _42773_ (_10441_, _10440_, _06850_);
  not _42774_ (_10442_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nand _42775_ (_10443_, _06845_, _10442_);
  nand _42776_ (_10444_, _06846_, _08419_);
  nand _42777_ (_10445_, _10444_, _10443_);
  nand _42778_ (_10446_, _10445_, _06849_);
  nand _42779_ (_10447_, _10446_, _10441_);
  nor _42780_ (_10449_, _10447_, _06855_);
  nor _42781_ (_10450_, _06846_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _42782_ (_10451_, _06845_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _42783_ (_10452_, _10451_, _10450_);
  nand _42784_ (_10453_, _10452_, _06969_);
  nor _42785_ (_10454_, _06846_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _42786_ (_10455_, _06845_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _42787_ (_10456_, _10455_, _10454_);
  nand _42788_ (_10457_, _10456_, _06959_);
  nand _42789_ (_10458_, _10457_, _10453_);
  nor _42790_ (_10459_, _10458_, _10449_);
  nor _42791_ (_10460_, _10459_, _06858_);
  nor _42792_ (_10461_, _10460_, _10436_);
  nand _42793_ (_10462_, _10461_, _10430_);
  nand _42794_ (_10464_, _10462_, _06944_);
  nand _42795_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _10464_, _10412_);
  nand _42796_ (_10465_, _07009_, word_in[4]);
  nor _42797_ (_10466_, _06846_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _42798_ (_10467_, _06845_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _42799_ (_10468_, _10467_, _10466_);
  nor _42800_ (_10469_, _10468_, _06850_);
  nor _42801_ (_10470_, _06846_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _42802_ (_10471_, _06845_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _42803_ (_10472_, _10471_, _10470_);
  nor _42804_ (_10473_, _10472_, _06849_);
  nor _42805_ (_10474_, _10473_, _10469_);
  nand _42806_ (_10475_, _10474_, _06863_);
  nand _42807_ (_10476_, _06845_, _08878_);
  not _42808_ (_10477_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nand _42809_ (_10478_, _06846_, _10477_);
  nand _42810_ (_10479_, _10478_, _10476_);
  nor _42811_ (_10480_, _10479_, _06970_);
  not _42812_ (_10481_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand _42813_ (_10482_, _06845_, _10481_);
  nand _42814_ (_10483_, _06846_, _09008_);
  nand _42815_ (_10485_, _10483_, _10482_);
  nor _42816_ (_10486_, _10485_, _06960_);
  nor _42817_ (_10487_, _10486_, _10480_);
  nand _42818_ (_10489_, _10487_, _10475_);
  nand _42819_ (_10490_, _10489_, _06864_);
  not _42820_ (_10491_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nand _42821_ (_10492_, _06845_, _10491_);
  not _42822_ (_10493_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nand _42823_ (_10494_, _06846_, _10493_);
  nand _42824_ (_10495_, _10494_, _10492_);
  nor _42825_ (_10497_, _10495_, _06850_);
  not _42826_ (_10498_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nand _42827_ (_10499_, _06845_, _10498_);
  not _42828_ (_10500_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nand _42829_ (_10501_, _06846_, _10500_);
  nand _42830_ (_10503_, _10501_, _10499_);
  nor _42831_ (_10504_, _10503_, _06849_);
  nor _42832_ (_10505_, _10504_, _10497_);
  nor _42833_ (_10506_, _10505_, _06855_);
  not _42834_ (_10507_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nand _42835_ (_10508_, _06845_, _10507_);
  not _42836_ (_10509_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand _42837_ (_10510_, _06846_, _10509_);
  nand _42838_ (_10511_, _10510_, _10508_);
  nor _42839_ (_10512_, _10511_, _06970_);
  nor _42840_ (_10514_, _10512_, _10506_);
  nor _42841_ (_10515_, _10514_, _06864_);
  not _42842_ (_10516_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand _42843_ (_10517_, _06845_, _10516_);
  not _42844_ (_10518_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nand _42845_ (_10519_, _06846_, _10518_);
  nand _42846_ (_10520_, _10519_, _10517_);
  nor _42847_ (_10522_, _10520_, _10255_);
  nor _42848_ (_10524_, _10522_, _10515_);
  nand _42849_ (_10526_, _10524_, _10490_);
  nand _42850_ (_10527_, _10526_, _06944_);
  nand _42851_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _10527_, _10465_);
  nand _42852_ (_10528_, _07009_, word_in[5]);
  nor _42853_ (_10529_, _06846_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _42854_ (_10530_, _06845_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _42855_ (_10531_, _10530_, _10529_);
  nor _42856_ (_10532_, _10531_, _06849_);
  nor _42857_ (_10533_, _06846_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _42858_ (_10534_, _06845_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _42859_ (_10535_, _10534_, _10533_);
  nor _42860_ (_10537_, _10535_, _06850_);
  nor _42861_ (_10538_, _10537_, _10532_);
  nand _42862_ (_10539_, _10538_, _06863_);
  nor _42863_ (_10540_, _06846_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _42864_ (_10541_, _06845_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _42865_ (_10542_, _10541_, _10540_);
  nand _42866_ (_10543_, _10542_, _06969_);
  nand _42867_ (_10544_, _10543_, _10539_);
  nand _42868_ (_10545_, _10544_, _06858_);
  not _42869_ (_10546_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nand _42870_ (_10547_, _06845_, _10546_);
  not _42871_ (_10548_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nand _42872_ (_10549_, _06846_, _10548_);
  nand _42873_ (_10550_, _10549_, _10547_);
  nor _42874_ (_10551_, _10550_, _10255_);
  nand _42875_ (_10552_, _06845_, _08269_);
  nand _42876_ (_10553_, _06846_, _08104_);
  nand _42877_ (_10554_, _10553_, _10552_);
  nand _42878_ (_10555_, _10554_, _06850_);
  nand _42879_ (_10557_, _06845_, _08604_);
  nand _42880_ (_10559_, _06846_, _08447_);
  nand _42881_ (_10560_, _10559_, _10557_);
  nand _42882_ (_10561_, _10560_, _06849_);
  nand _42883_ (_10563_, _10561_, _10555_);
  nor _42884_ (_10564_, _10563_, _06855_);
  nor _42885_ (_10565_, _06846_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _42886_ (_10566_, _06845_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _42887_ (_10567_, _10566_, _10565_);
  nand _42888_ (_10568_, _10567_, _06969_);
  nor _42889_ (_10569_, _06846_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _42890_ (_10570_, _06845_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _42891_ (_10571_, _10570_, _10569_);
  nand _42892_ (_10572_, _10571_, _06959_);
  nand _42893_ (_10573_, _10572_, _10568_);
  nor _42894_ (_10574_, _10573_, _10564_);
  nor _42895_ (_10575_, _10574_, _06858_);
  nor _42896_ (_10576_, _10575_, _10551_);
  nand _42897_ (_10577_, _10576_, _10545_);
  nand _42898_ (_10578_, _10577_, _06944_);
  nand _42899_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _10578_, _10528_);
  nand _42900_ (_10579_, _07009_, word_in[6]);
  nor _42901_ (_10580_, _06846_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _42902_ (_10581_, _06845_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _42903_ (_10582_, _10581_, _10580_);
  nand _42904_ (_10583_, _10582_, _06849_);
  nor _42905_ (_10584_, _06846_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _42906_ (_10585_, _06845_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _42907_ (_10586_, _10585_, _10584_);
  nand _42908_ (_10588_, _10586_, _06850_);
  nand _42909_ (_10589_, _10588_, _10583_);
  nand _42910_ (_10590_, _10589_, _06863_);
  nor _42911_ (_10591_, _06846_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _42912_ (_10592_, _06845_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _42913_ (_10593_, _10592_, _10591_);
  nand _42914_ (_10594_, _10593_, _06969_);
  nand _42915_ (_10595_, _10594_, _10590_);
  nand _42916_ (_10596_, _10595_, _06858_);
  nor _42917_ (_10597_, _06846_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _42918_ (_10598_, _06845_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _42919_ (_10599_, _10598_, _10597_);
  not _42920_ (_10600_, _10599_);
  nor _42921_ (_10602_, _10600_, _10255_);
  nor _42922_ (_10603_, _06846_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _42923_ (_10604_, _06845_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _42924_ (_10605_, _10604_, _10603_);
  not _42925_ (_10606_, _10605_);
  nor _42926_ (_10607_, _10606_, _06850_);
  nor _42927_ (_10608_, _06846_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _42928_ (_10609_, _06845_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _42929_ (_10611_, _10609_, _10608_);
  not _42930_ (_10613_, _10611_);
  nor _42931_ (_10615_, _10613_, _06849_);
  nor _42932_ (_10616_, _10615_, _10607_);
  nor _42933_ (_10617_, _10616_, _06855_);
  nor _42934_ (_10619_, _06846_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _42935_ (_10620_, _06845_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _42936_ (_10621_, _10620_, _10619_);
  nand _42937_ (_10622_, _10621_, _06959_);
  nor _42938_ (_10623_, _06846_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _42939_ (_10624_, _06845_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _42940_ (_10625_, _10624_, _10623_);
  nand _42941_ (_10626_, _10625_, _06969_);
  nand _42942_ (_10627_, _10626_, _10622_);
  nor _42943_ (_10628_, _10627_, _10617_);
  nor _42944_ (_10629_, _10628_, _06858_);
  nor _42945_ (_10630_, _10629_, _10602_);
  nand _42946_ (_10631_, _10630_, _10596_);
  nand _42947_ (_10632_, _10631_, _06944_);
  nand _42948_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _10632_, _10579_);
  nand _42949_ (_10633_, _07157_, word_in[8]);
  nor _42950_ (_10635_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor _42951_ (_10636_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _42952_ (_10638_, _10636_, _10635_);
  nand _42953_ (_10639_, _10638_, _07100_);
  nor _42954_ (_10641_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _42955_ (_10642_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _42956_ (_10643_, _10642_, _10641_);
  nand _42957_ (_10644_, _10643_, _07093_);
  nand _42958_ (_10645_, _10644_, _10639_);
  nor _42959_ (_10646_, _10645_, _07022_);
  nor _42960_ (_10648_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _42961_ (_10649_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _42962_ (_10650_, _10649_, _10648_);
  nand _42963_ (_10651_, _10650_, _07100_);
  nor _42964_ (_10652_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _42965_ (_10653_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _42966_ (_10654_, _10653_, _10652_);
  nand _42967_ (_10655_, _10654_, _07093_);
  nand _42968_ (_10657_, _10655_, _10651_);
  nor _42969_ (_10658_, _10657_, _07030_);
  nor _42970_ (_10659_, _10658_, _10646_);
  nand _42971_ (_10661_, _10659_, _07019_);
  nor _42972_ (_10662_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _42973_ (_10663_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _42974_ (_10664_, _10663_, _10662_);
  nand _42975_ (_10665_, _10664_, _07100_);
  nor _42976_ (_10666_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _42977_ (_10667_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _42978_ (_10668_, _10667_, _10666_);
  nand _42979_ (_10669_, _10668_, _07093_);
  nand _42980_ (_10671_, _10669_, _10665_);
  nand _42981_ (_10672_, _10671_, _07030_);
  nor _42982_ (_10673_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _42983_ (_10674_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _42984_ (_10675_, _10674_, _10673_);
  nand _42985_ (_10677_, _10675_, _07100_);
  nor _42986_ (_10679_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _42987_ (_10680_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _42988_ (_10681_, _10680_, _10679_);
  nand _42989_ (_10682_, _10681_, _07093_);
  nand _42990_ (_10683_, _10682_, _10677_);
  nand _42991_ (_10684_, _10683_, _07022_);
  nand _42992_ (_10686_, _10684_, _10672_);
  nand _42993_ (_10687_, _10686_, _07017_);
  nand _42994_ (_10688_, _10687_, _10661_);
  nand _42995_ (_10689_, _10688_, _07091_);
  nand _42996_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _10689_, _10633_);
  nand _42997_ (_10690_, _07157_, word_in[9]);
  nor _42998_ (_10692_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _42999_ (_10693_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _43000_ (_10694_, _10693_, _10692_);
  nand _43001_ (_10696_, _10694_, _07100_);
  nor _43002_ (_10697_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _43003_ (_10698_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _43004_ (_10699_, _10698_, _10697_);
  nand _43005_ (_10700_, _10699_, _07093_);
  nand _43006_ (_10702_, _10700_, _10696_);
  nor _43007_ (_10703_, _10702_, _07030_);
  nor _43008_ (_10704_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _43009_ (_10706_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _43010_ (_10707_, _10706_, _10704_);
  nand _43011_ (_10708_, _10707_, _07100_);
  nor _43012_ (_10710_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _43013_ (_10711_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _43014_ (_10712_, _10711_, _10710_);
  nand _43015_ (_10714_, _10712_, _07093_);
  nand _43016_ (_10715_, _10714_, _10708_);
  nor _43017_ (_10716_, _10715_, _07022_);
  nor _43018_ (_10717_, _10716_, _10703_);
  nand _43019_ (_10718_, _10717_, _07019_);
  nor _43020_ (_10720_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _43021_ (_10721_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _43022_ (_10722_, _10721_, _10720_);
  nand _43023_ (_10723_, _10722_, _07100_);
  nor _43024_ (_10725_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _43025_ (_10726_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _43026_ (_10728_, _10726_, _10725_);
  nand _43027_ (_10729_, _10728_, _07093_);
  nand _43028_ (_10731_, _10729_, _10723_);
  nand _43029_ (_10733_, _10731_, _07030_);
  nor _43030_ (_10734_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _43031_ (_10735_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _43032_ (_10736_, _10735_, _10734_);
  nand _43033_ (_10737_, _10736_, _07100_);
  nor _43034_ (_10738_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _43035_ (_10740_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _43036_ (_10741_, _10740_, _10738_);
  nand _43037_ (_10742_, _10741_, _07093_);
  nand _43038_ (_10743_, _10742_, _10737_);
  nand _43039_ (_10745_, _10743_, _07022_);
  nand _43040_ (_10746_, _10745_, _10733_);
  nand _43041_ (_10747_, _10746_, _07017_);
  nand _43042_ (_10748_, _10747_, _10718_);
  nand _43043_ (_10749_, _10748_, _07091_);
  nand _43044_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _10749_, _10690_);
  nand _43045_ (_10750_, _07157_, word_in[10]);
  nor _43046_ (_10751_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _43047_ (_10752_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _43048_ (_10753_, _10752_, _10751_);
  nand _43049_ (_10754_, _10753_, _07100_);
  nor _43050_ (_10755_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _43051_ (_10756_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _43052_ (_10758_, _10756_, _10755_);
  nand _43053_ (_10759_, _10758_, _07093_);
  nand _43054_ (_10760_, _10759_, _10754_);
  nor _43055_ (_10761_, _10760_, _07022_);
  nor _43056_ (_10762_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _43057_ (_10763_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _43058_ (_10764_, _10763_, _10762_);
  nand _43059_ (_10765_, _10764_, _07100_);
  nor _43060_ (_10767_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _43061_ (_10768_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _43062_ (_10769_, _10768_, _10767_);
  nand _43063_ (_10770_, _10769_, _07093_);
  nand _43064_ (_10771_, _10770_, _10765_);
  nor _43065_ (_10772_, _10771_, _07030_);
  nor _43066_ (_10774_, _10772_, _10761_);
  nand _43067_ (_10775_, _10774_, _07019_);
  nor _43068_ (_10776_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _43069_ (_10777_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _43070_ (_10778_, _10777_, _10776_);
  nand _43071_ (_10780_, _10778_, _07100_);
  nor _43072_ (_10781_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _43073_ (_10782_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _43074_ (_10783_, _10782_, _10781_);
  nand _43075_ (_10784_, _10783_, _07093_);
  nand _43076_ (_10785_, _10784_, _10780_);
  nand _43077_ (_10786_, _10785_, _07030_);
  nor _43078_ (_10787_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _43079_ (_10788_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _43080_ (_10789_, _10788_, _10787_);
  nand _43081_ (_10790_, _10789_, _07100_);
  nor _43082_ (_10791_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _43083_ (_10793_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _43084_ (_10794_, _10793_, _10791_);
  nand _43085_ (_10795_, _10794_, _07093_);
  nand _43086_ (_10796_, _10795_, _10790_);
  nand _43087_ (_10797_, _10796_, _07022_);
  nand _43088_ (_10798_, _10797_, _10786_);
  nand _43089_ (_10800_, _10798_, _07017_);
  nand _43090_ (_10801_, _10800_, _10775_);
  nand _43091_ (_10803_, _10801_, _07091_);
  nand _43092_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _10803_, _10750_);
  nand _43093_ (_10804_, _07157_, word_in[11]);
  nor _43094_ (_10805_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _43095_ (_10806_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _43096_ (_10808_, _10806_, _10805_);
  nand _43097_ (_10809_, _10808_, _07100_);
  nor _43098_ (_10811_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _43099_ (_10812_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _43100_ (_10813_, _10812_, _10811_);
  nand _43101_ (_10814_, _10813_, _07093_);
  nand _43102_ (_10815_, _10814_, _10809_);
  nor _43103_ (_10816_, _10815_, _07030_);
  nor _43104_ (_10817_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _43105_ (_10818_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _43106_ (_10819_, _10818_, _10817_);
  nand _43107_ (_10820_, _10819_, _07100_);
  nor _43108_ (_10821_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _43109_ (_10822_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _43110_ (_10824_, _10822_, _10821_);
  nand _43111_ (_10826_, _10824_, _07093_);
  nand _43112_ (_10827_, _10826_, _10820_);
  nor _43113_ (_10828_, _10827_, _07022_);
  nor _43114_ (_10830_, _10828_, _10816_);
  nand _43115_ (_10831_, _10830_, _07019_);
  nor _43116_ (_10833_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _43117_ (_10834_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _43118_ (_10835_, _10834_, _10833_);
  nand _43119_ (_10836_, _10835_, _07100_);
  nor _43120_ (_10837_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _43121_ (_10838_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _43122_ (_10839_, _10838_, _10837_);
  nand _43123_ (_10840_, _10839_, _07093_);
  nand _43124_ (_10841_, _10840_, _10836_);
  nand _43125_ (_10843_, _10841_, _07030_);
  nor _43126_ (_10844_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _43127_ (_10846_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _43128_ (_10847_, _10846_, _10844_);
  nand _43129_ (_10848_, _10847_, _07100_);
  nor _43130_ (_10849_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _43131_ (_10850_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _43132_ (_10851_, _10850_, _10849_);
  nand _43133_ (_10852_, _10851_, _07093_);
  nand _43134_ (_10853_, _10852_, _10848_);
  nand _43135_ (_10855_, _10853_, _07022_);
  nand _43136_ (_10856_, _10855_, _10843_);
  nand _43137_ (_10857_, _10856_, _07017_);
  nand _43138_ (_10858_, _10857_, _10831_);
  nand _43139_ (_10859_, _10858_, _07091_);
  nand _43140_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _10859_, _10804_);
  nand _43141_ (_10860_, _07157_, word_in[12]);
  nor _43142_ (_10862_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _43143_ (_10863_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _43144_ (_10864_, _10863_, _10862_);
  nand _43145_ (_10865_, _10864_, _07100_);
  nor _43146_ (_10866_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _43147_ (_10867_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _43148_ (_10868_, _10867_, _10866_);
  nand _43149_ (_10870_, _10868_, _07093_);
  nand _43150_ (_10871_, _10870_, _10865_);
  nor _43151_ (_10872_, _10871_, _07030_);
  nor _43152_ (_10873_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _43153_ (_10874_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _43154_ (_10875_, _10874_, _10873_);
  nand _43155_ (_10876_, _10875_, _07100_);
  nor _43156_ (_10877_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _43157_ (_10879_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _43158_ (_10880_, _10879_, _10877_);
  nand _43159_ (_10881_, _10880_, _07093_);
  nand _43160_ (_10882_, _10881_, _10876_);
  nor _43161_ (_10883_, _10882_, _07022_);
  nor _43162_ (_10884_, _10883_, _10872_);
  nand _43163_ (_10886_, _10884_, _07019_);
  nor _43164_ (_10887_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _43165_ (_10888_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _43166_ (_10889_, _10888_, _10887_);
  nand _43167_ (_10890_, _10889_, _07100_);
  nor _43168_ (_10892_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _43169_ (_10893_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _43170_ (_10894_, _10893_, _10892_);
  nand _43171_ (_10895_, _10894_, _07093_);
  nand _43172_ (_10896_, _10895_, _10890_);
  nand _43173_ (_10897_, _10896_, _07030_);
  nor _43174_ (_10899_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _43175_ (_10901_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _43176_ (_10902_, _10901_, _10899_);
  nand _43177_ (_10903_, _10902_, _07100_);
  nor _43178_ (_10905_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _43179_ (_10906_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _43180_ (_10907_, _10906_, _10905_);
  nand _43181_ (_10909_, _10907_, _07093_);
  nand _43182_ (_10910_, _10909_, _10903_);
  nand _43183_ (_10911_, _10910_, _07022_);
  nand _43184_ (_10912_, _10911_, _10897_);
  nand _43185_ (_10913_, _10912_, _07017_);
  nand _43186_ (_10915_, _10913_, _10886_);
  nand _43187_ (_10916_, _10915_, _07091_);
  nand _43188_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _10916_, _10860_);
  nand _43189_ (_10918_, _07157_, word_in[13]);
  nor _43190_ (_10920_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _43191_ (_10922_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _43192_ (_10923_, _10922_, _10920_);
  nand _43193_ (_10925_, _10923_, _07100_);
  nor _43194_ (_10926_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _43195_ (_10927_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _43196_ (_10928_, _10927_, _10926_);
  nand _43197_ (_10929_, _10928_, _07093_);
  nand _43198_ (_10931_, _10929_, _10925_);
  nor _43199_ (_10932_, _10931_, _07030_);
  nor _43200_ (_10933_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _43201_ (_10934_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _43202_ (_10935_, _10934_, _10933_);
  nand _43203_ (_10936_, _10935_, _07100_);
  nor _43204_ (_10937_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _43205_ (_10939_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _43206_ (_10940_, _10939_, _10937_);
  nand _43207_ (_10942_, _10940_, _07093_);
  nand _43208_ (_10944_, _10942_, _10936_);
  nor _43209_ (_10946_, _10944_, _07022_);
  nor _43210_ (_10948_, _10946_, _10932_);
  nand _43211_ (_10950_, _10948_, _07019_);
  nor _43212_ (_10951_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _43213_ (_10952_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _43214_ (_10953_, _10952_, _10951_);
  nand _43215_ (_10955_, _10953_, _07100_);
  nor _43216_ (_10956_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _43217_ (_10957_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _43218_ (_10958_, _10957_, _10956_);
  nand _43219_ (_10959_, _10958_, _07093_);
  nand _43220_ (_10961_, _10959_, _10955_);
  nand _43221_ (_10962_, _10961_, _07030_);
  nor _43222_ (_10964_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _43223_ (_10965_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _43224_ (_10966_, _10965_, _10964_);
  nand _43225_ (_10967_, _10966_, _07100_);
  nor _43226_ (_10969_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _43227_ (_10970_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _43228_ (_10971_, _10970_, _10969_);
  nand _43229_ (_10973_, _10971_, _07093_);
  nand _43230_ (_10974_, _10973_, _10967_);
  nand _43231_ (_10975_, _10974_, _07022_);
  nand _43232_ (_10977_, _10975_, _10962_);
  nand _43233_ (_10978_, _10977_, _07017_);
  nand _43234_ (_10979_, _10978_, _10950_);
  nand _43235_ (_10980_, _10979_, _07091_);
  nand _43236_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _10980_, _10918_);
  nand _43237_ (_10983_, _07157_, word_in[14]);
  nor _43238_ (_10984_, _06846_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _43239_ (_10986_, _06845_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _43240_ (_10988_, _10986_, _10984_);
  nand _43241_ (_10989_, _10988_, _07100_);
  nor _43242_ (_10990_, _06846_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _43243_ (_10991_, _06845_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _43244_ (_10992_, _10991_, _10990_);
  nand _43245_ (_10994_, _10992_, _07093_);
  nand _43246_ (_10995_, _10994_, _10989_);
  nor _43247_ (_10996_, _10995_, _07022_);
  nor _43248_ (_10998_, _06846_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _43249_ (_11000_, _06845_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _43250_ (_11002_, _11000_, _10998_);
  nand _43251_ (_11003_, _11002_, _07100_);
  nor _43252_ (_11004_, _06846_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _43253_ (_11006_, _06845_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _43254_ (_11007_, _11006_, _11004_);
  nand _43255_ (_11008_, _11007_, _07093_);
  nand _43256_ (_11009_, _11008_, _11003_);
  nor _43257_ (_11010_, _11009_, _07030_);
  nor _43258_ (_11011_, _11010_, _10996_);
  nand _43259_ (_11012_, _11011_, _07019_);
  nor _43260_ (_11014_, _06846_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _43261_ (_11015_, _06845_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _43262_ (_11016_, _11015_, _11014_);
  nand _43263_ (_11017_, _11016_, _07100_);
  nor _43264_ (_11018_, _06846_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _43265_ (_11020_, _06845_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _43266_ (_11021_, _11020_, _11018_);
  nand _43267_ (_11023_, _11021_, _07093_);
  nand _43268_ (_11025_, _11023_, _11017_);
  nand _43269_ (_11027_, _11025_, _07030_);
  nor _43270_ (_11029_, _06846_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _43271_ (_11031_, _06845_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _43272_ (_11033_, _11031_, _11029_);
  nand _43273_ (_11035_, _11033_, _07100_);
  nor _43274_ (_11037_, _06846_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _43275_ (_11038_, _06845_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _43276_ (_11040_, _11038_, _11037_);
  nand _43277_ (_11042_, _11040_, _07093_);
  nand _43278_ (_11044_, _11042_, _11035_);
  nand _43279_ (_11046_, _11044_, _07022_);
  nand _43280_ (_11048_, _11046_, _11027_);
  nand _43281_ (_11049_, _11048_, _07017_);
  nand _43282_ (_11050_, _11049_, _11012_);
  nand _43283_ (_11051_, _11050_, _07091_);
  nand _43284_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _11051_, _10983_);
  nor _43285_ (_11054_, _10240_, _06849_);
  nor _43286_ (_11055_, _10244_, _06850_);
  nor _43287_ (_11057_, _11055_, _11054_);
  nand _43288_ (_11058_, _11057_, _07166_);
  nor _43289_ (_11059_, _10259_, _06970_);
  not _43290_ (_11061_, _10250_);
  nor _43291_ (_11062_, _11061_, _07236_);
  nor _43292_ (_11063_, _11062_, _11059_);
  nand _43293_ (_11064_, _11063_, _11058_);
  nand _43294_ (_11065_, _11064_, _07178_);
  nor _43295_ (_11067_, _10264_, _06849_);
  nor _43296_ (_11069_, _10270_, _06850_);
  nor _43297_ (_11071_, _11069_, _11067_);
  nand _43298_ (_11073_, _11071_, _07166_);
  nand _43299_ (_11075_, _10283_, _06849_);
  nand _43300_ (_11076_, _10278_, _06850_);
  nand _43301_ (_11078_, _11076_, _11075_);
  nand _43302_ (_11079_, _11078_, _07167_);
  nand _43303_ (_11081_, _11079_, _11073_);
  nand _43304_ (_11083_, _11081_, _07163_);
  nand _43305_ (_11085_, _11083_, _11065_);
  nand _43306_ (_11086_, _11085_, _07226_);
  nand _43307_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _11086_, _08693_);
  nor _43308_ (_11087_, _10299_, _06849_);
  nor _43309_ (_11088_, _10294_, _06850_);
  nor _43310_ (_11089_, _11088_, _11087_);
  nand _43311_ (_11091_, _11089_, _07166_);
  nor _43312_ (_11092_, _10317_, _06970_);
  not _43313_ (_11093_, _10308_);
  nor _43314_ (_11094_, _11093_, _07236_);
  nor _43315_ (_11096_, _11094_, _11092_);
  nand _43316_ (_11098_, _11096_, _11091_);
  nand _43317_ (_11100_, _11098_, _07178_);
  nand _43318_ (_11101_, _10333_, _07164_);
  nand _43319_ (_11102_, _10327_, _06850_);
  nand _43320_ (_11104_, _10322_, _06849_);
  nand _43321_ (_11105_, _11104_, _11102_);
  nor _43322_ (_11107_, _11105_, _07167_);
  not _43323_ (_11109_, _10337_);
  nor _43324_ (_11111_, _11109_, _06970_);
  nor _43325_ (_11113_, _11111_, _11107_);
  nand _43326_ (_11114_, _11113_, _11101_);
  nand _43327_ (_11116_, _11114_, _07163_);
  nand _43328_ (_11118_, _11116_, _11100_);
  nand _43329_ (_11119_, _11118_, _07226_);
  nand _43330_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _11119_, _08401_);
  nand _43331_ (_11122_, _10388_, _06850_);
  nand _43332_ (_11124_, _10382_, _06849_);
  nand _43333_ (_11125_, _11124_, _11122_);
  nor _43334_ (_11126_, _11125_, _07167_);
  nand _43335_ (_11127_, _10395_, _06849_);
  nand _43336_ (_11129_, _10400_, _06850_);
  nand _43337_ (_11130_, _11129_, _11127_);
  nand _43338_ (_11131_, _11130_, _07167_);
  nand _43339_ (_11132_, _11131_, _07163_);
  nor _43340_ (_11134_, _11132_, _11126_);
  not _43341_ (_11135_, _10357_);
  nand _43342_ (_11137_, _11135_, _06850_);
  not _43343_ (_11139_, _10353_);
  nand _43344_ (_11141_, _11139_, _06849_);
  nand _43345_ (_11143_, _11141_, _11137_);
  nor _43346_ (_11144_, _11143_, _07167_);
  nor _43347_ (_11145_, _10377_, _06970_);
  not _43348_ (_11147_, _10366_);
  nor _43349_ (_11148_, _11147_, _07236_);
  nor _43350_ (_11150_, _11148_, _11145_);
  nand _43351_ (_11152_, _11150_, _07178_);
  nor _43352_ (_11153_, _11152_, _11144_);
  nor _43353_ (_11155_, _11153_, _11134_);
  nand _43354_ (_11156_, _11155_, _07226_);
  nand _43355_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _11156_, _08717_);
  nand _43356_ (_11158_, _10445_, _06850_);
  nand _43357_ (_11160_, _10440_, _06849_);
  nand _43358_ (_11162_, _11160_, _11158_);
  nor _43359_ (_11163_, _11162_, _07167_);
  nand _43360_ (_11165_, _10452_, _06849_);
  nand _43361_ (_11166_, _10456_, _06850_);
  nand _43362_ (_11167_, _11166_, _11165_);
  nand _43363_ (_11168_, _11167_, _07167_);
  nand _43364_ (_11170_, _11168_, _07163_);
  nor _43365_ (_11172_, _11170_, _11163_);
  not _43366_ (_11174_, _10421_);
  nand _43367_ (_11175_, _11174_, _06850_);
  not _43368_ (_11176_, _10416_);
  nand _43369_ (_11177_, _11176_, _06849_);
  nand _43370_ (_11180_, _11177_, _11175_);
  nor _43371_ (_11182_, _11180_, _07167_);
  nor _43372_ (_11184_, _10435_, _06970_);
  not _43373_ (_11186_, _10427_);
  nor _43374_ (_11188_, _11186_, _07236_);
  nor _43375_ (_11190_, _11188_, _11184_);
  nand _43376_ (_11191_, _11190_, _07178_);
  nor _43377_ (_11192_, _11191_, _11182_);
  nor _43378_ (_11194_, _11192_, _11172_);
  nand _43379_ (_11195_, _11194_, _07226_);
  nand _43380_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _11195_, _08247_);
  not _43381_ (_11197_, _10468_);
  nand _43382_ (_11198_, _11197_, _06850_);
  not _43383_ (_11199_, _10472_);
  nand _43384_ (_11200_, _11199_, _06849_);
  nand _43385_ (_11201_, _11200_, _11198_);
  nor _43386_ (_11202_, _11201_, _07167_);
  nor _43387_ (_11204_, _10485_, _06970_);
  nor _43388_ (_11205_, _10479_, _07236_);
  nor _43389_ (_11206_, _11205_, _11204_);
  nand _43390_ (_11207_, _11206_, _07163_);
  nor _43391_ (_11209_, _11207_, _11202_);
  nand _43392_ (_11211_, _10495_, _06850_);
  nand _43393_ (_11213_, _10503_, _06849_);
  nand _43394_ (_11215_, _11213_, _11211_);
  nor _43395_ (_11216_, _11215_, _07167_);
  nor _43396_ (_11217_, _10520_, _06970_);
  nor _43397_ (_11219_, _10511_, _07236_);
  nor _43398_ (_11220_, _11219_, _11217_);
  nand _43399_ (_11222_, _11220_, _07178_);
  nor _43400_ (_11224_, _11222_, _11216_);
  nor _43401_ (_11225_, _11224_, _11209_);
  nand _43402_ (_11227_, _11225_, _07226_);
  nand _43403_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _11227_, _08761_);
  nor _43404_ (_11229_, _10535_, _06849_);
  nor _43405_ (_11230_, _10531_, _06850_);
  nor _43406_ (_11232_, _11230_, _11229_);
  nand _43407_ (_11234_, _11232_, _07166_);
  nor _43408_ (_11235_, _10550_, _06970_);
  not _43409_ (_11236_, _10542_);
  nor _43410_ (_11237_, _11236_, _07236_);
  nor _43411_ (_11239_, _11237_, _11235_);
  nand _43412_ (_11241_, _11239_, _11234_);
  nand _43413_ (_11242_, _11241_, _07178_);
  nand _43414_ (_11243_, _10571_, _06969_);
  nand _43415_ (_11245_, _10560_, _06850_);
  nand _43416_ (_11246_, _10554_, _06849_);
  nand _43417_ (_11248_, _11246_, _11245_);
  nor _43418_ (_11250_, _11248_, _07167_);
  not _43419_ (_11251_, _10567_);
  nor _43420_ (_11253_, _11251_, _07236_);
  nor _43421_ (_11254_, _11253_, _11250_);
  nand _43422_ (_11255_, _11254_, _11243_);
  nand _43423_ (_11256_, _11255_, _07163_);
  nand _43424_ (_11258_, _11256_, _11242_);
  nand _43425_ (_11259_, _11258_, _07226_);
  nand _43426_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11259_, _08612_);
  nand _43427_ (_11260_, _10586_, _06849_);
  nand _43428_ (_11261_, _10582_, _06850_);
  nand _43429_ (_11263_, _11261_, _11260_);
  nand _43430_ (_11264_, _11263_, _07166_);
  not _43431_ (_11265_, _10593_);
  nor _43432_ (_11267_, _11265_, _07236_);
  nor _43433_ (_11269_, _10600_, _06970_);
  nor _43434_ (_11271_, _11269_, _11267_);
  nand _43435_ (_11273_, _11271_, _11264_);
  nand _43436_ (_11275_, _11273_, _07178_);
  nor _43437_ (_11276_, _10605_, _06849_);
  nor _43438_ (_11278_, _10611_, _06850_);
  nor _43439_ (_11279_, _11278_, _11276_);
  nand _43440_ (_11281_, _11279_, _07166_);
  nand _43441_ (_11283_, _10625_, _06849_);
  nand _43442_ (_11284_, _10621_, _06850_);
  nand _43443_ (_11286_, _11284_, _11283_);
  nand _43444_ (_11288_, _11286_, _07167_);
  nand _43445_ (_11289_, _11288_, _11281_);
  nand _43446_ (_11290_, _11289_, _07163_);
  nand _43447_ (_11291_, _11290_, _11275_);
  nand _43448_ (_11293_, _11291_, _07226_);
  nand _43449_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11293_, _08297_);
  nand _43450_ (_11296_, _10650_, _07093_);
  nand _43451_ (_11297_, _10654_, _07100_);
  nand _43452_ (_11299_, _11297_, _11296_);
  nand _43453_ (_11301_, _11299_, _07263_);
  nand _43454_ (_11303_, _10638_, _07093_);
  nand _43455_ (_11304_, _10643_, _07100_);
  nand _43456_ (_11306_, _11304_, _11303_);
  nand _43457_ (_11307_, _11306_, _07264_);
  nand _43458_ (_11309_, _11307_, _11301_);
  nand _43459_ (_11311_, _11309_, _07259_);
  nand _43460_ (_11312_, _10675_, _07093_);
  nand _43461_ (_11314_, _10681_, _07100_);
  nand _43462_ (_11316_, _11314_, _11312_);
  nand _43463_ (_11318_, _11316_, _07263_);
  nand _43464_ (_11319_, _10668_, _07100_);
  nand _43465_ (_11320_, _10664_, _07093_);
  nand _43466_ (_11322_, _11320_, _11319_);
  nand _43467_ (_11323_, _11322_, _07264_);
  nand _43468_ (_11325_, _11323_, _11318_);
  nand _43469_ (_11327_, _11325_, _07271_);
  nand _43470_ (_11329_, _11327_, _11311_);
  nand _43471_ (_11331_, _11329_, _07324_);
  nand _43472_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11331_, _08698_);
  nand _43473_ (_11333_, _10694_, _07093_);
  nand _43474_ (_11334_, _10699_, _07100_);
  nand _43475_ (_11336_, _11334_, _11333_);
  nand _43476_ (_11337_, _11336_, _07263_);
  nand _43477_ (_11338_, _10712_, _07100_);
  nand _43478_ (_11339_, _10707_, _07093_);
  nand _43479_ (_11341_, _11339_, _11338_);
  nand _43480_ (_11342_, _11341_, _07264_);
  nand _43481_ (_11344_, _11342_, _11337_);
  nand _43482_ (_11345_, _11344_, _07259_);
  nand _43483_ (_11347_, _10736_, _07093_);
  nand _43484_ (_11349_, _10741_, _07100_);
  nand _43485_ (_11350_, _11349_, _11347_);
  nand _43486_ (_11352_, _11350_, _07263_);
  nand _43487_ (_11354_, _10728_, _07100_);
  nand _43488_ (_11356_, _10722_, _07093_);
  nand _43489_ (_11357_, _11356_, _11354_);
  nand _43490_ (_11358_, _11357_, _07264_);
  nand _43491_ (_11359_, _11358_, _11352_);
  nand _43492_ (_11360_, _11359_, _07271_);
  nand _43493_ (_11361_, _11360_, _11345_);
  nand _43494_ (_11363_, _11361_, _07324_);
  nand _43495_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _11363_, _08037_);
  nand _43496_ (_11366_, _10764_, _07093_);
  nand _43497_ (_11368_, _10769_, _07100_);
  nand _43498_ (_11370_, _11368_, _11366_);
  nand _43499_ (_11372_, _11370_, _07263_);
  nand _43500_ (_11373_, _10758_, _07100_);
  nand _43501_ (_11374_, _10753_, _07093_);
  nand _43502_ (_11375_, _11374_, _11373_);
  nand _43503_ (_11376_, _11375_, _07264_);
  nand _43504_ (_11378_, _11376_, _11372_);
  nand _43505_ (_11379_, _11378_, _07259_);
  nand _43506_ (_11381_, _10789_, _07093_);
  nand _43507_ (_11382_, _10794_, _07100_);
  nand _43508_ (_11383_, _11382_, _11381_);
  nand _43509_ (_11385_, _11383_, _07263_);
  nand _43510_ (_11386_, _10783_, _07100_);
  nand _43511_ (_11387_, _10778_, _07093_);
  nand _43512_ (_11388_, _11387_, _11386_);
  nand _43513_ (_11389_, _11388_, _07264_);
  nand _43514_ (_11390_, _11389_, _11385_);
  nand _43515_ (_11391_, _11390_, _07271_);
  nand _43516_ (_11392_, _11391_, _11379_);
  nand _43517_ (_11393_, _11392_, _07324_);
  nand _43518_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _11393_, _08053_);
  nand _43519_ (_11394_, _10808_, _07093_);
  nand _43520_ (_11395_, _10813_, _07100_);
  nand _43521_ (_11397_, _11395_, _11394_);
  nand _43522_ (_11398_, _11397_, _07263_);
  nand _43523_ (_11400_, _10824_, _07100_);
  nand _43524_ (_11401_, _10819_, _07093_);
  nand _43525_ (_11402_, _11401_, _11400_);
  nand _43526_ (_11404_, _11402_, _07264_);
  nand _43527_ (_11405_, _11404_, _11398_);
  nand _43528_ (_11406_, _11405_, _07259_);
  nand _43529_ (_11407_, _10847_, _07093_);
  nand _43530_ (_11408_, _10851_, _07100_);
  nand _43531_ (_11409_, _11408_, _11407_);
  nand _43532_ (_11410_, _11409_, _07263_);
  nand _43533_ (_11411_, _10839_, _07100_);
  nand _43534_ (_11412_, _10835_, _07093_);
  nand _43535_ (_11413_, _11412_, _11411_);
  nand _43536_ (_11414_, _11413_, _07264_);
  nand _43537_ (_11416_, _11414_, _11410_);
  nand _43538_ (_11418_, _11416_, _07271_);
  nand _43539_ (_11419_, _11418_, _11406_);
  nand _43540_ (_11421_, _11419_, _07324_);
  nand _43541_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _11421_, _08234_);
  nand _43542_ (_11423_, _10864_, _07093_);
  nand _43543_ (_11424_, _10868_, _07100_);
  nand _43544_ (_11426_, _11424_, _11423_);
  nand _43545_ (_11427_, _11426_, _07263_);
  nand _43546_ (_11429_, _10875_, _07093_);
  nand _43547_ (_11430_, _10880_, _07100_);
  nand _43548_ (_11431_, _11430_, _11429_);
  nand _43549_ (_11432_, _11431_, _07264_);
  nand _43550_ (_11434_, _11432_, _11427_);
  nand _43551_ (_11435_, _11434_, _07259_);
  nand _43552_ (_11436_, _10902_, _07093_);
  nand _43553_ (_11437_, _10907_, _07100_);
  nand _43554_ (_11438_, _11437_, _11436_);
  nand _43555_ (_11439_, _11438_, _07263_);
  nand _43556_ (_11440_, _10894_, _07100_);
  nand _43557_ (_11441_, _10889_, _07093_);
  nand _43558_ (_11443_, _11441_, _11440_);
  nand _43559_ (_11445_, _11443_, _07264_);
  nand _43560_ (_11446_, _11445_, _11439_);
  nand _43561_ (_11447_, _11446_, _07271_);
  nand _43562_ (_11448_, _11447_, _11435_);
  nand _43563_ (_11449_, _11448_, _07324_);
  nand _43564_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _11449_, _08083_);
  nand _43565_ (_11450_, _10923_, _07093_);
  nand _43566_ (_11452_, _10928_, _07100_);
  nand _43567_ (_11454_, _11452_, _11450_);
  nand _43568_ (_11455_, _11454_, _07263_);
  nand _43569_ (_11456_, _10940_, _07100_);
  nand _43570_ (_11457_, _10935_, _07093_);
  nand _43571_ (_11458_, _11457_, _11456_);
  nand _43572_ (_11460_, _11458_, _07264_);
  nand _43573_ (_11462_, _11460_, _11455_);
  nand _43574_ (_11464_, _11462_, _07259_);
  nand _43575_ (_11465_, _10966_, _07093_);
  nand _43576_ (_11467_, _10971_, _07100_);
  nand _43577_ (_11468_, _11467_, _11465_);
  nand _43578_ (_11469_, _11468_, _07263_);
  nand _43579_ (_11470_, _10953_, _07093_);
  nand _43580_ (_11471_, _10958_, _07100_);
  nand _43581_ (_11473_, _11471_, _11470_);
  nand _43582_ (_11474_, _11473_, _07264_);
  nand _43583_ (_11475_, _11474_, _11469_);
  nand _43584_ (_11476_, _11475_, _07271_);
  nand _43585_ (_11477_, _11476_, _11464_);
  nand _43586_ (_11479_, _11477_, _07324_);
  nand _43587_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _11479_, _08101_);
  nand _43588_ (_11480_, _11002_, _07093_);
  nand _43589_ (_11482_, _11007_, _07100_);
  nand _43590_ (_11484_, _11482_, _11480_);
  nand _43591_ (_11485_, _11484_, _07263_);
  nand _43592_ (_11486_, _10988_, _07093_);
  nand _43593_ (_11488_, _10992_, _07100_);
  nand _43594_ (_11490_, _11488_, _11486_);
  nand _43595_ (_11491_, _11490_, _07264_);
  nand _43596_ (_11492_, _11491_, _11485_);
  nand _43597_ (_11494_, _11492_, _07259_);
  nand _43598_ (_11496_, _11033_, _07093_);
  nand _43599_ (_11498_, _11040_, _07100_);
  nand _43600_ (_11500_, _11498_, _11496_);
  nand _43601_ (_11502_, _11500_, _07263_);
  nand _43602_ (_11503_, _11021_, _07100_);
  nand _43603_ (_11505_, _11016_, _07093_);
  nand _43604_ (_11506_, _11505_, _11503_);
  nand _43605_ (_11508_, _11506_, _07264_);
  nand _43606_ (_11510_, _11508_, _11502_);
  nand _43607_ (_11511_, _11510_, _07271_);
  nand _43608_ (_11512_, _11511_, _11494_);
  nand _43609_ (_11513_, _11512_, _07324_);
  nand _43610_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _11513_, _08282_);
  nand _43611_ (_11516_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _43612_ (_11517_, _11516_, _01075_);
  nand _43613_ (_11518_, _11517_, _26487_);
  nand _43614_ (_11520_, _01032_, _25329_);
  nand _43615_ (_11522_, _11520_, _01045_);
  nor _43616_ (_11524_, _11522_, _25421_);
  nand _43617_ (_11526_, _11524_, _01073_);
  nand _43618_ (_11528_, _11526_, _00883_);
  nand _43619_ (_28190_[1], _11528_, _11518_);
  nand _43620_ (_11530_, _10222_, _28096_);
  nand _43621_ (_11531_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nand _43622_ (_03339_, _11531_, _11530_);
  nor _43623_ (_11533_, _00954_, _25159_);
  nand _43624_ (_11534_, _11533_, _24789_);
  not _43625_ (_11535_, _11533_);
  nand _43626_ (_11537_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand _43627_ (_03342_, _11537_, _11534_);
  nand _43628_ (_11540_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  nand _43629_ (_11541_, _08149_, _24830_);
  nand _43630_ (_03379_, _11541_, _11540_);
  nor _43631_ (_11542_, _00415_, _24889_);
  nand _43632_ (_11543_, _11542_, _28096_);
  not _43633_ (_11545_, _11542_);
  nand _43634_ (_11547_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  nand _43635_ (_03386_, _11547_, _11543_);
  nand _43636_ (_11549_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nand _43637_ (_11551_, _08149_, _25039_);
  nand _43638_ (_03401_, _11551_, _11549_);
  nand _43639_ (_11554_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nand _43640_ (_11556_, _25039_, _24796_);
  nand _43641_ (_03403_, _11556_, _11554_);
  nor _43642_ (_11558_, _08142_, _24059_);
  not _43643_ (_11560_, _11558_);
  nand _43644_ (_11562_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  nand _43645_ (_11564_, _11558_, _25039_);
  nand _43646_ (_03406_, _11564_, _11562_);
  nand _43647_ (_11565_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nand _43648_ (_11566_, _11558_, _25099_);
  nand _43649_ (_03419_, _11566_, _11565_);
  nand _43650_ (_11568_, _06437_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _43651_ (_11570_, _06526_, _06458_);
  nor _43652_ (_11571_, _26212_, _26790_);
  nand _43653_ (_11572_, _11571_, _11570_);
  nand _43654_ (_11573_, _00874_, _25329_);
  nor _43655_ (_11575_, _25578_, _25532_);
  nand _43656_ (_11577_, _11575_, _11573_);
  nor _43657_ (_11579_, _11577_, _11572_);
  nand _43658_ (_11581_, _11579_, _25544_);
  nand _43659_ (_11582_, _11581_, _00883_);
  nand _43660_ (_28187_, _11582_, _11568_);
  nand _43661_ (_11583_, _01371_, _24830_);
  nand _43662_ (_11584_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  nand _43663_ (_03425_, _11584_, _11583_);
  nand _43664_ (_11585_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nand _43665_ (_11586_, _08144_, _24830_);
  nand _43666_ (_03430_, _11586_, _11585_);
  nor _43667_ (_11588_, _08142_, _00926_);
  not _43668_ (_11589_, _11588_);
  nand _43669_ (_11590_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  nand _43670_ (_11591_, _11588_, _25099_);
  nand _43671_ (_03435_, _11591_, _11590_);
  nand _43672_ (_11594_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  nand _43673_ (_11595_, _06807_, _25203_);
  nand _43674_ (_03438_, _11595_, _11594_);
  nand _43675_ (_11596_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  nand _43676_ (_11597_, _08144_, _24789_);
  nand _43677_ (_03441_, _11597_, _11596_);
  nand _43678_ (_11599_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  nand _43679_ (_11601_, _11588_, _24789_);
  nand _43680_ (_03448_, _11601_, _11599_);
  nand _43681_ (_11604_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  nand _43682_ (_11606_, _11588_, _25039_);
  nand _43683_ (_03452_, _11606_, _11604_);
  nor _43684_ (_11607_, _00114_, _24073_);
  not _43685_ (_11609_, _11607_);
  nand _43686_ (_11611_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  nand _43687_ (_11612_, _11607_, _25203_);
  nand _43688_ (_03544_, _11612_, _11611_);
  nand _43689_ (_11615_, _00479_, _24927_);
  nand _43690_ (_11616_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  nand _43691_ (_03574_, _11616_, _11615_);
  nor _43692_ (_11619_, _05824_, _25194_);
  not _43693_ (_11621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  nand _43694_ (_11623_, _05824_, _11621_);
  nand _43695_ (_11625_, _11623_, _26487_);
  nor _43696_ (_03580_, _11625_, _11619_);
  nor _43697_ (_11627_, _05824_, _25680_);
  not _43698_ (_11628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nand _43699_ (_11629_, _05824_, _11628_);
  nand _43700_ (_11631_, _11629_, _26487_);
  nor _43701_ (_03590_, _11631_, _11627_);
  nor _43702_ (_11633_, _00114_, _28057_);
  nand _43703_ (_11634_, _11633_, _28096_);
  not _43704_ (_11636_, _11633_);
  nand _43705_ (_11637_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nand _43706_ (_03594_, _11637_, _11634_);
  nor _43707_ (_11638_, _28104_, _24882_);
  nand _43708_ (_11639_, _11638_, _25099_);
  not _43709_ (_11640_, _11638_);
  nand _43710_ (_11642_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nand _43711_ (_03606_, _11642_, _11639_);
  nand _43712_ (_11643_, _04624_, _25039_);
  nand _43713_ (_11644_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  nand _43714_ (_03608_, _11644_, _11643_);
  nand _43715_ (_11646_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  nand _43716_ (_11647_, _11588_, _25203_);
  nand _43717_ (_03610_, _11647_, _11646_);
  nand _43718_ (_11648_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  nand _43719_ (_11649_, _11588_, _28096_);
  nand _43720_ (_03622_, _11649_, _11648_);
  nand _43721_ (_11652_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  nand _43722_ (_11654_, _03547_, _24789_);
  nand _43723_ (_03625_, _11654_, _11652_);
  nand _43724_ (_11657_, _01402_, _25150_);
  nand _43725_ (_11658_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nand _43726_ (_03636_, _11658_, _11657_);
  nor _43727_ (_11659_, _00629_, _28104_);
  nand _43728_ (_11660_, _11659_, _25150_);
  not _43729_ (_11661_, _11659_);
  nand _43730_ (_11662_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  nand _43731_ (_03648_, _11662_, _11660_);
  nand _43732_ (_11663_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  nand _43733_ (_11665_, _11607_, _24830_);
  nand _43734_ (_03661_, _11665_, _11663_);
  nand _43735_ (_11666_, _04624_, _25203_);
  nand _43736_ (_11668_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  nand _43737_ (_03663_, _11668_, _11666_);
  nand _43738_ (_11669_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  nand _43739_ (_11670_, _11607_, _25150_);
  nand _43740_ (_03677_, _11670_, _11669_);
  nand _43741_ (_11671_, _03446_, _25099_);
  nand _43742_ (_11672_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nand _43743_ (_03681_, _11672_, _11671_);
  nand _43744_ (_11673_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  nand _43745_ (_11674_, _11588_, _25150_);
  nand _43746_ (_03683_, _11674_, _11673_);
  nand _43747_ (_11675_, _09944_, _24789_);
  nand _43748_ (_11676_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  nand _43749_ (_03696_, _11676_, _11675_);
  nand _43750_ (_11677_, _07742_, _04181_);
  nor _43751_ (_11678_, _04192_, _07747_);
  nand _43752_ (_11679_, _11678_, _11677_);
  nor _43753_ (_11680_, _07728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _43754_ (_11681_, _07730_, _01617_);
  nor _43755_ (_11682_, _11681_, _11680_);
  nor _43756_ (_11683_, _09321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _43757_ (_11684_, _07736_, _01574_);
  nor _43758_ (_11685_, _11684_, _11683_);
  nor _43759_ (_11686_, _11685_, _11682_);
  nand _43760_ (_11687_, _11686_, _11679_);
  nand _43761_ (_11688_, _11687_, _01642_);
  nand _43762_ (_11690_, _01644_, _25194_);
  nand _43763_ (_11692_, _11690_, _11688_);
  nor _43764_ (_11693_, _11692_, _01573_);
  nand _43765_ (_11694_, _01573_, _04181_);
  nand _43766_ (_11695_, _11694_, _26487_);
  nor _43767_ (_03700_, _11695_, _11693_);
  nand _43768_ (_11696_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  nand _43769_ (_11697_, _11607_, _24927_);
  nand _43770_ (_03712_, _11697_, _11696_);
  nand _43771_ (_11698_, _11638_, _25203_);
  nand _43772_ (_11699_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  nand _43773_ (_03721_, _11699_, _11698_);
  nand _43774_ (_11700_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  nand _43775_ (_11701_, _11588_, _24927_);
  nand _43776_ (_03723_, _11701_, _11700_);
  nor _43777_ (_11702_, _05824_, _25089_);
  nand _43778_ (_11703_, _05824_, _01609_);
  nand _43779_ (_11705_, _11703_, _26487_);
  nor _43780_ (_03730_, _11705_, _11702_);
  nand _43781_ (_11706_, _11638_, _24927_);
  nand _43782_ (_11708_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  nand _43783_ (_03733_, _11708_, _11706_);
  nand _43784_ (_11711_, _03850_, _24927_);
  nand _43785_ (_11713_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  nand _43786_ (_03745_, _11713_, _11711_);
  nand _43787_ (_11716_, _11638_, _24789_);
  nand _43788_ (_11718_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  nand _43789_ (_03747_, _11718_, _11716_);
  nor _43790_ (_11720_, _00393_, _28104_);
  nand _43791_ (_11722_, _11720_, _24830_);
  not _43792_ (_11724_, _11720_);
  nand _43793_ (_11726_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  nand _43794_ (_03754_, _11726_, _11722_);
  nand _43795_ (_11729_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  nand _43796_ (_11731_, _11607_, _24789_);
  nand _43797_ (_03758_, _11731_, _11729_);
  nand _43798_ (_11734_, _00979_, _24927_);
  nand _43799_ (_11736_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  nand _43800_ (_03776_, _11736_, _11734_);
  nor _43801_ (_11738_, _25165_, _24795_);
  nand _43802_ (_11739_, _11738_, _25039_);
  not _43803_ (_11741_, _11738_);
  nand _43804_ (_11742_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  nand _43805_ (_03784_, _11742_, _11739_);
  not _43806_ (_11744_, _01073_);
  not _43807_ (_11745_, _11573_);
  nor _43808_ (_11746_, _11745_, _11744_);
  nor _43809_ (_11747_, _11746_, _25530_);
  not _43810_ (_11749_, _06664_);
  nor _43811_ (_11750_, _01074_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _43812_ (_11751_, _11750_, _11749_);
  nor _43813_ (_11753_, _11751_, _11747_);
  nand _43814_ (_11755_, _24100_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _43815_ (_11756_, _11755_, _26487_);
  nor _43816_ (_28191_[2], _11756_, _11753_);
  nand _43817_ (_11758_, _11738_, _25203_);
  nand _43818_ (_11759_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nand _43819_ (_03799_, _11759_, _11758_);
  nand _43820_ (_11761_, _03850_, _25039_);
  nand _43821_ (_11762_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  nand _43822_ (_03802_, _11762_, _11761_);
  nand _43823_ (_11764_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nand _43824_ (_11765_, _08144_, _25150_);
  nand _43825_ (_03821_, _11765_, _11764_);
  nand _43826_ (_11767_, _11738_, _28096_);
  nand _43827_ (_11769_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  nand _43828_ (_03823_, _11769_, _11767_);
  nand _43829_ (_11770_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  nand _43830_ (_11771_, _08144_, _24927_);
  nand _43831_ (_03833_, _11771_, _11770_);
  nor _43832_ (_11772_, _00926_, _25165_);
  nand _43833_ (_11774_, _11772_, _24830_);
  not _43834_ (_11776_, _11772_);
  nand _43835_ (_11778_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  nand _43836_ (_03860_, _11778_, _11774_);
  nor _43837_ (_11781_, _07814_, _24016_);
  nand _43838_ (_11782_, _25156_, _11781_);
  nor _43839_ (_11783_, _11782_, _24978_);
  nand _43840_ (_11784_, _11783_, _24830_);
  not _43841_ (_11785_, _11783_);
  nand _43842_ (_11786_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nand _43843_ (_03863_, _11786_, _11784_);
  nand _43844_ (_11787_, _11783_, _24927_);
  nand _43845_ (_11788_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  nand _43846_ (_03864_, _11788_, _11787_);
  nand _43847_ (_11789_, _11783_, _25150_);
  nand _43848_ (_11790_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  nand _43849_ (_03875_, _11790_, _11789_);
  nand _43850_ (_11791_, _01371_, _25099_);
  nand _43851_ (_11792_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  nand _43852_ (_03885_, _11792_, _11791_);
  nand _43853_ (_11793_, _11738_, _24789_);
  nand _43854_ (_11794_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  nand _43855_ (_03887_, _11794_, _11793_);
  nor _43856_ (_11795_, _01260_, _05327_);
  nand _43857_ (_11796_, _01253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _43858_ (_11797_, _11796_, _01261_);
  nor _43859_ (_11798_, _11797_, _11795_);
  nor _43860_ (_03899_, _11798_, rst);
  nand _43861_ (_11800_, _11738_, _25150_);
  nand _43862_ (_11802_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nand _43863_ (_03901_, _11802_, _11800_);
  nor _43864_ (_11805_, _05775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _43865_ (_11807_, _05076_, _00259_);
  nor _43866_ (_11809_, _11807_, _05779_);
  not _43867_ (_11811_, _11809_);
  nor _43868_ (_11813_, _11811_, _11805_);
  nor _43869_ (_11815_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _43870_ (_11818_, _11815_, _11813_);
  nor _43871_ (_11820_, _11818_, _11813_);
  nor _43872_ (_11822_, _11820_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _43873_ (_11824_, _11818_, _05730_);
  nand _43874_ (_11826_, _11824_, _26487_);
  nor _43875_ (_03909_, _11826_, _11822_);
  nor _43876_ (_11827_, _00926_, _00631_);
  nand _43877_ (_11828_, _11827_, _25039_);
  not _43878_ (_11829_, _11827_);
  nand _43879_ (_11831_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nand _43880_ (_03922_, _11831_, _11828_);
  nand _43881_ (_11834_, _11738_, _24927_);
  nand _43882_ (_11835_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  nand _43883_ (_03927_, _11835_, _11834_);
  nand _43884_ (_11836_, _07670_, _25039_);
  nand _43885_ (_11837_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  nand _43886_ (_03941_, _11837_, _11836_);
  nor _43887_ (_11839_, _28104_, _28080_);
  nand _43888_ (_11840_, _11839_, _24927_);
  not _43889_ (_11841_, _11839_);
  nand _43890_ (_11842_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  nand _43891_ (_03950_, _11842_, _11840_);
  nand _43892_ (_11843_, _11589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  nand _43893_ (_11844_, _11588_, _24830_);
  nand _43894_ (_03963_, _11844_, _11843_);
  nand _43895_ (_11845_, _11839_, _24830_);
  nand _43896_ (_11846_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  nand _43897_ (_03965_, _11846_, _11845_);
  nor _43898_ (_11848_, _28104_, _28073_);
  nand _43899_ (_11849_, _11848_, _25039_);
  not _43900_ (_11850_, _11848_);
  nand _43901_ (_11852_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  nand _43902_ (_03970_, _11852_, _11849_);
  nand _43903_ (_11853_, _11848_, _28096_);
  nand _43904_ (_11854_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  nand _43905_ (_03972_, _11854_, _11853_);
  nor _43906_ (_11855_, _00122_, _28104_);
  nand _43907_ (_11856_, _11855_, _24927_);
  not _43908_ (_11857_, _11855_);
  nand _43909_ (_11858_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  nand _43910_ (_03982_, _11858_, _11856_);
  nand _43911_ (_11859_, _11855_, _25203_);
  nand _43912_ (_11861_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  nand _43913_ (_03984_, _11861_, _11859_);
  nor _43914_ (_11862_, _25165_, _24059_);
  nand _43915_ (_11863_, _11862_, _25039_);
  not _43916_ (_11864_, _11862_);
  nand _43917_ (_11865_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nand _43918_ (_03993_, _11865_, _11863_);
  nor _43919_ (_11867_, _28104_, _25047_);
  nand _43920_ (_11869_, _11867_, _24927_);
  not _43921_ (_11870_, _11867_);
  nand _43922_ (_11871_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  nand _43923_ (_03996_, _11871_, _11869_);
  nand _43924_ (_11872_, _11867_, _25203_);
  nand _43925_ (_11873_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  nand _43926_ (_03997_, _11873_, _11872_);
  nor _43927_ (_11874_, _00415_, _28104_);
  nand _43928_ (_11875_, _11874_, _25150_);
  not _43929_ (_11876_, _11874_);
  nand _43930_ (_11877_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  nand _43931_ (_04002_, _11877_, _11875_);
  nand _43932_ (_11879_, _11874_, _25039_);
  nand _43933_ (_11880_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nand _43934_ (_04004_, _11880_, _11879_);
  nand _43935_ (_11882_, _11862_, _24927_);
  nand _43936_ (_11884_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  nand _43937_ (_04010_, _11884_, _11882_);
  nor _43938_ (_11886_, _23870_, _24077_);
  nand _43939_ (_11887_, _11886_, _26487_);
  nand _43940_ (_11889_, _01048_, _25391_);
  nor _43941_ (_11891_, _04965_, _01050_);
  nand _43942_ (_11892_, _11891_, _11889_);
  nand _43943_ (_11894_, _06524_, _04969_);
  nor _43944_ (_11895_, _11894_, _11892_);
  nor _43945_ (_11896_, _26202_, _25490_);
  nand _43946_ (_11898_, _06441_, _04282_);
  nor _43947_ (_11899_, _11898_, _11896_);
  nor _43948_ (_11900_, _04953_, _25566_);
  nand _43949_ (_11901_, _11900_, _11899_);
  nor _43950_ (_11902_, _06557_, _25491_);
  nand _43951_ (_11903_, _11902_, _06543_);
  nor _43952_ (_11904_, _11903_, _11901_);
  nand _43953_ (_11905_, _11904_, _11895_);
  nand _43954_ (_11906_, _11905_, _00883_);
  nand _43955_ (_28193_[3], _11906_, _11887_);
  nor _43956_ (_11907_, _00954_, _28104_);
  nand _43957_ (_11908_, _11907_, _25203_);
  not _43958_ (_11909_, _11907_);
  nand _43959_ (_11910_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nand _43960_ (_04029_, _11910_, _11908_);
  nand _43961_ (_11911_, _11827_, _25203_);
  nand _43962_ (_11912_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nand _43963_ (_04032_, _11912_, _11911_);
  nand _43964_ (_11913_, _11720_, _25039_);
  nand _43965_ (_11914_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nand _43966_ (_04039_, _11914_, _11913_);
  nand _43967_ (_11915_, _11659_, _28096_);
  nand _43968_ (_11916_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nand _43969_ (_04049_, _11916_, _11915_);
  nand _43970_ (_11917_, _11659_, _24830_);
  nand _43971_ (_11918_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  nand _43972_ (_04051_, _11918_, _11917_);
  nor _43973_ (_11919_, _00114_, _28104_);
  nand _43974_ (_11920_, _11919_, _24789_);
  not _43975_ (_11921_, _11919_);
  nand _43976_ (_11922_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  nand _43977_ (_04064_, _11922_, _11920_);
  nand _43978_ (_11923_, _11919_, _25203_);
  nand _43979_ (_11924_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  nand _43980_ (_04073_, _11924_, _11923_);
  nand _43981_ (_11925_, _11919_, _25099_);
  nand _43982_ (_11926_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nand _43983_ (_04075_, _11926_, _11925_);
  nand _43984_ (_11927_, _11862_, _24789_);
  nand _43985_ (_11928_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  nand _43986_ (_04077_, _11928_, _11927_);
  nand _43987_ (_11929_, _11738_, _24830_);
  nand _43988_ (_11930_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  nand _43989_ (_04092_, _11930_, _11929_);
  nor _43990_ (_11931_, _11782_, _00926_);
  nand _43991_ (_11932_, _11931_, _25039_);
  not _43992_ (_11933_, _11931_);
  nand _43993_ (_11934_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nand _43994_ (_04100_, _11934_, _11932_);
  nand _43995_ (_11935_, _11931_, _28096_);
  nand _43996_ (_11936_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nand _43997_ (_04102_, _11936_, _11935_);
  nor _43998_ (_11937_, _11782_, _24795_);
  nand _43999_ (_11938_, _11937_, _24927_);
  not _44000_ (_11939_, _11937_);
  nand _44001_ (_11940_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  nand _44002_ (_04108_, _11940_, _11938_);
  nand _44003_ (_11941_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  nand _44004_ (_11942_, _11558_, _24789_);
  nand _44005_ (_04112_, _11942_, _11941_);
  nand _44006_ (_11943_, _11937_, _25203_);
  nand _44007_ (_11944_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  nand _44008_ (_04115_, _11944_, _11943_);
  nand _44009_ (_11945_, _11638_, _25039_);
  nand _44010_ (_11946_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nand _44011_ (_04124_, _11946_, _11945_);
  nand _44012_ (_11947_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  nand _44013_ (_11948_, _11558_, _25150_);
  nand _44014_ (_04126_, _11948_, _11947_);
  nand _44015_ (_11949_, _11638_, _24830_);
  nand _44016_ (_11950_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  nand _44017_ (_04128_, _11950_, _11949_);
  nand _44018_ (_11951_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  nand _44019_ (_11952_, _11558_, _24927_);
  nand _44020_ (_04135_, _11952_, _11951_);
  nand _44021_ (_11953_, _11659_, _24789_);
  nand _44022_ (_11954_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  nand _44023_ (_04137_, _11954_, _11953_);
  nand _44024_ (_11955_, _11638_, _28096_);
  nand _44025_ (_11956_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  nand _44026_ (_04143_, _11956_, _11955_);
  nand _44027_ (_11957_, _07670_, _25099_);
  nand _44028_ (_11958_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nand _44029_ (_04147_, _11958_, _11957_);
  nand _44030_ (_11959_, _11839_, _28096_);
  nand _44031_ (_11960_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  nand _44032_ (_04161_, _11960_, _11959_);
  not _44033_ (_11961_, _04591_);
  nand _44034_ (_11962_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nand _44035_ (_04164_, _11962_, _11961_);
  nand _44036_ (_11963_, _11848_, _25150_);
  nand _44037_ (_11964_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  nand _44038_ (_04179_, _11964_, _11963_);
  nand _44039_ (_11966_, _11855_, _24789_);
  nand _44040_ (_11967_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  nand _44041_ (_04184_, _11967_, _11966_);
  nand _44042_ (_11968_, _11783_, _25039_);
  nand _44043_ (_11969_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nand _44044_ (_04190_, _11969_, _11968_);
  nand _44045_ (_11971_, _11867_, _24789_);
  nand _44046_ (_11972_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  nand _44047_ (_04197_, _11972_, _11971_);
  nor _44048_ (_11973_, _11782_, _24059_);
  nand _44049_ (_11974_, _11973_, _25039_);
  not _44050_ (_11975_, _11973_);
  nand _44051_ (_11976_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  nand _44052_ (_04200_, _11976_, _11974_);
  nand _44053_ (_11977_, _11973_, _25099_);
  nand _44054_ (_11978_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nand _44055_ (_04202_, _11978_, _11977_);
  nand _44056_ (_11979_, _11874_, _24830_);
  nand _44057_ (_11980_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  nand _44058_ (_04211_, _11980_, _11979_);
  nand _44059_ (_11981_, _11907_, _24927_);
  nand _44060_ (_11982_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  nand _44061_ (_04213_, _11982_, _11981_);
  nand _44062_ (_11983_, _11907_, _25099_);
  nand _44063_ (_11984_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  nand _44064_ (_04216_, _11984_, _11983_);
  nand _44065_ (_11985_, _11720_, _25150_);
  nand _44066_ (_11986_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  nand _44067_ (_04218_, _11986_, _11985_);
  nand _44068_ (_11987_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nand _44069_ (_11988_, _08144_, _28096_);
  nand _44070_ (_04224_, _11988_, _11987_);
  nand _44071_ (_11989_, _11659_, _25039_);
  nand _44072_ (_11990_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  nand _44073_ (_04227_, _11990_, _11989_);
  nand _44074_ (_11991_, _11919_, _24927_);
  nand _44075_ (_11992_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  nand _44076_ (_04229_, _11992_, _11991_);
  nand _44077_ (_11993_, _11973_, _28096_);
  nand _44078_ (_11994_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  nand _44079_ (_04239_, _11994_, _11993_);
  nand _44080_ (_11995_, _11931_, _25150_);
  nand _44081_ (_11996_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  nand _44082_ (_04241_, _11996_, _11995_);
  nand _44083_ (_11997_, _11937_, _24789_);
  nand _44084_ (_11998_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  nand _44085_ (_04260_, _11998_, _11997_);
  nand _44086_ (_11999_, _11937_, _24830_);
  nand _44087_ (_12000_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  nand _44088_ (_04263_, _12000_, _11999_);
  nand _44089_ (_12001_, _11720_, _25099_);
  nand _44090_ (_12002_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nand _44091_ (_04268_, _12002_, _12001_);
  nand _44092_ (_12003_, _11638_, _25150_);
  nand _44093_ (_12004_, _11640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nand _44094_ (_04272_, _12004_, _12003_);
  nand _44095_ (_12005_, _07670_, _24927_);
  nand _44096_ (_12006_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  nand _44097_ (_04278_, _12006_, _12005_);
  nand _44098_ (_12008_, _11839_, _25150_);
  nand _44099_ (_12009_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nand _44100_ (_04281_, _12009_, _12008_);
  nor _44101_ (_12010_, _28057_, _28080_);
  nand _44102_ (_12011_, _12010_, _24830_);
  not _44103_ (_12012_, _12010_);
  nand _44104_ (_12013_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nand _44105_ (_04284_, _12013_, _12011_);
  nand _44106_ (_12014_, _11973_, _24927_);
  nand _44107_ (_12015_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  nand _44108_ (_04287_, _12015_, _12014_);
  nand _44109_ (_12016_, _08146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  nand _44110_ (_12017_, _08144_, _25099_);
  nand _44111_ (_04294_, _12017_, _12016_);
  nand _44112_ (_12018_, _11867_, _24830_);
  nand _44113_ (_12019_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  nand _44114_ (_04295_, _12019_, _12018_);
  nand _44115_ (_12020_, _11973_, _25150_);
  nand _44116_ (_12021_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  nand _44117_ (_04297_, _12021_, _12020_);
  not _44118_ (_12022_, _01430_);
  nand _44119_ (_12023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _03739_);
  nor _44120_ (_12024_, _12023_, _12022_);
  nand _44121_ (_12025_, _01429_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not _44122_ (_12027_, _01436_);
  nand _44123_ (_12028_, _12027_, _01431_);
  nand _44124_ (_12029_, _01433_, _01241_);
  nand _44125_ (_12030_, _12029_, _12028_);
  nand _44126_ (_12031_, _12030_, _12025_);
  nor _44127_ (_12032_, _12031_, _12024_);
  nor _44128_ (_04300_, _12032_, _01460_);
  nand _44129_ (_12034_, _11973_, _24830_);
  nand _44130_ (_12035_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nand _44131_ (_04330_, _12035_, _12034_);
  nand _44132_ (_12036_, _11848_, _24789_);
  nand _44133_ (_12037_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  nand _44134_ (_04334_, _12037_, _12036_);
  nor _44135_ (_12038_, _11782_, _00114_);
  nand _44136_ (_12039_, _12038_, _25203_);
  not _44137_ (_12040_, _12038_);
  nand _44138_ (_12041_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  nand _44139_ (_04339_, _12041_, _12039_);
  nand _44140_ (_12043_, _11874_, _25099_);
  nand _44141_ (_12044_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  nand _44142_ (_04343_, _12044_, _12043_);
  nand _44143_ (_12045_, _11659_, _24927_);
  nand _44144_ (_12046_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  nand _44145_ (_04345_, _12046_, _12045_);
  nand _44146_ (_12047_, _11931_, _24789_);
  nand _44147_ (_12048_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nand _44148_ (_04349_, _12048_, _12047_);
  nand _44149_ (_12049_, _12038_, _28096_);
  nand _44150_ (_12050_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nand _44151_ (_04351_, _12050_, _12049_);
  nand _44152_ (_12051_, _11720_, _28096_);
  nand _44153_ (_12052_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  nand _44154_ (_04353_, _12052_, _12051_);
  nand _44155_ (_12053_, _07670_, _25150_);
  nand _44156_ (_12054_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  nand _44157_ (_04355_, _12054_, _12053_);
  nand _44158_ (_12055_, _11855_, _24830_);
  nand _44159_ (_12056_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  nand _44160_ (_04357_, _12056_, _12055_);
  nand _44161_ (_12058_, _11937_, _25099_);
  nand _44162_ (_12059_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  nand _44163_ (_04359_, _12059_, _12058_);
  nand _44164_ (_12060_, _12038_, _25099_);
  nand _44165_ (_12061_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  nand _44166_ (_04361_, _12061_, _12060_);
  nor _44167_ (_12062_, _04173_, _24782_);
  nand _44168_ (_12063_, _04233_, _01609_);
  nor _44169_ (_12064_, _12063_, _07998_);
  nand _44170_ (_12066_, _12063_, _07998_);
  nand _44171_ (_12067_, _12066_, _01617_);
  nor _44172_ (_12068_, _12067_, _12064_);
  nand _44173_ (_12069_, _04194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _44174_ (_12070_, _12069_, _07998_);
  nor _44175_ (_12072_, _12069_, _07998_);
  nor _44176_ (_12073_, _12072_, _07747_);
  nand _44177_ (_12074_, _12073_, _12070_);
  nand _44178_ (_12076_, _04207_, _07998_);
  nor _44179_ (_12077_, _08000_, _01597_);
  nor _44180_ (_12078_, _12077_, _04208_);
  nand _44181_ (_12079_, _12078_, _12076_);
  nand _44182_ (_12080_, _12079_, _12074_);
  nor _44183_ (_12081_, _12080_, _12068_);
  nand _44184_ (_12083_, _12081_, _04173_);
  nand _44185_ (_12084_, _12083_, _04175_);
  nor _44186_ (_12085_, _12084_, _12062_);
  nor _44187_ (_12086_, _04175_, _07998_);
  nor _44188_ (_12088_, _12086_, _12085_);
  nor _44189_ (_04365_, _12088_, rst);
  nor _44190_ (_12089_, _25165_, _24999_);
  nand _44191_ (_12090_, _12089_, _28096_);
  not _44192_ (_12092_, _12089_);
  nand _44193_ (_12093_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  nand _44194_ (_04368_, _12093_, _12090_);
  nand _44195_ (_12094_, _03850_, _24789_);
  nand _44196_ (_12095_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  nand _44197_ (_04374_, _12095_, _12094_);
  nor _44198_ (_12096_, _00122_, _25165_);
  nand _44199_ (_12097_, _12096_, _24927_);
  not _44200_ (_12098_, _12096_);
  nand _44201_ (_12099_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  nand _44202_ (_04381_, _12099_, _12097_);
  nor _44203_ (_12100_, _25165_, _25047_);
  nand _44204_ (_12101_, _12100_, _28096_);
  not _44205_ (_12102_, _12100_);
  nand _44206_ (_12103_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  nand _44207_ (_04388_, _12103_, _12101_);
  nor _44208_ (_12104_, _00415_, _25165_);
  nand _44209_ (_12105_, _12104_, _25203_);
  not _44210_ (_12107_, _12104_);
  nand _44211_ (_12108_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  nand _44212_ (_04404_, _12108_, _12105_);
  nand _44213_ (_12109_, _06826_, _25039_);
  nand _44214_ (_12110_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  nand _44215_ (_04406_, _12110_, _12109_);
  nand _44216_ (_12112_, _03876_, _24927_);
  nand _44217_ (_12114_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  nand _44218_ (_04408_, _12114_, _12112_);
  nand _44219_ (_12116_, _12038_, _25150_);
  nand _44220_ (_12117_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  nand _44221_ (_04414_, _12117_, _12116_);
  nand _44222_ (_12118_, _00115_, _25039_);
  nand _44223_ (_12120_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  nand _44224_ (_04417_, _12120_, _12118_);
  nand _44225_ (_12122_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  nand _44226_ (_12123_, _01388_, _24789_);
  nand _44227_ (_04422_, _12123_, _12122_);
  nand _44228_ (_12124_, _12038_, _24927_);
  nand _44229_ (_12125_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  nand _44230_ (_04432_, _12125_, _12124_);
  nand _44231_ (_12127_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  nand _44232_ (_12128_, _11558_, _24830_);
  nand _44233_ (_04433_, _12128_, _12127_);
  nand _44234_ (_12129_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  nand _44235_ (_12131_, _00330_, _24830_);
  nand _44236_ (_04436_, _12131_, _12129_);
  nand _44237_ (_12132_, _12038_, _25039_);
  nand _44238_ (_12133_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  nand _44239_ (_04438_, _12133_, _12132_);
  nand _44240_ (_12134_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  nand _44241_ (_12135_, _00408_, _28096_);
  nand _44242_ (_04439_, _12135_, _12134_);
  nand _44243_ (_12136_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nand _44244_ (_12137_, _00636_, _25039_);
  nand _44245_ (_04441_, _12137_, _12136_);
  nand _44246_ (_12138_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  nand _44247_ (_12139_, _01174_, _25150_);
  nand _44248_ (_04448_, _12139_, _12138_);
  nand _44249_ (_12140_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  nand _44250_ (_12141_, _03547_, _25150_);
  nand _44251_ (_04463_, _12141_, _12140_);
  nand _44252_ (_12142_, _11772_, _25203_);
  nand _44253_ (_12143_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  nand _44254_ (_04469_, _12143_, _12142_);
  nand _44255_ (_12144_, _03830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  nand _44256_ (_12145_, _03829_, _28096_);
  nand _44257_ (_04472_, _12145_, _12144_);
  nand _44258_ (_12146_, _11772_, _24927_);
  nand _44259_ (_12147_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  nand _44260_ (_04474_, _12147_, _12146_);
  nor _44261_ (_12148_, _04175_, _25680_);
  not _44262_ (_12149_, _07561_);
  nor _44263_ (_12150_, _12149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _44264_ (_12151_, _12150_, _07562_);
  nor _44265_ (_12152_, _07637_, _04182_);
  nor _44266_ (_12153_, _12152_, _12151_);
  nor _44267_ (_12154_, _12153_, _01644_);
  nor _44268_ (_12155_, _01642_, _07558_);
  nor _44269_ (_12156_, _12155_, _12154_);
  nand _44270_ (_12157_, _12156_, _04175_);
  nand _44271_ (_12158_, _12157_, _26487_);
  nor _44272_ (_04481_, _12158_, _12148_);
  nand _44273_ (_12159_, _11772_, _25039_);
  nand _44274_ (_12160_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nand _44275_ (_04483_, _12160_, _12159_);
  nand _44276_ (_12161_, _09547_, _25150_);
  nand _44277_ (_12162_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nand _44278_ (_04489_, _12162_, _12161_);
  nand _44279_ (_12163_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  nand _44280_ (_12164_, _04299_, _28096_);
  nand _44281_ (_04501_, _12164_, _12163_);
  nand _44282_ (_12165_, _09547_, _24927_);
  nand _44283_ (_12166_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  nand _44284_ (_04504_, _12166_, _12165_);
  nand _44285_ (_12167_, _08354_, _28096_);
  nand _44286_ (_12168_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nand _44287_ (_04507_, _12168_, _12167_);
  nand _44288_ (_12169_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  nand _44289_ (_12170_, _11558_, _28096_);
  nand _44290_ (_04512_, _12170_, _12169_);
  nand _44291_ (_12171_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nand _44292_ (_12172_, _05735_, _24830_);
  nand _44293_ (_04516_, _12172_, _12171_);
  nand _44294_ (_12173_, _28096_, _24890_);
  nand _44295_ (_12174_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nand _44296_ (_04519_, _12174_, _12173_);
  nand _44297_ (_12175_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  nand _44298_ (_12176_, _05847_, _24927_);
  nand _44299_ (_04527_, _12176_, _12175_);
  nand _44300_ (_12177_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  nand _44301_ (_12178_, _05864_, _25203_);
  nand _44302_ (_04535_, _12178_, _12177_);
  nand _44303_ (_12179_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  nand _44304_ (_12180_, _05864_, _24830_);
  nand _44305_ (_04540_, _12180_, _12179_);
  nand _44306_ (_12181_, _11560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nand _44307_ (_12182_, _11558_, _25203_);
  nand _44308_ (_04551_, _12182_, _12181_);
  nand _44309_ (_12183_, _11772_, _24789_);
  nand _44310_ (_12184_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  nand _44311_ (_04565_, _12184_, _12183_);
  nand _44312_ (_12185_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  nand _44313_ (_12186_, _11607_, _25039_);
  nand _44314_ (_04568_, _12186_, _12185_);
  nor _44315_ (_12187_, _24768_, _26812_);
  nand _44316_ (_12188_, _12187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44317_ (_12189_, _12187_);
  nand _44318_ (_12190_, _12189_, _26816_);
  nand _44319_ (_12191_, _12190_, _12188_);
  nor _44320_ (_04572_, _12191_, rst);
  nor _44321_ (_04574_, _02791_, rst);
  nor _44322_ (_04578_, _27087_, rst);
  nand _44323_ (_12192_, _03911_, _25039_);
  nand _44324_ (_12193_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  nand _44325_ (_04582_, _12193_, _12192_);
  nand _44326_ (_12194_, _25166_, _24830_);
  nand _44327_ (_12195_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  nand _44328_ (_04593_, _12195_, _12194_);
  nand _44329_ (_12196_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nand _44330_ (_12197_, _25150_, _24074_);
  nand _44331_ (_04595_, _12197_, _12196_);
  nand _44332_ (_12198_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nand _44333_ (_12199_, _00843_, _25039_);
  nand _44334_ (_04605_, _12199_, _12198_);
  nand _44335_ (_12200_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  nand _44336_ (_12201_, _01129_, _25203_);
  nand _44337_ (_04612_, _12201_, _12200_);
  nor _44338_ (_12202_, _07560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _44339_ (_12203_, _12202_, _12149_);
  nand _44340_ (_12204_, _01614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _44341_ (_12205_, _12204_, _01632_);
  nor _44342_ (_12206_, _12205_, _12203_);
  nor _44343_ (_12207_, _12206_, _01644_);
  nor _44344_ (_12208_, _01642_, _01588_);
  nor _44345_ (_12209_, _12208_, _12207_);
  nor _44346_ (_12210_, _12209_, _01573_);
  nor _44347_ (_12211_, _04175_, _25088_);
  nor _44348_ (_12212_, _12211_, _12210_);
  nor _44349_ (_04619_, _12212_, rst);
  nand _44350_ (_12213_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  nand _44351_ (_12214_, _04166_, _24789_);
  nand _44352_ (_04636_, _12214_, _12213_);
  nand _44353_ (_12215_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nand _44354_ (_12216_, _04255_, _25039_);
  nand _44355_ (_04641_, _12216_, _12215_);
  nand _44356_ (_12217_, _11772_, _25099_);
  nand _44357_ (_12218_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nand _44358_ (_04645_, _12218_, _12217_);
  nand _44359_ (_12219_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nand _44360_ (_12220_, _08149_, _25203_);
  nand _44361_ (_04649_, _12220_, _12219_);
  nand _44362_ (_12221_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  nand _44363_ (_12222_, _04322_, _25203_);
  nand _44364_ (_04651_, _12222_, _12221_);
  nand _44365_ (_12223_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nand _44366_ (_12224_, _08149_, _28096_);
  nand _44367_ (_04658_, _12224_, _12223_);
  nand _44368_ (_12225_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nand _44369_ (_12226_, _08149_, _25099_);
  nand _44370_ (_04661_, _12226_, _12225_);
  nand _44371_ (_12227_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  nand _44372_ (_12228_, _05864_, _24789_);
  nand _44373_ (_04663_, _12228_, _12227_);
  nand _44374_ (_12229_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nand _44375_ (_12230_, _05847_, _25099_);
  nand _44376_ (_04665_, _12230_, _12229_);
  nand _44377_ (_12231_, _11633_, _24927_);
  nand _44378_ (_12232_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  nand _44379_ (_04674_, _12232_, _12231_);
  nor _44380_ (_04677_, _07953_, rst);
  nand _44381_ (_12233_, _12104_, _25039_);
  nand _44382_ (_12234_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  nand _44383_ (_04688_, _12234_, _12233_);
  nor _44384_ (_12235_, _25165_, _24978_);
  nand _44385_ (_12236_, _12235_, _25099_);
  not _44386_ (_12237_, _12235_);
  nand _44387_ (_12238_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nand _44388_ (_04691_, _12238_, _12236_);
  nand _44389_ (_12239_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  nand _44390_ (_12240_, _01388_, _24830_);
  nand _44391_ (_04699_, _12240_, _12239_);
  nand _44392_ (_12241_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nand _44393_ (_12242_, _00330_, _25099_);
  nand _44394_ (_04705_, _12242_, _12241_);
  nand _44395_ (_12243_, _12235_, _24830_);
  nand _44396_ (_12244_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nand _44397_ (_04709_, _12244_, _12243_);
  nand _44398_ (_12245_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nand _44399_ (_12246_, _08149_, _24927_);
  nand _44400_ (_04735_, _12246_, _12245_);
  nand _44401_ (_12247_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nand _44402_ (_12248_, _04299_, _25203_);
  nand _44403_ (_04741_, _12248_, _12247_);
  nand _44404_ (_12249_, _08150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nand _44405_ (_12250_, _08149_, _25150_);
  nand _44406_ (_04743_, _12250_, _12249_);
  nand _44407_ (_12251_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nand _44408_ (_12252_, _06807_, _25099_);
  nand _44409_ (_04748_, _12252_, _12251_);
  nand _44410_ (_12254_, _12235_, _24927_);
  nand _44411_ (_12255_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  nand _44412_ (_04758_, _12255_, _12254_);
  nand _44413_ (_12256_, _12235_, _25039_);
  nand _44414_ (_12257_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nand _44415_ (_04765_, _12257_, _12256_);
  nand _44416_ (_12258_, _12235_, _25203_);
  nand _44417_ (_12259_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  nand _44418_ (_04798_, _12259_, _12258_);
  nor _44419_ (_12260_, _11782_, _24999_);
  nand _44420_ (_12261_, _12260_, _28096_);
  not _44421_ (_12262_, _12260_);
  nand _44422_ (_12263_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  nand _44423_ (_04816_, _12263_, _12261_);
  nor _44424_ (_12264_, _04172_, _01587_);
  nor _44425_ (_12265_, _12264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _44426_ (_12266_, _01630_, _01575_);
  nand _44427_ (_12267_, _12266_, _01614_);
  nand _44428_ (_12268_, _12267_, _07560_);
  nor _44429_ (_12269_, _12268_, _04172_);
  nor _44430_ (_12270_, _12269_, _12265_);
  nor _44431_ (_12271_, _12270_, _01573_);
  nand _44432_ (_12272_, _01573_, _24820_);
  nand _44433_ (_12273_, _12272_, _26487_);
  nor _44434_ (_04825_, _12273_, _12271_);
  nor _44435_ (_12274_, _25351_, _24862_);
  not _44436_ (_12275_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nand _44437_ (_12276_, _24862_, _12275_);
  nand _44438_ (_12277_, _12276_, _26487_);
  nor _44439_ (_28186_[7], _12277_, _12274_);
  nand _44440_ (_12278_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  nand _44441_ (_12279_, _24796_, _24789_);
  nand _44442_ (_04832_, _12279_, _12278_);
  nand _44443_ (_12280_, _03520_, _24830_);
  nand _44444_ (_12281_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nand _44445_ (_04838_, _12281_, _12280_);
  nor _44446_ (_12282_, _11782_, _25057_);
  nand _44447_ (_12283_, _12282_, _25203_);
  not _44448_ (_12284_, _12282_);
  nand _44449_ (_12285_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nand _44450_ (_04840_, _12285_, _12283_);
  nand _44451_ (_12286_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  nand _44452_ (_12287_, _08153_, _24927_);
  nand _44453_ (_04843_, _12287_, _12286_);
  nand _44454_ (_12288_, _12089_, _25039_);
  nand _44455_ (_12289_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  nand _44456_ (_04846_, _12289_, _12288_);
  nand _44457_ (_12290_, _12089_, _25203_);
  nand _44458_ (_12291_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nand _44459_ (_04857_, _12291_, _12290_);
  nand _44460_ (_12292_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  nand _44461_ (_12293_, _08153_, _25039_);
  nand _44462_ (_04859_, _12293_, _12292_);
  nor _44463_ (_12294_, _11782_, _28080_);
  nand _44464_ (_12295_, _12294_, _24927_);
  not _44465_ (_12296_, _12294_);
  nand _44466_ (_12297_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  nand _44467_ (_04863_, _12297_, _12295_);
  nand _44468_ (_12298_, _00115_, _24789_);
  nand _44469_ (_12299_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  nand _44470_ (_04866_, _12299_, _12298_);
  nand _44471_ (_12300_, _12294_, _25203_);
  nand _44472_ (_12301_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  nand _44473_ (_04869_, _12301_, _12300_);
  nand _44474_ (_12302_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  nand _44475_ (_12303_, _08153_, _25203_);
  nand _44476_ (_04890_, _12303_, _12302_);
  nor _44477_ (_12304_, _11782_, _28073_);
  nand _44478_ (_12305_, _12304_, _24830_);
  not _44479_ (_12306_, _12304_);
  nand _44480_ (_12307_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  nand _44481_ (_04896_, _12307_, _12305_);
  nand _44482_ (_12308_, _12089_, _24789_);
  nand _44483_ (_12309_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  nand _44484_ (_04918_, _12309_, _12308_);
  nand _44485_ (_12310_, _04308_, _25203_);
  nand _44486_ (_12311_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nand _44487_ (_04921_, _12311_, _12310_);
  nor _44488_ (_12312_, _11782_, _00122_);
  nand _44489_ (_12313_, _12312_, _24789_);
  not _44490_ (_12314_, _12312_);
  nand _44491_ (_12315_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  nand _44492_ (_04925_, _12315_, _12313_);
  nand _44493_ (_12316_, _12312_, _25203_);
  nand _44494_ (_12317_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  nand _44495_ (_04935_, _12317_, _12316_);
  nand _44496_ (_12318_, _12089_, _25150_);
  nand _44497_ (_12319_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nand _44498_ (_04938_, _12319_, _12318_);
  nand _44499_ (_12320_, _12089_, _24927_);
  nand _44500_ (_12321_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  nand _44501_ (_04943_, _12321_, _12320_);
  nand _44502_ (_12322_, _08354_, _25039_);
  nand _44503_ (_12323_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nand _44504_ (_04946_, _12323_, _12322_);
  nor _44505_ (_12324_, _11782_, _25047_);
  nand _44506_ (_12325_, _12324_, _25203_);
  not _44507_ (_12326_, _12324_);
  nand _44508_ (_12327_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nand _44509_ (_04951_, _12327_, _12325_);
  nand _44510_ (_12328_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  nand _44511_ (_12329_, _08153_, _24789_);
  nand _44512_ (_04956_, _12329_, _12328_);
  nor _44513_ (_12330_, _11782_, _00415_);
  nand _44514_ (_12331_, _12330_, _24789_);
  not _44515_ (_12332_, _12330_);
  nand _44516_ (_12333_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  nand _44517_ (_04963_, _12333_, _12331_);
  nand _44518_ (_12334_, _12330_, _25039_);
  nand _44519_ (_12335_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  nand _44520_ (_04966_, _12335_, _12334_);
  nand _44521_ (_12336_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nand _44522_ (_12337_, _08153_, _25150_);
  nand _44523_ (_04970_, _12337_, _12336_);
  nor _44524_ (_12338_, _11782_, _00393_);
  nand _44525_ (_12339_, _12338_, _24789_);
  not _44526_ (_12340_, _12338_);
  nand _44527_ (_12341_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  nand _44528_ (_04975_, _12341_, _12339_);
  nand _44529_ (_12342_, _12235_, _24789_);
  nand _44530_ (_12343_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  nand _44531_ (_04981_, _12343_, _12342_);
  nand _44532_ (_12344_, _01178_, _28096_);
  nand _44533_ (_12345_, _01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand _44534_ (_04983_, _12345_, _12344_);
  nand _44535_ (_12346_, _12235_, _25150_);
  nand _44536_ (_12347_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  nand _44537_ (_04987_, _12347_, _12346_);
  nor _44538_ (_12348_, _11782_, _24882_);
  nand _44539_ (_12349_, _12348_, _24789_);
  not _44540_ (_12350_, _12348_);
  nand _44541_ (_12351_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  nand _44542_ (_04993_, _12351_, _12349_);
  nand _44543_ (_12352_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nand _44544_ (_12353_, _08158_, _25203_);
  nand _44545_ (_04997_, _12353_, _12352_);
  nand _44546_ (_12354_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  nand _44547_ (_12355_, _08158_, _24927_);
  nand _44548_ (_05016_, _12355_, _12354_);
  nand _44549_ (_12356_, _12348_, _28096_);
  nand _44550_ (_12357_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  nand _44551_ (_05018_, _12357_, _12356_);
  nand _44552_ (_12358_, _12348_, _24830_);
  nand _44553_ (_12359_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nand _44554_ (_05024_, _12359_, _12358_);
  nand _44555_ (_12360_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nand _44556_ (_12361_, _08158_, _25039_);
  nand _44557_ (_05028_, _12361_, _12360_);
  nor _44558_ (_12362_, _11782_, _00629_);
  nand _44559_ (_12363_, _12362_, _24789_);
  not _44560_ (_12365_, _12362_);
  nand _44561_ (_12366_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  nand _44562_ (_05033_, _12366_, _12363_);
  nand _44563_ (_12367_, _11862_, _28096_);
  nand _44564_ (_12368_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nand _44565_ (_05040_, _12368_, _12367_);
  nand _44566_ (_12369_, _12362_, _25099_);
  nand _44567_ (_12370_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nand _44568_ (_05042_, _12370_, _12369_);
  nand _44569_ (_12371_, _12330_, _25099_);
  nand _44570_ (_12372_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  nand _44571_ (_05045_, _12372_, _12371_);
  nor _44572_ (_12373_, _11782_, _00954_);
  nand _44573_ (_12374_, _12373_, _25150_);
  not _44574_ (_12375_, _12373_);
  nand _44575_ (_12376_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  nand _44576_ (_05054_, _12376_, _12374_);
  nand _44577_ (_12377_, _11862_, _25099_);
  nand _44578_ (_12378_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  nand _44579_ (_05057_, _12378_, _12377_);
  nand _44580_ (_12379_, _12373_, _25203_);
  nand _44581_ (_12380_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  nand _44582_ (_05068_, _12380_, _12379_);
  nand _44583_ (_12381_, _12282_, _24927_);
  nand _44584_ (_12382_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  nand _44585_ (_05078_, _12382_, _12381_);
  nand _44586_ (_12383_, _12294_, _24789_);
  nand _44587_ (_12384_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  nand _44588_ (_05086_, _12384_, _12383_);
  nand _44589_ (_12385_, _12294_, _24830_);
  nand _44590_ (_12386_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nand _44591_ (_05096_, _12386_, _12385_);
  nand _44592_ (_12387_, _11862_, _25203_);
  nand _44593_ (_12388_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  nand _44594_ (_05099_, _12388_, _12387_);
  nand _44595_ (_12389_, _08154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nand _44596_ (_12390_, _08153_, _24830_);
  nand _44597_ (_05105_, _12390_, _12389_);
  nand _44598_ (_12391_, _12304_, _24927_);
  nand _44599_ (_12392_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  nand _44600_ (_05107_, _12392_, _12391_);
  nand _44601_ (_12393_, _12304_, _28096_);
  nand _44602_ (_12394_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nand _44603_ (_05110_, _12394_, _12393_);
  nand _44604_ (_12395_, _12312_, _24830_);
  nand _44605_ (_12396_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nand _44606_ (_05142_, _12396_, _12395_);
  nand _44607_ (_12397_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  nand _44608_ (_12398_, _08158_, _24789_);
  nand _44609_ (_05144_, _12398_, _12397_);
  nor _44610_ (_05147_, _01577_, rst);
  nand _44611_ (_12399_, _12324_, _24927_);
  nand _44612_ (_12400_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  nand _44613_ (_05150_, _12400_, _12399_);
  nor _44614_ (_12401_, _07818_, _28080_);
  nand _44615_ (_12402_, _12401_, _25039_);
  not _44616_ (_12403_, _12401_);
  nand _44617_ (_12404_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  nand _44618_ (_05154_, _12404_, _12402_);
  nand _44619_ (_12405_, _12401_, _25203_);
  nand _44620_ (_12406_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  nand _44621_ (_05163_, _12406_, _12405_);
  nand _44622_ (_12407_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  nand _44623_ (_12408_, _08158_, _25150_);
  nand _44624_ (_05165_, _12408_, _12407_);
  nand _44625_ (_12409_, _12338_, _28096_);
  nand _44626_ (_12410_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  nand _44627_ (_05168_, _12410_, _12409_);
  nand _44628_ (_12411_, _12362_, _25203_);
  nand _44629_ (_12412_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  nand _44630_ (_05200_, _12412_, _12411_);
  nor _44631_ (_12413_, _07818_, _00926_);
  nand _44632_ (_12414_, _12413_, _24830_);
  not _44633_ (_12415_, _12413_);
  nand _44634_ (_12416_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nand _44635_ (_05224_, _12416_, _12414_);
  not _44636_ (_12417_, _00305_);
  nor _44637_ (_12418_, _12417_, _00170_);
  nor _44638_ (_12419_, _00170_, _00184_);
  nor _44639_ (_12420_, _12419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor _44640_ (_12421_, _12420_, _12418_);
  nand _44641_ (_12422_, _00205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nor _44642_ (_12423_, _12422_, _00244_);
  nor _44643_ (_12424_, _12423_, _12421_);
  nor _44644_ (_12425_, _12424_, _00157_);
  not _44645_ (_12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nor _44646_ (_12427_, _00158_, _12426_);
  nor _44647_ (_12428_, _12427_, _12425_);
  nor _44648_ (_12429_, _12428_, _00150_);
  nor _44649_ (_12430_, _00302_, _25088_);
  nor _44650_ (_12431_, _12430_, _12429_);
  nor _44651_ (_12432_, _12431_, _00140_);
  nor _44652_ (_12433_, _00141_, _00176_);
  nor _44653_ (_12434_, _12433_, _12432_);
  nor _44654_ (_05251_, _12434_, rst);
  nor _44655_ (_12435_, _00302_, _25703_);
  nor _44656_ (_12436_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand _44657_ (_12437_, _12418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  not _44658_ (_12438_, _12418_);
  nand _44659_ (_12439_, _12438_, _00180_);
  nand _44660_ (_12440_, _12439_, _12437_);
  nand _44661_ (_12441_, _12440_, _00158_);
  nand _44662_ (_12442_, _00205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor _44663_ (_12443_, _12442_, _00244_);
  nor _44664_ (_12444_, _12443_, _12441_);
  nor _44665_ (_12445_, _12444_, _12436_);
  nand _44666_ (_12446_, _12445_, _00240_);
  nand _44667_ (_12447_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand _44668_ (_12448_, _12447_, _12446_);
  nor _44669_ (_12449_, _12448_, _12435_);
  nor _44670_ (_05254_, _12449_, rst);
  nand _44671_ (_12450_, _12312_, _25039_);
  nand _44672_ (_12451_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  nand _44673_ (_05256_, _12451_, _12450_);
  nor _44674_ (_12452_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _44675_ (_12453_, _12452_, _12419_);
  nor _44676_ (_12454_, _12453_, _00157_);
  nor _44677_ (_12455_, _00204_, _05904_);
  nand _44678_ (_12456_, _12455_, _00245_);
  nand _44679_ (_12457_, _12456_, _12454_);
  nand _44680_ (_12458_, _00157_, _05904_);
  nand _44681_ (_12459_, _12458_, _12457_);
  nor _44682_ (_12460_, _12459_, _00241_);
  nand _44683_ (_12461_, _00150_, _24821_);
  nand _44684_ (_12462_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _44685_ (_12463_, _12462_, _12461_);
  nor _44686_ (_12464_, _12463_, _12460_);
  nor _44687_ (_05262_, _12464_, rst);
  nor _44688_ (_12465_, _07818_, _24795_);
  nand _44689_ (_12466_, _12465_, _25099_);
  not _44690_ (_12467_, _12465_);
  nand _44691_ (_12468_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  nand _44692_ (_05265_, _12468_, _12466_);
  nand _44693_ (_12469_, _12465_, _25203_);
  nand _44694_ (_12470_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  nand _44695_ (_05268_, _12470_, _12469_);
  nand _44696_ (_12471_, _12465_, _24927_);
  nand _44697_ (_12472_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  nand _44698_ (_05272_, _12472_, _12471_);
  nand _44699_ (_12473_, _12465_, _25150_);
  nand _44700_ (_12474_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  nand _44701_ (_05280_, _12474_, _12473_);
  nand _44702_ (_12475_, _12348_, _25039_);
  nand _44703_ (_12476_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nand _44704_ (_05283_, _12476_, _12475_);
  nand _44705_ (_12477_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  nand _44706_ (_12478_, _08163_, _25150_);
  nand _44707_ (_05289_, _12478_, _12477_);
  nand _44708_ (_12479_, _07819_, _24927_);
  nand _44709_ (_12480_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  nand _44710_ (_05294_, _12480_, _12479_);
  nand _44711_ (_12481_, _07819_, _25150_);
  nand _44712_ (_12482_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  nand _44713_ (_05303_, _12482_, _12481_);
  nor _44714_ (_12483_, _07818_, _24999_);
  nand _44715_ (_12484_, _12483_, _24830_);
  not _44716_ (_12485_, _12483_);
  nand _44717_ (_12486_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  nand _44718_ (_05310_, _12486_, _12484_);
  nor _44719_ (_05312_, _26940_, rst);
  nor _44720_ (_05315_, _02586_, rst);
  nor _44721_ (_05317_, _27076_, rst);
  nand _44722_ (_12487_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  nand _44723_ (_12488_, _08163_, _24927_);
  nand _44724_ (_05321_, _12488_, _12487_);
  nor _44725_ (_05324_, _02710_, rst);
  nor _44726_ (_05326_, _02641_, rst);
  nand _44727_ (_12489_, _12483_, _25099_);
  nand _44728_ (_12490_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nand _44729_ (_05330_, _12490_, _12489_);
  nand _44730_ (_12492_, _12483_, _25039_);
  nand _44731_ (_12493_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  nand _44732_ (_05332_, _12493_, _12492_);
  nand _44733_ (_12494_, _12483_, _24927_);
  nand _44734_ (_12495_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  nand _44735_ (_05335_, _12495_, _12494_);
  nand _44736_ (_12496_, _12483_, _24789_);
  nand _44737_ (_12497_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  nand _44738_ (_05353_, _12497_, _12496_);
  nor _44739_ (_12498_, _07818_, _24978_);
  nand _44740_ (_12499_, _12498_, _24830_);
  not _44741_ (_12500_, _12498_);
  nand _44742_ (_12501_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nand _44743_ (_05358_, _12501_, _12499_);
  nand _44744_ (_12502_, _24768_, _26812_);
  nand _44745_ (_12503_, _12502_, _26487_);
  nor _44746_ (_05360_, _12503_, _12187_);
  nand _44747_ (_12504_, _12498_, _25203_);
  nand _44748_ (_12505_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nand _44749_ (_05363_, _12505_, _12504_);
  nand _44750_ (_12506_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  nand _44751_ (_12507_, _08163_, _25039_);
  nand _44752_ (_05366_, _12507_, _12506_);
  nand _44753_ (_12508_, _12498_, _25039_);
  nand _44754_ (_12509_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  nand _44755_ (_05369_, _12509_, _12508_);
  nand _44756_ (_12510_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  nand _44757_ (_12511_, _06807_, _24830_);
  nand _44758_ (_05373_, _12511_, _12510_);
  nand _44759_ (_12512_, _12498_, _25150_);
  nand _44760_ (_12513_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nand _44761_ (_05375_, _12513_, _12512_);
  nand _44762_ (_12514_, _12373_, _28096_);
  nand _44763_ (_12515_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nand _44764_ (_05377_, _12515_, _12514_);
  nor _44765_ (_05381_, _02445_, rst);
  nand _44766_ (_12516_, _12373_, _24830_);
  nand _44767_ (_12517_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  nand _44768_ (_05385_, _12517_, _12516_);
  not _44769_ (_12518_, _02061_);
  nor _44770_ (_05387_, _12518_, rst);
  not _44771_ (_12519_, _02007_);
  nor _44772_ (_05389_, _12519_, rst);
  nand _44773_ (_12520_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nand _44774_ (_12521_, _11607_, _25099_);
  nand _44775_ (_05391_, _12521_, _12520_);
  nor _44776_ (_05395_, _02194_, rst);
  nor _44777_ (_05397_, _02265_, rst);
  nor _44778_ (_12522_, _07818_, _24059_);
  nand _44779_ (_12523_, _12522_, _28096_);
  not _44780_ (_12524_, _12522_);
  nand _44781_ (_12525_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nand _44782_ (_05400_, _12525_, _12523_);
  nor _44783_ (_05402_, _02128_, rst);
  nand _44784_ (_12526_, _12373_, _25099_);
  nand _44785_ (_12527_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  nand _44786_ (_05409_, _12527_, _12526_);
  nor _44787_ (_05412_, _02336_, rst);
  nand _44788_ (_12528_, _11609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  nand _44789_ (_12529_, _11607_, _28096_);
  nand _44790_ (_05420_, _12529_, _12528_);
  nand _44791_ (_12530_, _12373_, _25039_);
  nand _44792_ (_12531_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nand _44793_ (_05422_, _12531_, _12530_);
  nand _44794_ (_12532_, _12522_, _25203_);
  nand _44795_ (_12533_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nand _44796_ (_05424_, _12533_, _12532_);
  nand _44797_ (_12534_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nand _44798_ (_12535_, _06807_, _25039_);
  nand _44799_ (_05429_, _12535_, _12534_);
  nand _44800_ (_12536_, _06808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nand _44801_ (_12537_, _06807_, _28096_);
  nand _44802_ (_05432_, _12537_, _12536_);
  nand _44803_ (_12538_, _12522_, _24927_);
  nand _44804_ (_12539_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  nand _44805_ (_05434_, _12539_, _12538_);
  nand _44806_ (_12540_, _12522_, _24789_);
  nand _44807_ (_12541_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  nand _44808_ (_05449_, _12541_, _12540_);
  nand _44809_ (_12542_, _12373_, _24927_);
  nand _44810_ (_12543_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  nand _44811_ (_05451_, _12543_, _12542_);
  nand _44812_ (_12544_, _12413_, _28096_);
  nand _44813_ (_12545_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nand _44814_ (_05458_, _12545_, _12544_);
  nand _44815_ (_12546_, _12373_, _24789_);
  nand _44816_ (_12547_, _12375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  nand _44817_ (_05471_, _12547_, _12546_);
  nand _44818_ (_12548_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  nand _44819_ (_12549_, _05864_, _28096_);
  nand _44820_ (_05474_, _12549_, _12548_);
  nand _44821_ (_12550_, _12413_, _25203_);
  nand _44822_ (_12551_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  nand _44823_ (_05477_, _12551_, _12550_);
  nand _44824_ (_12552_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  nand _44825_ (_12553_, _05864_, _25150_);
  nand _44826_ (_05483_, _12553_, _12552_);
  nand _44827_ (_12554_, _12330_, _24830_);
  nand _44828_ (_12555_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  nand _44829_ (_05485_, _12555_, _12554_);
  nand _44830_ (_12556_, _12413_, _24927_);
  nand _44831_ (_12557_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  nand _44832_ (_05490_, _12557_, _12556_);
  nand _44833_ (_12558_, _12413_, _24789_);
  nand _44834_ (_12559_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  nand _44835_ (_05491_, _12559_, _12558_);
  nand _44836_ (_12560_, _05865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  nand _44837_ (_12561_, _05864_, _24927_);
  nand _44838_ (_05494_, _12561_, _12560_);
  nand _44839_ (_12562_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nand _44840_ (_12563_, _08158_, _25099_);
  nand _44841_ (_05496_, _12563_, _12562_);
  nand _44842_ (_12564_, _12362_, _24830_);
  nand _44843_ (_12565_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  nand _44844_ (_05504_, _12565_, _12564_);
  nor _44845_ (_12566_, _03546_, _00114_);
  not _44846_ (_12567_, _12566_);
  nand _44847_ (_12568_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  nand _44848_ (_12569_, _12566_, _24830_);
  nand _44849_ (_05510_, _12569_, _12568_);
  nand _44850_ (_12570_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  nand _44851_ (_12571_, _12566_, _28096_);
  nand _44852_ (_05514_, _12571_, _12570_);
  nand _44853_ (_12572_, _12362_, _28096_);
  nand _44854_ (_12573_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  nand _44855_ (_05519_, _12573_, _12572_);
  nand _44856_ (_12574_, _12362_, _25039_);
  nand _44857_ (_12575_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  nand _44858_ (_05525_, _12575_, _12574_);
  nand _44859_ (_12576_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  nand _44860_ (_12577_, _12566_, _25039_);
  nand _44861_ (_05527_, _12577_, _12576_);
  nand _44862_ (_12578_, _08159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nand _44863_ (_12579_, _08158_, _24830_);
  nand _44864_ (_05529_, _12579_, _12578_);
  nand _44865_ (_12580_, _05736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  nand _44866_ (_12581_, _05735_, _24927_);
  nand _44867_ (_05532_, _12581_, _12580_);
  nand _44868_ (_12582_, _12362_, _24927_);
  nand _44869_ (_12583_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  nand _44870_ (_05543_, _12583_, _12582_);
  nand _44871_ (_12584_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  nand _44872_ (_12585_, _12566_, _24927_);
  nand _44873_ (_05545_, _12585_, _12584_);
  nand _44874_ (_12586_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  nand _44875_ (_12587_, _05685_, _24830_);
  nand _44876_ (_05549_, _12587_, _12586_);
  nand _44877_ (_12588_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  nand _44878_ (_12589_, _12566_, _24789_);
  nand _44879_ (_05569_, _12589_, _12588_);
  nor _44880_ (_12590_, _03546_, _00629_);
  not _44881_ (_12591_, _12590_);
  nand _44882_ (_12592_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nand _44883_ (_12593_, _12590_, _24830_);
  nand _44884_ (_05573_, _12593_, _12592_);
  nand _44885_ (_12594_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  nand _44886_ (_12595_, _12590_, _28096_);
  nand _44887_ (_05576_, _12595_, _12594_);
  nand _44888_ (_12596_, _05686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  nand _44889_ (_12597_, _05685_, _25150_);
  nand _44890_ (_05580_, _12597_, _12596_);
  nand _44891_ (_12598_, _12362_, _25150_);
  nand _44892_ (_12599_, _12365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  nand _44893_ (_05583_, _12599_, _12598_);
  nand _44894_ (_12600_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nand _44895_ (_12601_, _04322_, _28096_);
  nand _44896_ (_05591_, _12601_, _12600_);
  nand _44897_ (_12602_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nand _44898_ (_12603_, _12590_, _25203_);
  nand _44899_ (_05594_, _12603_, _12602_);
  nand _44900_ (_12604_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  nand _44901_ (_12605_, _12590_, _25150_);
  nand _44902_ (_05596_, _12605_, _12604_);
  nand _44903_ (_12606_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  nand _44904_ (_12607_, _08163_, _24789_);
  nand _44905_ (_05598_, _12607_, _12606_);
  nand _44906_ (_12608_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  nand _44907_ (_12609_, _04322_, _25150_);
  nand _44908_ (_05603_, _12609_, _12608_);
  nand _44909_ (_12610_, _12348_, _25099_);
  nand _44910_ (_12611_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  nand _44911_ (_05608_, _12611_, _12610_);
  nand _44912_ (_12612_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  nand _44913_ (_12613_, _12590_, _24789_);
  nand _44914_ (_05610_, _12613_, _12612_);
  nand _44915_ (_12614_, _04323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  nand _44916_ (_12615_, _04322_, _24927_);
  nand _44917_ (_05613_, _12615_, _12614_);
  nand _44918_ (_12616_, _12348_, _25203_);
  nand _44919_ (_12617_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  nand _44920_ (_05615_, _12617_, _12616_);
  nor _44921_ (_12618_, _03546_, _24882_);
  not _44922_ (_12619_, _12618_);
  nand _44923_ (_12620_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  nand _44924_ (_12621_, _12618_, _25099_);
  nand _44925_ (_05623_, _12621_, _12620_);
  nand _44926_ (_12622_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  nand _44927_ (_12623_, _04299_, _24830_);
  nand _44928_ (_05626_, _12623_, _12622_);
  nand _44929_ (_12624_, _12348_, _24927_);
  nand _44930_ (_12625_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  nand _44931_ (_05631_, _12625_, _12624_);
  nand _44932_ (_12626_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  nand _44933_ (_12627_, _12618_, _28096_);
  nand _44934_ (_05635_, _12627_, _12626_);
  nand _44935_ (_12628_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  nand _44936_ (_12629_, _04299_, _24789_);
  nand _44937_ (_05647_, _12629_, _12628_);
  nand _44938_ (_12630_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  nand _44939_ (_12631_, _12618_, _24927_);
  nand _44940_ (_05673_, _12631_, _12630_);
  nand _44941_ (_12632_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  nand _44942_ (_12633_, _12618_, _24789_);
  nand _44943_ (_05674_, _12633_, _12632_);
  nand _44944_ (_12634_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  nand _44945_ (_12635_, _04255_, _25203_);
  nand _44946_ (_05677_, _12635_, _12634_);
  nand _44947_ (_12636_, _12348_, _25150_);
  nand _44948_ (_12637_, _12350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nand _44949_ (_05681_, _12637_, _12636_);
  nand _44950_ (_12638_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nand _44951_ (_12639_, _04255_, _25099_);
  nand _44952_ (_05687_, _12639_, _12638_);
  nand _44953_ (_12640_, _12338_, _24830_);
  nand _44954_ (_12641_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nand _44955_ (_05689_, _12641_, _12640_);
  nor _44956_ (_12642_, _03546_, _00393_);
  not _44957_ (_12643_, _12642_);
  nand _44958_ (_12644_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nand _44959_ (_12645_, _12642_, _24830_);
  nand _44960_ (_05692_, _12645_, _12644_);
  nand _44961_ (_12646_, _04257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nand _44962_ (_12647_, _04255_, _25150_);
  nand _44963_ (_05694_, _12647_, _12646_);
  nand _44964_ (_12648_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  nand _44965_ (_12649_, _12642_, _28096_);
  nand _44966_ (_05696_, _12649_, _12648_);
  nand _44967_ (_12650_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  nand _44968_ (_12651_, _04166_, _25150_);
  nand _44969_ (_05703_, _12651_, _12650_);
  nand _44970_ (_12652_, _12338_, _25099_);
  nand _44971_ (_12653_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nand _44972_ (_05707_, _12653_, _12652_);
  nand _44973_ (_12654_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nand _44974_ (_12655_, _12642_, _25039_);
  nand _44975_ (_05710_, _12655_, _12654_);
  nand _44976_ (_12656_, _04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nand _44977_ (_12657_, _04166_, _25203_);
  nand _44978_ (_05713_, _12657_, _12656_);
  nand _44979_ (_12658_, _12338_, _25203_);
  nand _44980_ (_12660_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  nand _44981_ (_05714_, _12660_, _12658_);
  nand _44982_ (_12661_, _03886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nand _44983_ (_12662_, _03884_, _25039_);
  nand _44984_ (_05717_, _12662_, _12661_);
  nor _44985_ (_12663_, _00415_, _25159_);
  nand _44986_ (_12664_, _12663_, _24789_);
  not _44987_ (_12665_, _12663_);
  nand _44988_ (_12666_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand _44989_ (_05720_, _12666_, _12664_);
  nand _44990_ (_12667_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nand _44991_ (_12668_, _12642_, _25150_);
  nand _44992_ (_05723_, _12668_, _12667_);
  nand _44993_ (_12669_, _12338_, _25039_);
  nand _44994_ (_12670_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  nand _44995_ (_05728_, _12670_, _12669_);
  nor _44996_ (_12671_, _03546_, _00954_);
  not _44997_ (_12672_, _12671_);
  nand _44998_ (_12673_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  nand _44999_ (_12674_, _12671_, _25099_);
  nand _45000_ (_05732_, _12674_, _12673_);
  nand _45001_ (_12676_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  nand _45002_ (_12677_, _12671_, _25039_);
  nand _45003_ (_05752_, _12677_, _12676_);
  nand _45004_ (_12678_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nand _45005_ (_12679_, _10214_, _25150_);
  nand _45006_ (_05755_, _12679_, _12678_);
  nand _45007_ (_12680_, _10226_, _24789_);
  nand _45008_ (_12681_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand _45009_ (_05758_, _12681_, _12680_);
  nand _45010_ (_12682_, _04111_, _24830_);
  nand _45011_ (_12683_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand _45012_ (_05760_, _12683_, _12682_);
  nand _45013_ (_12684_, _12338_, _24927_);
  nand _45014_ (_12685_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  nand _45015_ (_05765_, _12685_, _12684_);
  nand _45016_ (_12686_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  nand _45017_ (_12687_, _12671_, _24927_);
  nand _45018_ (_05768_, _12687_, _12686_);
  nor _45019_ (_12688_, _25159_, _25047_);
  nand _45020_ (_12689_, _12688_, _25203_);
  not _45021_ (_12690_, _12688_);
  nand _45022_ (_12691_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nand _45023_ (_05773_, _12691_, _12689_);
  nand _45024_ (_12692_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  nand _45025_ (_12693_, _12671_, _24789_);
  nand _45026_ (_05776_, _12693_, _12692_);
  nand _45027_ (_12694_, _12688_, _28096_);
  nand _45028_ (_12695_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nand _45029_ (_05778_, _12695_, _12694_);
  nand _45030_ (_12696_, _12688_, _25099_);
  nand _45031_ (_12697_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand _45032_ (_05782_, _12697_, _12696_);
  nor _45033_ (_12698_, _03546_, _00415_);
  not _45034_ (_12699_, _12698_);
  nand _45035_ (_12700_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nand _45036_ (_12701_, _12698_, _24830_);
  nand _45037_ (_05787_, _12701_, _12700_);
  nand _45038_ (_12702_, _12338_, _25150_);
  nand _45039_ (_12703_, _12340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nand _45040_ (_05789_, _12703_, _12702_);
  nand _45041_ (_12704_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nand _45042_ (_12705_, _12698_, _25203_);
  nand _45043_ (_05793_, _12705_, _12704_);
  nand _45044_ (_12706_, _03548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  nand _45045_ (_12707_, _03547_, _28096_);
  nand _45046_ (_05796_, _12707_, _12706_);
  nand _45047_ (_12708_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  nand _45048_ (_12709_, _10214_, _24789_);
  nand _45049_ (_05804_, _12709_, _12708_);
  nor _45050_ (_12710_, _28057_, _25047_);
  nand _45051_ (_12711_, _12710_, _24789_);
  not _45052_ (_12712_, _12710_);
  nand _45053_ (_12713_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  nand _45054_ (_05807_, _12713_, _12711_);
  nand _45055_ (_12714_, _12330_, _28096_);
  nand _45056_ (_12715_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nand _45057_ (_05809_, _12715_, _12714_);
  nand _45058_ (_12716_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  nand _45059_ (_12717_, _12698_, _25039_);
  nand _45060_ (_05811_, _12717_, _12716_);
  nand _45061_ (_12719_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  nand _45062_ (_12720_, _12698_, _25150_);
  nand _45063_ (_05814_, _12720_, _12719_);
  nand _45064_ (_12721_, _12663_, _24830_);
  nand _45065_ (_12722_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand _45066_ (_05823_, _12722_, _12721_);
  nand _45067_ (_12723_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  nand _45068_ (_12724_, _12698_, _24789_);
  nand _45069_ (_05827_, _12724_, _12723_);
  nand _45070_ (_12725_, _01175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  nand _45071_ (_12726_, _01174_, _24830_);
  nand _45072_ (_05833_, _12726_, _12725_);
  nand _45073_ (_12727_, _12663_, _25099_);
  nand _45074_ (_12728_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand _45075_ (_05835_, _12728_, _12727_);
  nand _45076_ (_12729_, _12330_, _25203_);
  nand _45077_ (_12730_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  nand _45078_ (_05839_, _12730_, _12729_);
  nand _45079_ (_12731_, _12401_, _24789_);
  nand _45080_ (_12732_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  nand _45081_ (_05843_, _12732_, _12731_);
  nand _45082_ (_12733_, _01521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nand _45083_ (_12734_, _01520_, _25150_);
  nand _45084_ (_05846_, _12734_, _12733_);
  nand _45085_ (_12735_, _12330_, _24927_);
  nand _45086_ (_12736_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  nand _45087_ (_05860_, _12736_, _12735_);
  nand _45088_ (_12737_, _12401_, _25150_);
  nand _45089_ (_12738_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nand _45090_ (_05866_, _12738_, _12737_);
  nand _45091_ (_12739_, _12401_, _24927_);
  nand _45092_ (_12740_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  nand _45093_ (_05869_, _12740_, _12739_);
  nand _45094_ (_12741_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nand _45095_ (_12742_, _01129_, _28096_);
  nand _45096_ (_05878_, _12742_, _12741_);
  nand _45097_ (_12743_, _12330_, _25150_);
  nand _45098_ (_12744_, _12332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  nand _45099_ (_05882_, _12744_, _12743_);
  nand _45100_ (_12745_, _01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  nand _45101_ (_12746_, _01129_, _24830_);
  nand _45102_ (_05888_, _12746_, _12745_);
  nand _45103_ (_12747_, _12324_, _24830_);
  nand _45104_ (_12748_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  nand _45105_ (_05890_, _12748_, _12747_);
  nand _45106_ (_12749_, _12663_, _25203_);
  nand _45107_ (_12750_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand _45108_ (_05893_, _12750_, _12749_);
  nand _45109_ (_12751_, _12663_, _24927_);
  nand _45110_ (_12752_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nand _45111_ (_05897_, _12752_, _12751_);
  nand _45112_ (_12753_, _12663_, _25039_);
  nand _45113_ (_12754_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nand _45114_ (_05905_, _12754_, _12753_);
  nand _45115_ (_12755_, _12324_, _25099_);
  nand _45116_ (_12756_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nand _45117_ (_05913_, _12756_, _12755_);
  nand _45118_ (_12757_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  nand _45119_ (_12758_, _01085_, _24789_);
  nand _45120_ (_05916_, _12758_, _12757_);
  nand _45121_ (_12759_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  nand _45122_ (_12760_, _08163_, _24830_);
  nand _45123_ (_05918_, _12760_, _12759_);
  nand _45124_ (_12761_, _01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nand _45125_ (_12762_, _01085_, _25039_);
  nand _45126_ (_05923_, _12762_, _12761_);
  nor _45127_ (_12763_, _07818_, _28073_);
  nand _45128_ (_12764_, _12763_, _24789_);
  not _45129_ (_12765_, _12763_);
  nand _45130_ (_12766_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  nand _45131_ (_05930_, _12766_, _12764_);
  nand _45132_ (_12767_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  nand _45133_ (_12768_, _00933_, _24927_);
  nand _45134_ (_05936_, _12768_, _12767_);
  nand _45135_ (_12769_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  nand _45136_ (_12770_, _08163_, _28096_);
  nand _45137_ (_05938_, _12770_, _12769_);
  nand _45138_ (_12771_, _12763_, _25150_);
  nand _45139_ (_12772_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nand _45140_ (_05940_, _12772_, _12771_);
  nand _45141_ (_12773_, _12324_, _28096_);
  nand _45142_ (_12774_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  nand _45143_ (_05945_, _12774_, _12773_);
  nand _45144_ (_12775_, _00934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nand _45145_ (_12776_, _00933_, _25203_);
  nand _45146_ (_05948_, _12776_, _12775_);
  nand _45147_ (_12777_, _12324_, _25039_);
  nand _45148_ (_12778_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nand _45149_ (_05951_, _12778_, _12777_);
  nand _45150_ (_12779_, _04111_, _25039_);
  nand _45151_ (_12780_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nand _45152_ (_05954_, _12780_, _12779_);
  nand _45153_ (_12781_, _08164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  nand _45154_ (_12782_, _08163_, _25099_);
  nand _45155_ (_05957_, _12782_, _12781_);
  nand _45156_ (_12783_, _04111_, _25099_);
  nand _45157_ (_12784_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand _45158_ (_05960_, _12784_, _12783_);
  nand _45159_ (_12785_, _00844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  nand _45160_ (_12786_, _00843_, _25203_);
  nand _45161_ (_05976_, _12786_, _12785_);
  nand _45162_ (_12787_, _04111_, _25203_);
  nand _45163_ (_12788_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nand _45164_ (_05978_, _12788_, _12787_);
  nand _45165_ (_12789_, _12324_, _25150_);
  nand _45166_ (_12790_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  nand _45167_ (_05993_, _12790_, _12789_);
  nand _45168_ (_12791_, _04111_, _24927_);
  nand _45169_ (_12792_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nand _45170_ (_05995_, _12792_, _12791_);
  nor _45171_ (_28182_[7], _27729_, rst);
  nand _45172_ (_12793_, _04111_, _24789_);
  nand _45173_ (_12794_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand _45174_ (_06004_, _12794_, _12793_);
  nand _45175_ (_12795_, _03858_, _25039_);
  nand _45176_ (_12796_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nand _45177_ (_06008_, _12796_, _12795_);
  nand _45178_ (_12797_, _12324_, _24789_);
  nand _45179_ (_12798_, _12326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  nand _45180_ (_06014_, _12798_, _12797_);
  nand _45181_ (_12799_, _00637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  nand _45182_ (_12800_, _00636_, _25150_);
  nand _45183_ (_06019_, _12800_, _12799_);
  nand _45184_ (_12801_, _12312_, _25099_);
  nand _45185_ (_12802_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  nand _45186_ (_06021_, _12802_, _12801_);
  nand _45187_ (_12803_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  nand _45188_ (_12804_, _00360_, _25099_);
  nand _45189_ (_06023_, _12804_, _12803_);
  nand _45190_ (_12805_, _00409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  nand _45191_ (_12806_, _00408_, _25150_);
  nand _45192_ (_06028_, _12806_, _12805_);
  nor _45193_ (_12807_, _00122_, _25159_);
  nand _45194_ (_12808_, _12807_, _24789_);
  not _45195_ (_12809_, _12807_);
  nand _45196_ (_12810_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nand _45197_ (_06034_, _12810_, _12808_);
  nand _45198_ (_12811_, _12312_, _28096_);
  nand _45199_ (_12812_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  nand _45200_ (_06041_, _12812_, _12811_);
  nand _45201_ (_12813_, _00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  nand _45202_ (_12814_, _00360_, _24927_);
  nand _45203_ (_06043_, _12814_, _12813_);
  nand _45204_ (_12815_, _12401_, _25099_);
  nand _45205_ (_12816_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nand _45206_ (_06046_, _12816_, _12815_);
  nand _45207_ (_12817_, _12312_, _24927_);
  nand _45208_ (_12818_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  nand _45209_ (_06063_, _12818_, _12817_);
  nand _45210_ (_12819_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  nand _45211_ (_12820_, _24830_, _24074_);
  nand _45212_ (_06066_, _12820_, _12819_);
  nand _45213_ (_12821_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  nand _45214_ (_12822_, _08492_, _24789_);
  nand _45215_ (_06069_, _12822_, _12821_);
  nand _45216_ (_12823_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  nand _45217_ (_12824_, _10214_, _25099_);
  nand _45218_ (_06071_, _12824_, _12823_);
  nand _45219_ (_12825_, _12401_, _24830_);
  nand _45220_ (_12826_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nand _45221_ (_06073_, _12826_, _12825_);
  nand _45222_ (_12827_, _00331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  nand _45223_ (_12828_, _00330_, _24927_);
  nand _45224_ (_06075_, _12828_, _12827_);
  nand _45225_ (_12829_, _10226_, _28096_);
  nand _45226_ (_12830_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand _45227_ (_06079_, _12830_, _12829_);
  nand _45228_ (_12831_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  nand _45229_ (_12832_, _24927_, _24074_);
  nand _45230_ (_06081_, _12832_, _12831_);
  nand _45231_ (_12833_, _12312_, _25150_);
  nand _45232_ (_12834_, _12314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nand _45233_ (_06083_, _12834_, _12833_);
  nand _45234_ (_12835_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nand _45235_ (_12836_, _10214_, _24830_);
  nand _45236_ (_06085_, _12836_, _12835_);
  nand _45237_ (_12837_, _10226_, _25099_);
  nand _45238_ (_12838_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nand _45239_ (_06091_, _12838_, _12837_);
  nand _45240_ (_12839_, _11937_, _28096_);
  nand _45241_ (_12840_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nand _45242_ (_06094_, _12840_, _12839_);
  nand _45243_ (_12841_, _24075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  nand _45244_ (_12842_, _25203_, _24074_);
  nand _45245_ (_06097_, _12842_, _12841_);
  nand _45246_ (_12843_, _10226_, _24830_);
  nand _45247_ (_12844_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nand _45248_ (_06099_, _12844_, _12843_);
  nand _45249_ (_12845_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  nand _45250_ (_12846_, _28096_, _24796_);
  nand _45251_ (_06105_, _12846_, _12845_);
  nand _45252_ (_12847_, _12763_, _25099_);
  nand _45253_ (_12848_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nand _45254_ (_06112_, _12848_, _12847_);
  nand _45255_ (_12849_, _12304_, _25099_);
  nand _45256_ (_12850_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nand _45257_ (_06118_, _12850_, _12849_);
  nand _45258_ (_12851_, _12763_, _24830_);
  nand _45259_ (_12852_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nand _45260_ (_06120_, _12852_, _12851_);
  nand _45261_ (_12853_, _12807_, _28096_);
  nand _45262_ (_12854_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nand _45263_ (_06123_, _12854_, _12853_);
  nand _45264_ (_12855_, _12807_, _25099_);
  nand _45265_ (_12856_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nand _45266_ (_06129_, _12856_, _12855_);
  nor _45267_ (_12857_, _07818_, _00122_);
  nand _45268_ (_12858_, _12857_, _24789_);
  not _45269_ (_12859_, _12857_);
  nand _45270_ (_12860_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  nand _45271_ (_06134_, _12860_, _12858_);
  nand _45272_ (_12861_, _12807_, _24830_);
  nand _45273_ (_12862_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nand _45274_ (_06137_, _12862_, _12861_);
  nand _45275_ (_12863_, _12304_, _25203_);
  nand _45276_ (_12864_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nand _45277_ (_06140_, _12864_, _12863_);
  nand _45278_ (_12865_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  nand _45279_ (_12866_, _10214_, _28096_);
  nand _45280_ (_06151_, _12866_, _12865_);
  nand _45281_ (_12868_, _12304_, _25039_);
  nand _45282_ (_12869_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nand _45283_ (_06156_, _12869_, _12868_);
  nand _45284_ (_12870_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nand _45285_ (_12871_, _10214_, _25039_);
  nand _45286_ (_06158_, _12871_, _12870_);
  nand _45287_ (_12872_, _12763_, _25039_);
  nand _45288_ (_12873_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nand _45289_ (_06165_, _12873_, _12872_);
  nand _45290_ (_12874_, _00115_, _25099_);
  nand _45291_ (_12875_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  nand _45292_ (_06168_, _12875_, _12874_);
  nand _45293_ (_12876_, _12807_, _24927_);
  nand _45294_ (_12877_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand _45295_ (_06170_, _12877_, _12876_);
  nand _45296_ (_12878_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  nand _45297_ (_12879_, _10214_, _25203_);
  nand _45298_ (_06174_, _12879_, _12878_);
  nand _45299_ (_12880_, _12807_, _25039_);
  nand _45300_ (_12881_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand _45301_ (_06181_, _12881_, _12880_);
  nand _45302_ (_12882_, _12807_, _25203_);
  nand _45303_ (_12883_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nand _45304_ (_06198_, _12883_, _12882_);
  nand _45305_ (_12884_, _12304_, _25150_);
  nand _45306_ (_12885_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  nand _45307_ (_06200_, _12885_, _12884_);
  nand _45308_ (_12886_, _00979_, _25099_);
  nand _45309_ (_12887_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  nand _45310_ (_06206_, _12887_, _12886_);
  nand _45311_ (_12888_, _12763_, _25203_);
  nand _45312_ (_12889_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nand _45313_ (_06211_, _12889_, _12888_);
  nand _45314_ (_12890_, _12304_, _24789_);
  nand _45315_ (_12891_, _12306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  nand _45316_ (_06214_, _12891_, _12890_);
  nand _45317_ (_12892_, _12294_, _25099_);
  nand _45318_ (_12893_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  nand _45319_ (_06219_, _12893_, _12892_);
  nand _45320_ (_12894_, _25166_, _24789_);
  nand _45321_ (_12895_, _25168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  nand _45322_ (_06227_, _12895_, _12894_);
  nand _45323_ (_12896_, _12688_, _24789_);
  nand _45324_ (_12897_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nand _45325_ (_06232_, _12897_, _12896_);
  nand _45326_ (_12898_, _12688_, _25150_);
  nand _45327_ (_12899_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nand _45328_ (_06240_, _12899_, _12898_);
  nand _45329_ (_12900_, _12294_, _28096_);
  nand _45330_ (_12901_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nand _45331_ (_06244_, _12901_, _12900_);
  nand _45332_ (_12902_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  nand _45333_ (_12903_, _08343_, _24789_);
  nand _45334_ (_06250_, _12903_, _12902_);
  nand _45335_ (_12904_, _25203_, _25152_);
  nand _45336_ (_12905_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  nand _45337_ (_06262_, _12905_, _12904_);
  nand _45338_ (_12906_, _12294_, _25039_);
  nand _45339_ (_12907_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  nand _45340_ (_06265_, _12907_, _12906_);
  nand _45341_ (_12908_, _12857_, _25203_);
  nand _45342_ (_12909_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  nand _45343_ (_06267_, _12909_, _12908_);
  nor _45344_ (_12910_, _00393_, _25159_);
  nand _45345_ (_12911_, _12910_, _24927_);
  not _45346_ (_12912_, _12910_);
  nand _45347_ (_12913_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand _45348_ (_06270_, _12913_, _12911_);
  nand _45349_ (_12914_, _06826_, _24830_);
  nand _45350_ (_12915_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nand _45351_ (_06275_, _12915_, _12914_);
  nand _45352_ (_12916_, _12910_, _25039_);
  nand _45353_ (_12917_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand _45354_ (_06278_, _12917_, _12916_);
  nand _45355_ (_12918_, _12294_, _25150_);
  nand _45356_ (_12919_, _12296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  nand _45357_ (_06284_, _12919_, _12918_);
  nand _45358_ (_12920_, _12857_, _28096_);
  nand _45359_ (_12921_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  nand _45360_ (_06286_, _12921_, _12920_);
  nand _45361_ (_12922_, _12910_, _25203_);
  nand _45362_ (_12923_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nand _45363_ (_06288_, _12923_, _12922_);
  nand _45364_ (_12924_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nand _45365_ (_12925_, _08492_, _25099_);
  nand _45366_ (_06298_, _12925_, _12924_);
  nand _45367_ (_12926_, _12282_, _24830_);
  nand _45368_ (_12927_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  nand _45369_ (_06302_, _12927_, _12926_);
  nand _45370_ (_12928_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  nand _45371_ (_12929_, _08492_, _24830_);
  nand _45372_ (_06326_, _12929_, _12928_);
  nand _45373_ (_12930_, _12104_, _24789_);
  nand _45374_ (_12931_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  nand _45375_ (_06330_, _12931_, _12930_);
  nand _45376_ (_12932_, _12282_, _25099_);
  nand _45377_ (_12933_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nand _45378_ (_06343_, _12933_, _12932_);
  nand _45379_ (_12934_, _12910_, _24789_);
  nand _45380_ (_12935_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nand _45381_ (_06354_, _12935_, _12934_);
  nand _45382_ (_12936_, _12910_, _25150_);
  nand _45383_ (_12937_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand _45384_ (_06363_, _12937_, _12936_);
  nand _45385_ (_12938_, _12282_, _28096_);
  nand _45386_ (_12939_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  nand _45387_ (_06365_, _12939_, _12938_);
  nand _45388_ (_12940_, _12282_, _25039_);
  nand _45389_ (_12941_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  nand _45390_ (_06374_, _12941_, _12940_);
  nand _45391_ (_12942_, _03911_, _25203_);
  nand _45392_ (_12943_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nand _45393_ (_06380_, _12943_, _12942_);
  nand _45394_ (_12944_, _12857_, _25150_);
  nand _45395_ (_12945_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  nand _45396_ (_06389_, _12945_, _12944_);
  nand _45397_ (_12946_, _25053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  nand _45398_ (_12947_, _25052_, _24927_);
  nand _45399_ (_06391_, _12947_, _12946_);
  nand _45400_ (_12948_, _00955_, _25099_);
  nand _45401_ (_12949_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  nand _45402_ (_06394_, _12949_, _12948_);
  nand _45403_ (_12950_, _12282_, _25150_);
  nand _45404_ (_12951_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  nand _45405_ (_06396_, _12951_, _12950_);
  nand _45406_ (_12952_, _03850_, _25099_);
  nand _45407_ (_12953_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  nand _45408_ (_06399_, _12953_, _12952_);
  nand _45409_ (_12954_, _12857_, _24927_);
  nand _45410_ (_12955_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  nand _45411_ (_06401_, _12955_, _12954_);
  nand _45412_ (_12956_, _12857_, _25039_);
  nand _45413_ (_12957_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  nand _45414_ (_06403_, _12957_, _12956_);
  nand _45415_ (_12958_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  nand _45416_ (_12959_, _04015_, _24830_);
  nand _45417_ (_06408_, _12959_, _12958_);
  nand _45418_ (_12960_, _03911_, _24789_);
  nand _45419_ (_12961_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  nand _45420_ (_06410_, _12961_, _12960_);
  nand _45421_ (_12962_, _01905_, _24789_);
  nand _45422_ (_12963_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nand _45423_ (_06413_, _12963_, _12962_);
  nand _45424_ (_12964_, _12282_, _24789_);
  nand _45425_ (_12965_, _12284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  nand _45426_ (_06415_, _12965_, _12964_);
  nand _45427_ (_12966_, _12260_, _24830_);
  nand _45428_ (_12967_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  nand _45429_ (_06421_, _12967_, _12966_);
  nand _45430_ (_12968_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  nand _45431_ (_12969_, _08492_, _25039_);
  nand _45432_ (_06423_, _12969_, _12968_);
  nand _45433_ (_12970_, _08387_, _25039_);
  nand _45434_ (_12971_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nand _45435_ (_06424_, _12971_, _12970_);
  nand _45436_ (_12972_, _08494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nand _45437_ (_12973_, _08492_, _25203_);
  nand _45438_ (_06444_, _12973_, _12972_);
  nand _45439_ (_12974_, _12260_, _25099_);
  nand _45440_ (_12975_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nand _45441_ (_06448_, _12975_, _12974_);
  nor _45442_ (_12976_, _07818_, _25047_);
  nand _45443_ (_12977_, _12976_, _25039_);
  not _45444_ (_12978_, _12976_);
  nand _45445_ (_12979_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  nand _45446_ (_06453_, _12979_, _12977_);
  nand _45447_ (_12980_, _08387_, _24789_);
  nand _45448_ (_12981_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  nand _45449_ (_06455_, _12981_, _12980_);
  nand _45450_ (_12982_, _12910_, _25099_);
  nand _45451_ (_12983_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nand _45452_ (_06467_, _12983_, _12982_);
  nand _45453_ (_12984_, _12976_, _25150_);
  nand _45454_ (_12985_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nand _45455_ (_06469_, _12985_, _12984_);
  nand _45456_ (_12986_, _12910_, _24830_);
  nand _45457_ (_12987_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nand _45458_ (_06471_, _12987_, _12986_);
  nand _45459_ (_12988_, _12976_, _24927_);
  nand _45460_ (_12989_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  nand _45461_ (_06474_, _12989_, _12988_);
  nor _45462_ (_12990_, _00591_, _00588_);
  not _45463_ (_12991_, _00601_);
  nand _45464_ (_12992_, _12991_, _00591_);
  nand _45465_ (_12993_, _12992_, _00538_);
  nor _45466_ (_12994_, _12993_, _12990_);
  nor _45467_ (_12995_, _12994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _45468_ (_12996_, _00609_);
  nand _45469_ (_12997_, _00668_, _12996_);
  nand _45470_ (_12998_, _00590_, _00570_);
  nand _45471_ (_12999_, _12998_, _12997_);
  nand _45472_ (_13000_, _12999_, _00538_);
  nand _45473_ (_13001_, _13000_, _26487_);
  nor _45474_ (_06487_, _13001_, _12995_);
  not _45475_ (_13002_, _11818_);
  nor _45476_ (_06502_, _13002_, rst);
  nand _45477_ (_13003_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nand _45478_ (_13004_, _08167_, _25203_);
  nand _45479_ (_06508_, _13004_, _13003_);
  nand _45480_ (_13005_, _11533_, _28096_);
  nand _45481_ (_13006_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand _45482_ (_06510_, _13006_, _13005_);
  not _45483_ (_13007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nor _45484_ (_13008_, _01383_, _13007_);
  nor _45485_ (_13009_, _01384_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nor _45486_ (_13010_, _13009_, _13008_);
  nor _45487_ (_06512_, _13010_, _01377_);
  nand _45488_ (_13011_, _01454_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _45489_ (_13012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _45490_ (_13013_, _13012_, _03739_);
  not _45491_ (_13014_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  not _45492_ (_13015_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _45493_ (_13016_, _13015_, _13014_);
  nand _45494_ (_13017_, _13016_, _01461_);
  nand _45495_ (_13018_, _13017_, _01503_);
  nand _45496_ (_13019_, _13018_, _13013_);
  nand _45497_ (_13020_, _13019_, _13011_);
  nor _45498_ (_13021_, _01503_, rxd_i);
  nor _45499_ (_13022_, _13021_, _01460_);
  nand _45500_ (_13023_, _13022_, _13020_);
  nand _45501_ (_13024_, _01410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _45502_ (_06514_, _13024_, _13023_);
  nand _45503_ (_13025_, _11533_, _25099_);
  nand _45504_ (_13026_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nand _45505_ (_06527_, _13026_, _13025_);
  nand _45506_ (_13027_, _12857_, _24830_);
  nand _45507_ (_13028_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  nand _45508_ (_06529_, _13028_, _13027_);
  nand _45509_ (_13029_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  nand _45510_ (_13030_, _08167_, _28096_);
  nand _45511_ (_06531_, _13030_, _13029_);
  nand _45512_ (_13031_, _00955_, _28096_);
  nand _45513_ (_13032_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  nand _45514_ (_06549_, _13032_, _13031_);
  nand _45515_ (_13033_, _12976_, _24789_);
  nand _45516_ (_13034_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nand _45517_ (_06552_, _13034_, _13033_);
  nor _45518_ (_06561_, _03971_, rst);
  nand _45519_ (_13035_, _11533_, _24927_);
  nand _45520_ (_13036_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand _45521_ (_06563_, _13036_, _13035_);
  nand _45522_ (_13037_, _11533_, _25039_);
  nand _45523_ (_13038_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand _45524_ (_06572_, _13038_, _13037_);
  nor _45525_ (_13039_, _26256_, _26241_);
  not _45526_ (_13040_, _13039_);
  nor _45527_ (_13041_, _13040_, _25723_);
  not _45528_ (_13042_, _13041_);
  nor _45529_ (_13043_, _13042_, _02415_);
  not _45530_ (_13044_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _45531_ (_13045_, _13042_, _13044_);
  nand _45532_ (_13046_, _13045_, _25630_);
  nor _45533_ (_13047_, _13046_, _13043_);
  nand _45534_ (_13048_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor _45535_ (_13049_, _13040_, _00227_);
  nand _45536_ (_13050_, _13049_, _24717_);
  nor _45537_ (_13051_, _13049_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor _45538_ (_13052_, _13051_, _26245_);
  nand _45539_ (_13053_, _13052_, _13050_);
  nand _45540_ (_13054_, _13053_, _13048_);
  nor _45541_ (_13055_, _13054_, _13047_);
  nor _45542_ (_06574_, _13055_, rst);
  nor _45543_ (_13056_, _07818_, _00415_);
  nand _45544_ (_13057_, _13056_, _25150_);
  not _45545_ (_13058_, _13056_);
  nand _45546_ (_13059_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  nand _45547_ (_06578_, _13059_, _13057_);
  nand _45548_ (_13060_, _13056_, _24789_);
  nand _45549_ (_13061_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  nand _45550_ (_06583_, _13061_, _13060_);
  nand _45551_ (_13062_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nand _45552_ (_13063_, _08167_, _25150_);
  nand _45553_ (_06591_, _13063_, _13062_);
  nand _45554_ (_13064_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  nand _45555_ (_13065_, _08167_, _24927_);
  nand _45556_ (_06595_, _13065_, _13064_);
  nand _45557_ (_13066_, _12976_, _28096_);
  nand _45558_ (_13067_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  nand _45559_ (_06602_, _13067_, _13066_);
  nor _45560_ (_13068_, _00942_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nand _45561_ (_13069_, _00944_, _00537_);
  nand _45562_ (_13070_, _13069_, _26487_);
  nor _45563_ (_06627_, _13070_, _13068_);
  nand _45564_ (_13071_, _00840_, _12992_);
  nor _45565_ (_13072_, _13071_, _12990_);
  nor _45566_ (_13073_, _13072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand _45567_ (_13074_, _12999_, _00840_);
  nand _45568_ (_13075_, _13074_, _26487_);
  nor _45569_ (_06631_, _13075_, _13073_);
  nor _45570_ (_06634_, _03915_, rst);
  nand _45571_ (_13076_, _12688_, _25039_);
  nand _45572_ (_13077_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nand _45573_ (_06638_, _13077_, _13076_);
  nand _45574_ (_13078_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  nand _45575_ (_13079_, _03867_, _25150_);
  nand _45576_ (_06643_, _13079_, _13078_);
  nor _45577_ (_13080_, _28057_, _24059_);
  nand _45578_ (_13081_, _13080_, _25099_);
  not _45579_ (_13082_, _13080_);
  nand _45580_ (_13084_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nand _45581_ (_06646_, _13084_, _13081_);
  nand _45582_ (_13085_, _11937_, _25039_);
  nand _45583_ (_13086_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  nand _45584_ (_06650_, _13086_, _13085_);
  nand _45585_ (_13087_, _11937_, _25150_);
  nand _45586_ (_13088_, _11939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nand _45587_ (_06652_, _13088_, _13087_);
  nand _45588_ (_13089_, _12663_, _25150_);
  nand _45589_ (_13090_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nand _45590_ (_06655_, _13090_, _13089_);
  nor _45591_ (_13091_, _00287_, _25139_);
  not _45592_ (_13092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _45593_ (_13093_, _00271_, _13092_);
  nor _45594_ (_13094_, _00272_, _00304_);
  nor _45595_ (_13095_, _13094_, _13093_);
  nand _45596_ (_13096_, _13095_, _00287_);
  nand _45597_ (_13097_, _13096_, _00269_);
  nor _45598_ (_13098_, _13097_, _13091_);
  nor _45599_ (_13099_, _00297_, _13092_);
  nor _45600_ (_13100_, _13099_, _13098_);
  nor _45601_ (_06661_, _13100_, rst);
  nand _45602_ (_13101_, _04016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  nand _45603_ (_13102_, _04015_, _24927_);
  nand _45604_ (_06666_, _13102_, _13101_);
  nand _45605_ (_13103_, _11931_, _24830_);
  nand _45606_ (_13104_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nand _45607_ (_06669_, _13104_, _13103_);
  not _45608_ (_13105_, _06790_);
  not _45609_ (_13106_, _06723_);
  nor _45610_ (_13107_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  not _45611_ (_13108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nand _45612_ (_13109_, _06771_, _13108_);
  nand _45613_ (_13110_, _13109_, _06717_);
  nor _45614_ (_13111_, _13110_, _13107_);
  not _45615_ (_13112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  nor _45616_ (_13113_, _06774_, _13112_);
  not _45617_ (_13114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  nor _45618_ (_13115_, _06771_, _13114_);
  nor _45619_ (_13116_, _13115_, _13113_);
  nor _45620_ (_13117_, _13116_, _06717_);
  nor _45621_ (_13118_, _13117_, _13111_);
  nor _45622_ (_13119_, _13118_, _06751_);
  nand _45623_ (_13120_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  nand _45624_ (_13121_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nand _45625_ (_13122_, _13121_, _13120_);
  nand _45626_ (_13123_, _13122_, _06717_);
  nand _45627_ (_13124_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nand _45628_ (_13125_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  nand _45629_ (_13126_, _13125_, _13124_);
  nand _45630_ (_13127_, _13126_, _06716_);
  nand _45631_ (_13128_, _13127_, _13123_);
  nand _45632_ (_13129_, _13128_, _06751_);
  nand _45633_ (_13130_, _13129_, _06761_);
  nor _45634_ (_13131_, _13130_, _13119_);
  nor _45635_ (_13132_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  not _45636_ (_13133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  nand _45637_ (_13134_, _06774_, _13133_);
  nand _45638_ (_13135_, _13134_, _06716_);
  nor _45639_ (_13136_, _13135_, _13132_);
  nor _45640_ (_13137_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  not _45641_ (_13138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nand _45642_ (_13139_, _06771_, _13138_);
  nand _45643_ (_13140_, _13139_, _06717_);
  nor _45644_ (_13141_, _13140_, _13137_);
  nor _45645_ (_13142_, _13141_, _13136_);
  nor _45646_ (_13143_, _13142_, _06751_);
  nor _45647_ (_13144_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  nor _45648_ (_13145_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  nor _45649_ (_13146_, _13145_, _13144_);
  nand _45650_ (_13147_, _13146_, _06716_);
  nand _45651_ (_13148_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nand _45652_ (_13149_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nand _45653_ (_13150_, _13149_, _13148_);
  nand _45654_ (_13151_, _13150_, _06717_);
  nand _45655_ (_13152_, _13151_, _13147_);
  nand _45656_ (_13153_, _13152_, _06751_);
  nand _45657_ (_13154_, _13153_, _06760_);
  nor _45658_ (_13155_, _13154_, _13143_);
  nor _45659_ (_13156_, _13155_, _13131_);
  nand _45660_ (_13157_, _13156_, _06780_);
  nand _45661_ (_13158_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nand _45662_ (_13159_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nand _45663_ (_13160_, _13159_, _13158_);
  nand _45664_ (_13161_, _13160_, _06717_);
  nand _45665_ (_13162_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nand _45666_ (_13163_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  nand _45667_ (_13164_, _13163_, _13162_);
  nand _45668_ (_13165_, _13164_, _06716_);
  nand _45669_ (_13166_, _13165_, _13161_);
  nand _45670_ (_13167_, _13166_, _06748_);
  nand _45671_ (_13168_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  nand _45672_ (_13169_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nand _45673_ (_13170_, _13169_, _13168_);
  nand _45674_ (_13171_, _13170_, _06717_);
  nand _45675_ (_13172_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nand _45676_ (_13173_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  nand _45677_ (_13174_, _13173_, _13172_);
  nand _45678_ (_13175_, _13174_, _06716_);
  nand _45679_ (_13176_, _13175_, _13171_);
  nand _45680_ (_13177_, _13176_, _06751_);
  nand _45681_ (_13178_, _13177_, _13167_);
  nand _45682_ (_13179_, _13178_, _06761_);
  nor _45683_ (_13180_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  nor _45684_ (_13181_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  nor _45685_ (_13182_, _13181_, _13180_);
  nand _45686_ (_13183_, _13182_, _06717_);
  nor _45687_ (_13184_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  nor _45688_ (_13185_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nor _45689_ (_13186_, _13185_, _13184_);
  nand _45690_ (_13187_, _13186_, _06716_);
  nand _45691_ (_13188_, _13187_, _13183_);
  nand _45692_ (_13189_, _13188_, _06748_);
  not _45693_ (_13190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  nand _45694_ (_13191_, _06774_, _13190_);
  nor _45695_ (_13192_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nor _45696_ (_13193_, _13192_, _06716_);
  nand _45697_ (_13194_, _13193_, _13191_);
  nor _45698_ (_13195_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nor _45699_ (_13196_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nor _45700_ (_13197_, _13196_, _13195_);
  nand _45701_ (_13198_, _13197_, _06716_);
  nand _45702_ (_13199_, _13198_, _13194_);
  nand _45703_ (_13200_, _13199_, _06751_);
  nand _45704_ (_13201_, _13200_, _13189_);
  nand _45705_ (_13202_, _13201_, _06760_);
  nand _45706_ (_13203_, _13202_, _13179_);
  nand _45707_ (_13204_, _13203_, _06731_);
  nand _45708_ (_13205_, _13204_, _13157_);
  nand _45709_ (_13206_, _13205_, _06733_);
  nand _45710_ (_13207_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  nand _45711_ (_13208_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  nand _45712_ (_13209_, _13208_, _13207_);
  nand _45713_ (_13210_, _13209_, _06717_);
  nand _45714_ (_13211_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  nand _45715_ (_13212_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nand _45716_ (_13213_, _13212_, _13211_);
  nand _45717_ (_13214_, _13213_, _06716_);
  nand _45718_ (_13215_, _13214_, _13210_);
  nor _45719_ (_13216_, _13215_, _06751_);
  nor _45720_ (_13217_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  not _45721_ (_13218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  nand _45722_ (_13219_, _06771_, _13218_);
  nand _45723_ (_13220_, _13219_, _06717_);
  nor _45724_ (_13221_, _13220_, _13217_);
  not _45725_ (_13222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  nor _45726_ (_13223_, _06774_, _13222_);
  not _45727_ (_13224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nor _45728_ (_13225_, _06771_, _13224_);
  nor _45729_ (_13226_, _13225_, _13223_);
  nor _45730_ (_13227_, _13226_, _06717_);
  nor _45731_ (_13228_, _13227_, _13221_);
  nand _45732_ (_13229_, _13228_, _06751_);
  nand _45733_ (_13230_, _13229_, _06761_);
  nor _45734_ (_13231_, _13230_, _13216_);
  nor _45735_ (_13232_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nor _45736_ (_13233_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  nor _45737_ (_13234_, _13233_, _13232_);
  nand _45738_ (_13235_, _13234_, _06716_);
  nand _45739_ (_13236_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  nand _45740_ (_13237_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  nand _45741_ (_13238_, _13237_, _13236_);
  nand _45742_ (_13239_, _13238_, _06717_);
  nand _45743_ (_13240_, _13239_, _13235_);
  nor _45744_ (_13241_, _13240_, _06751_);
  nor _45745_ (_13242_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  not _45746_ (_13243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nand _45747_ (_13244_, _06774_, _13243_);
  nand _45748_ (_13245_, _13244_, _06716_);
  nor _45749_ (_13246_, _13245_, _13242_);
  nor _45750_ (_13247_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  not _45751_ (_13248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  nand _45752_ (_13249_, _06771_, _13248_);
  nand _45753_ (_13250_, _13249_, _06717_);
  nor _45754_ (_13251_, _13250_, _13247_);
  nor _45755_ (_13252_, _13251_, _13246_);
  nand _45756_ (_13253_, _13252_, _06751_);
  nand _45757_ (_13254_, _13253_, _06760_);
  nor _45758_ (_13255_, _13254_, _13241_);
  nor _45759_ (_13256_, _13255_, _13231_);
  nand _45760_ (_13258_, _13256_, _06780_);
  nand _45761_ (_13259_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  nand _45762_ (_13260_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  nand _45763_ (_13261_, _13260_, _13259_);
  nand _45764_ (_13262_, _13261_, _06717_);
  nand _45765_ (_13263_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  nand _45766_ (_13264_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nand _45767_ (_13265_, _13264_, _13263_);
  nand _45768_ (_13266_, _13265_, _06716_);
  nand _45769_ (_13267_, _13266_, _13262_);
  nand _45770_ (_13268_, _13267_, _06748_);
  nand _45771_ (_13269_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  nand _45772_ (_13270_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  nand _45773_ (_13271_, _13270_, _13269_);
  nand _45774_ (_13272_, _13271_, _06717_);
  nand _45775_ (_13273_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  nand _45776_ (_13274_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nand _45777_ (_13275_, _13274_, _13273_);
  nand _45778_ (_13276_, _13275_, _06716_);
  nand _45779_ (_13277_, _13276_, _13272_);
  nand _45780_ (_13279_, _13277_, _06751_);
  nand _45781_ (_13280_, _13279_, _13268_);
  nand _45782_ (_13281_, _13280_, _06761_);
  nor _45783_ (_13282_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nor _45784_ (_13283_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  nor _45785_ (_13284_, _13283_, _13282_);
  nand _45786_ (_13285_, _13284_, _06717_);
  nor _45787_ (_13286_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nor _45788_ (_13287_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  nor _45789_ (_13288_, _13287_, _13286_);
  nand _45790_ (_13289_, _13288_, _06716_);
  nand _45791_ (_13290_, _13289_, _13285_);
  nand _45792_ (_13291_, _13290_, _06748_);
  nor _45793_ (_13292_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  nor _45794_ (_13293_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  nor _45795_ (_13294_, _13293_, _13292_);
  nand _45796_ (_13295_, _13294_, _06717_);
  nor _45797_ (_13296_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  nor _45798_ (_13297_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nor _45799_ (_13298_, _13297_, _13296_);
  nand _45800_ (_13299_, _13298_, _06716_);
  nand _45801_ (_13300_, _13299_, _13295_);
  nand _45802_ (_13301_, _13300_, _06751_);
  nand _45803_ (_13302_, _13301_, _13291_);
  nand _45804_ (_13303_, _13302_, _06760_);
  nand _45805_ (_13304_, _13303_, _13281_);
  nor _45806_ (_13305_, _13304_, _06780_);
  nor _45807_ (_13306_, _13305_, _06733_);
  nand _45808_ (_13307_, _13306_, _13258_);
  nand _45809_ (_13308_, _13307_, _13206_);
  nand _45810_ (_13309_, _13308_, _13106_);
  nand _45811_ (_13310_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  nand _45812_ (_13311_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  nand _45813_ (_13312_, _13311_, _13310_);
  nand _45814_ (_13313_, _13312_, _06717_);
  nand _45815_ (_13314_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nand _45816_ (_13315_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  nand _45817_ (_13316_, _13315_, _13314_);
  nand _45818_ (_13317_, _13316_, _06716_);
  nand _45819_ (_13318_, _13317_, _13313_);
  nand _45820_ (_13319_, _13318_, _06751_);
  nand _45821_ (_13320_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  nand _45822_ (_13321_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  nand _45823_ (_13322_, _13321_, _13320_);
  nand _45824_ (_13323_, _13322_, _06717_);
  nand _45825_ (_13324_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  nand _45826_ (_13325_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  nand _45827_ (_13326_, _13325_, _13324_);
  nand _45828_ (_13327_, _13326_, _06716_);
  nand _45829_ (_13328_, _13327_, _13323_);
  nand _45830_ (_13329_, _13328_, _06748_);
  nand _45831_ (_13330_, _13329_, _13319_);
  nand _45832_ (_13331_, _13330_, _06761_);
  nor _45833_ (_13332_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  nor _45834_ (_13333_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  nor _45835_ (_13334_, _13333_, _13332_);
  nand _45836_ (_13335_, _13334_, _06716_);
  nand _45837_ (_13336_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nand _45838_ (_13337_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nand _45839_ (_13338_, _13337_, _13336_);
  nand _45840_ (_13339_, _13338_, _06717_);
  nand _45841_ (_13340_, _13339_, _13335_);
  nand _45842_ (_13341_, _13340_, _06751_);
  nor _45843_ (_13342_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nor _45844_ (_13343_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  nor _45845_ (_13344_, _13343_, _13342_);
  nand _45846_ (_13345_, _13344_, _06716_);
  nand _45847_ (_13346_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nand _45848_ (_13347_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  nand _45849_ (_13348_, _13347_, _13346_);
  nand _45850_ (_13349_, _13348_, _06717_);
  nand _45851_ (_13350_, _13349_, _13345_);
  nand _45852_ (_13351_, _13350_, _06748_);
  nand _45853_ (_13352_, _13351_, _13341_);
  nand _45854_ (_13353_, _13352_, _06760_);
  nand _45855_ (_13354_, _13353_, _13331_);
  nand _45856_ (_13355_, _13354_, _06780_);
  nand _45857_ (_13356_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nand _45858_ (_13357_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nand _45859_ (_13358_, _13357_, _13356_);
  nand _45860_ (_13360_, _13358_, _06717_);
  nand _45861_ (_13361_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  nand _45862_ (_13362_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  nand _45863_ (_13363_, _13362_, _13361_);
  nand _45864_ (_13364_, _13363_, _06716_);
  nand _45865_ (_13365_, _13364_, _13360_);
  nand _45866_ (_13366_, _13365_, _06751_);
  nand _45867_ (_13367_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  nand _45868_ (_13368_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  nand _45869_ (_13369_, _13368_, _13367_);
  nand _45870_ (_13370_, _13369_, _06717_);
  nand _45871_ (_13371_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  nand _45872_ (_13372_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  nand _45873_ (_13373_, _13372_, _13371_);
  nand _45874_ (_13374_, _13373_, _06716_);
  nand _45875_ (_13375_, _13374_, _13370_);
  nand _45876_ (_13376_, _13375_, _06748_);
  nand _45877_ (_13377_, _13376_, _13366_);
  nand _45878_ (_13378_, _13377_, _06761_);
  not _45879_ (_13379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nand _45880_ (_13380_, _06774_, _13379_);
  nor _45881_ (_13381_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  nor _45882_ (_13382_, _13381_, _06716_);
  nand _45883_ (_13383_, _13382_, _13380_);
  nor _45884_ (_13384_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  nor _45885_ (_13385_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  nor _45886_ (_13386_, _13385_, _13384_);
  nand _45887_ (_13387_, _13386_, _06716_);
  nand _45888_ (_13388_, _13387_, _13383_);
  nand _45889_ (_13389_, _13388_, _06751_);
  not _45890_ (_13390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nand _45891_ (_13391_, _06774_, _13390_);
  nor _45892_ (_13392_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nor _45893_ (_13393_, _13392_, _06716_);
  nand _45894_ (_13394_, _13393_, _13391_);
  nor _45895_ (_13395_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nor _45896_ (_13396_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  nor _45897_ (_13397_, _13396_, _13395_);
  nand _45898_ (_13398_, _13397_, _06716_);
  nand _45899_ (_13399_, _13398_, _13394_);
  nand _45900_ (_13400_, _13399_, _06748_);
  nand _45901_ (_13401_, _13400_, _13389_);
  nand _45902_ (_13402_, _13401_, _06760_);
  nand _45903_ (_13403_, _13402_, _13378_);
  nand _45904_ (_13404_, _13403_, _06731_);
  nand _45905_ (_13405_, _13404_, _13355_);
  nand _45906_ (_13406_, _13405_, _06733_);
  nand _45907_ (_13407_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  nand _45908_ (_13408_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nand _45909_ (_13409_, _13408_, _13407_);
  nand _45910_ (_13410_, _13409_, _06717_);
  nand _45911_ (_13411_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nand _45912_ (_13412_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  nand _45913_ (_13413_, _13412_, _13411_);
  nand _45914_ (_13414_, _13413_, _06716_);
  nand _45915_ (_13415_, _13414_, _13410_);
  nand _45916_ (_13416_, _13415_, _06748_);
  nand _45917_ (_13417_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  nand _45918_ (_13418_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nand _45919_ (_13419_, _13418_, _13417_);
  nand _45920_ (_13420_, _13419_, _06717_);
  nand _45921_ (_13421_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nand _45922_ (_13422_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  nand _45923_ (_13423_, _13422_, _13421_);
  nand _45924_ (_13424_, _13423_, _06716_);
  nand _45925_ (_13425_, _13424_, _13420_);
  nand _45926_ (_13426_, _13425_, _06751_);
  nand _45927_ (_13427_, _13426_, _13416_);
  nand _45928_ (_13428_, _13427_, _06761_);
  nor _45929_ (_13429_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nor _45930_ (_13430_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nor _45931_ (_13431_, _13430_, _13429_);
  nand _45932_ (_13432_, _13431_, _06716_);
  nand _45933_ (_13433_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nand _45934_ (_13434_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  nand _45935_ (_13435_, _13434_, _13433_);
  nand _45936_ (_13436_, _13435_, _06717_);
  nand _45937_ (_13437_, _13436_, _13432_);
  nand _45938_ (_13438_, _13437_, _06748_);
  nor _45939_ (_13439_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nor _45940_ (_13440_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  nor _45941_ (_13441_, _13440_, _13439_);
  nand _45942_ (_13442_, _13441_, _06716_);
  nand _45943_ (_13443_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  nand _45944_ (_13444_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  nand _45945_ (_13445_, _13444_, _13443_);
  nand _45946_ (_13446_, _13445_, _06717_);
  nand _45947_ (_13447_, _13446_, _13442_);
  nand _45948_ (_13448_, _13447_, _06751_);
  nand _45949_ (_13449_, _13448_, _13438_);
  nand _45950_ (_13450_, _13449_, _06760_);
  nand _45951_ (_13451_, _13450_, _13428_);
  nand _45952_ (_13452_, _13451_, _06780_);
  nand _45953_ (_13453_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nand _45954_ (_13454_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  nand _45955_ (_13455_, _13454_, _13453_);
  nand _45956_ (_13456_, _13455_, _06717_);
  nand _45957_ (_13457_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nand _45958_ (_13458_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nand _45959_ (_13459_, _13458_, _13457_);
  nand _45960_ (_13460_, _13459_, _06716_);
  nand _45961_ (_13461_, _13460_, _13456_);
  nand _45962_ (_13462_, _13461_, _06748_);
  nand _45963_ (_13463_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  nand _45964_ (_13464_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  nand _45965_ (_13465_, _13464_, _13463_);
  nand _45966_ (_13466_, _13465_, _06717_);
  nand _45967_ (_13467_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nand _45968_ (_13468_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nand _45969_ (_13469_, _13468_, _13467_);
  nand _45970_ (_13470_, _13469_, _06716_);
  nand _45971_ (_13471_, _13470_, _13466_);
  nand _45972_ (_13472_, _13471_, _06751_);
  nand _45973_ (_13473_, _13472_, _13462_);
  nand _45974_ (_13474_, _13473_, _06761_);
  nor _45975_ (_13475_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  nor _45976_ (_13476_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  nor _45977_ (_13477_, _13476_, _13475_);
  nand _45978_ (_13478_, _13477_, _06717_);
  nor _45979_ (_13479_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  nor _45980_ (_13480_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nor _45981_ (_13481_, _13480_, _13479_);
  nand _45982_ (_13482_, _13481_, _06716_);
  nand _45983_ (_13483_, _13482_, _13478_);
  nand _45984_ (_13484_, _13483_, _06748_);
  nor _45985_ (_13485_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nor _45986_ (_13486_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nor _45987_ (_13487_, _13486_, _13485_);
  nand _45988_ (_13488_, _13487_, _06717_);
  nor _45989_ (_13489_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  nor _45990_ (_13490_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  nor _45991_ (_13491_, _13490_, _13489_);
  nand _45992_ (_13492_, _13491_, _06716_);
  nand _45993_ (_13493_, _13492_, _13488_);
  nand _45994_ (_13494_, _13493_, _06751_);
  nand _45995_ (_13495_, _13494_, _13484_);
  nand _45996_ (_13496_, _13495_, _06760_);
  nand _45997_ (_13497_, _13496_, _13474_);
  nand _45998_ (_13498_, _13497_, _06731_);
  nand _45999_ (_13499_, _13498_, _13452_);
  nand _46000_ (_13500_, _13499_, _06734_);
  nand _46001_ (_13501_, _13500_, _13406_);
  nand _46002_ (_13502_, _13501_, _06723_);
  nand _46003_ (_13503_, _13502_, _13309_);
  nand _46004_ (_13504_, _13503_, _25929_);
  nor _46005_ (_13505_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  nor _46006_ (_13506_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nor _46007_ (_13507_, _13506_, _13505_);
  nand _46008_ (_13508_, _13507_, _06717_);
  nor _46009_ (_13509_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  nor _46010_ (_13510_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  nor _46011_ (_13511_, _13510_, _13509_);
  nand _46012_ (_13512_, _13511_, _06716_);
  nand _46013_ (_13513_, _13512_, _13508_);
  nand _46014_ (_13514_, _13513_, _06751_);
  nor _46015_ (_13515_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  nor _46016_ (_13516_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nor _46017_ (_13517_, _13516_, _13515_);
  nand _46018_ (_13518_, _13517_, _06717_);
  nor _46019_ (_13519_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nor _46020_ (_13520_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  nor _46021_ (_13521_, _13520_, _13519_);
  nand _46022_ (_13522_, _13521_, _06716_);
  nand _46023_ (_13523_, _13522_, _13518_);
  nand _46024_ (_13524_, _13523_, _06748_);
  nand _46025_ (_13525_, _13524_, _13514_);
  nand _46026_ (_13526_, _13525_, _06760_);
  nand _46027_ (_13527_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  nand _46028_ (_13528_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nand _46029_ (_13529_, _13528_, _13527_);
  nand _46030_ (_13530_, _13529_, _06717_);
  nand _46031_ (_13531_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nand _46032_ (_13532_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  nand _46033_ (_13533_, _13532_, _13531_);
  nand _46034_ (_13534_, _13533_, _06716_);
  nand _46035_ (_13535_, _13534_, _13530_);
  nand _46036_ (_13536_, _13535_, _06751_);
  nand _46037_ (_13537_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  nand _46038_ (_13538_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nand _46039_ (_13539_, _13538_, _13537_);
  nand _46040_ (_13540_, _13539_, _06717_);
  nand _46041_ (_13541_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nand _46042_ (_13542_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  nand _46043_ (_13543_, _13542_, _13541_);
  nand _46044_ (_13544_, _13543_, _06716_);
  nand _46045_ (_13545_, _13544_, _13540_);
  nand _46046_ (_13546_, _13545_, _06748_);
  nand _46047_ (_13547_, _13546_, _13536_);
  nand _46048_ (_13548_, _13547_, _06761_);
  nand _46049_ (_13549_, _13548_, _13526_);
  nand _46050_ (_13550_, _13549_, _06731_);
  nor _46051_ (_13551_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _46052_ (_13552_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor _46053_ (_13553_, _13552_, _13551_);
  nand _46054_ (_13554_, _13553_, _06716_);
  nand _46055_ (_13555_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nand _46056_ (_13556_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nand _46057_ (_13557_, _13556_, _13555_);
  nand _46058_ (_13558_, _13557_, _06717_);
  nand _46059_ (_13559_, _13558_, _13554_);
  nand _46060_ (_13560_, _13559_, _06751_);
  nor _46061_ (_13561_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _46062_ (_13562_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _46063_ (_13563_, _13562_, _13561_);
  nand _46064_ (_13564_, _13563_, _06716_);
  nand _46065_ (_13565_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nand _46066_ (_13566_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nand _46067_ (_13567_, _13566_, _13565_);
  nand _46068_ (_13568_, _13567_, _06717_);
  nand _46069_ (_13569_, _13568_, _13564_);
  nand _46070_ (_13570_, _13569_, _06748_);
  nand _46071_ (_13571_, _13570_, _13560_);
  nand _46072_ (_13572_, _13571_, _06760_);
  nand _46073_ (_13573_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand _46074_ (_13574_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nand _46075_ (_13575_, _13574_, _13573_);
  nand _46076_ (_13576_, _13575_, _06717_);
  nand _46077_ (_13577_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nand _46078_ (_13578_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nand _46079_ (_13579_, _13578_, _13577_);
  nand _46080_ (_13580_, _13579_, _06716_);
  nand _46081_ (_13581_, _13580_, _13576_);
  nand _46082_ (_13582_, _13581_, _06751_);
  nand _46083_ (_13583_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nand _46084_ (_13584_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nand _46085_ (_13585_, _13584_, _13583_);
  nand _46086_ (_13586_, _13585_, _06717_);
  nand _46087_ (_13587_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nand _46088_ (_13588_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nand _46089_ (_13589_, _13588_, _13587_);
  nand _46090_ (_13591_, _13589_, _06716_);
  nand _46091_ (_13592_, _13591_, _13586_);
  nand _46092_ (_13593_, _13592_, _06748_);
  nand _46093_ (_13594_, _13593_, _13582_);
  nand _46094_ (_13595_, _13594_, _06761_);
  nand _46095_ (_13596_, _13595_, _13572_);
  nand _46096_ (_13597_, _13596_, _06780_);
  nand _46097_ (_13598_, _13597_, _13550_);
  nand _46098_ (_13599_, _13598_, _06733_);
  nand _46099_ (_13600_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nand _46100_ (_13601_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nand _46101_ (_13602_, _13601_, _13600_);
  nand _46102_ (_13603_, _13602_, _06717_);
  nand _46103_ (_13604_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  nand _46104_ (_13605_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  nand _46105_ (_13606_, _13605_, _13604_);
  nand _46106_ (_13607_, _13606_, _06716_);
  nand _46107_ (_13608_, _13607_, _13603_);
  nand _46108_ (_13609_, _13608_, _06748_);
  nand _46109_ (_13610_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nand _46110_ (_13612_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nand _46111_ (_13613_, _13612_, _13610_);
  nand _46112_ (_13614_, _13613_, _06717_);
  nand _46113_ (_13615_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  nand _46114_ (_13616_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nand _46115_ (_13617_, _13616_, _13615_);
  nand _46116_ (_13618_, _13617_, _06716_);
  nand _46117_ (_13619_, _13618_, _13614_);
  nand _46118_ (_13620_, _13619_, _06751_);
  nand _46119_ (_13621_, _13620_, _13609_);
  nand _46120_ (_13622_, _13621_, _06761_);
  nor _46121_ (_13623_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nor _46122_ (_13624_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  nor _46123_ (_13625_, _13624_, _13623_);
  nand _46124_ (_13626_, _13625_, _06716_);
  nand _46125_ (_13627_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  nand _46126_ (_13628_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  nand _46127_ (_13629_, _13628_, _13627_);
  nand _46128_ (_13630_, _13629_, _06717_);
  nand _46129_ (_13631_, _13630_, _13626_);
  nand _46130_ (_13633_, _13631_, _06748_);
  nor _46131_ (_13634_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nor _46132_ (_13635_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nor _46133_ (_13636_, _13635_, _13634_);
  nand _46134_ (_13637_, _13636_, _06716_);
  nand _46135_ (_13638_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nand _46136_ (_13639_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  nand _46137_ (_13640_, _13639_, _13638_);
  nand _46138_ (_13641_, _13640_, _06717_);
  nand _46139_ (_13642_, _13641_, _13637_);
  nand _46140_ (_13643_, _13642_, _06751_);
  nand _46141_ (_13644_, _13643_, _13633_);
  nand _46142_ (_13645_, _13644_, _06760_);
  nand _46143_ (_13646_, _13645_, _13622_);
  nand _46144_ (_13647_, _13646_, _06780_);
  nand _46145_ (_13648_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  nand _46146_ (_13649_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nand _46147_ (_13650_, _13649_, _13648_);
  nand _46148_ (_13651_, _13650_, _06717_);
  nand _46149_ (_13652_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  nand _46150_ (_13654_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  nand _46151_ (_13655_, _13654_, _13652_);
  nand _46152_ (_13656_, _13655_, _06716_);
  nand _46153_ (_13657_, _13656_, _13651_);
  nand _46154_ (_13658_, _13657_, _06748_);
  nand _46155_ (_13659_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nand _46156_ (_13660_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  nand _46157_ (_13661_, _13660_, _13659_);
  nand _46158_ (_13662_, _13661_, _06717_);
  nand _46159_ (_13663_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nand _46160_ (_13664_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nand _46161_ (_13665_, _13664_, _13663_);
  nand _46162_ (_13666_, _13665_, _06716_);
  nand _46163_ (_13667_, _13666_, _13662_);
  nand _46164_ (_13668_, _13667_, _06751_);
  nand _46165_ (_13669_, _13668_, _13658_);
  nand _46166_ (_13670_, _13669_, _06761_);
  nor _46167_ (_13671_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  nor _46168_ (_13672_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nor _46169_ (_13673_, _13672_, _13671_);
  nand _46170_ (_13675_, _13673_, _06717_);
  nor _46171_ (_13676_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nor _46172_ (_13677_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  nor _46173_ (_13678_, _13677_, _13676_);
  nand _46174_ (_13679_, _13678_, _06716_);
  nand _46175_ (_13680_, _13679_, _13675_);
  nand _46176_ (_13681_, _13680_, _06748_);
  nor _46177_ (_13682_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  nor _46178_ (_13683_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nor _46179_ (_13684_, _13683_, _13682_);
  nand _46180_ (_13685_, _13684_, _06717_);
  nor _46181_ (_13686_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  nor _46182_ (_13687_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  nor _46183_ (_13688_, _13687_, _13686_);
  nand _46184_ (_13689_, _13688_, _06716_);
  nand _46185_ (_13690_, _13689_, _13685_);
  nand _46186_ (_13691_, _13690_, _06751_);
  nand _46187_ (_13692_, _13691_, _13681_);
  nand _46188_ (_13693_, _13692_, _06760_);
  nand _46189_ (_13694_, _13693_, _13670_);
  nand _46190_ (_13696_, _13694_, _06731_);
  nand _46191_ (_13697_, _13696_, _13647_);
  nand _46192_ (_13698_, _13697_, _06734_);
  nand _46193_ (_13699_, _13698_, _13599_);
  nand _46194_ (_13700_, _13699_, _13106_);
  nand _46195_ (_13701_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nand _46196_ (_13702_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  nand _46197_ (_13703_, _13702_, _13701_);
  nand _46198_ (_13704_, _13703_, _06716_);
  nand _46199_ (_13705_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  nand _46200_ (_13706_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  nand _46201_ (_13707_, _13706_, _13705_);
  nand _46202_ (_13708_, _13707_, _06717_);
  nand _46203_ (_13709_, _13708_, _13704_);
  nand _46204_ (_13710_, _13709_, _06748_);
  nand _46205_ (_13711_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  nand _46206_ (_13712_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nand _46207_ (_13713_, _13712_, _13711_);
  nand _46208_ (_13714_, _13713_, _06716_);
  nand _46209_ (_13715_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nand _46210_ (_13716_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nand _46211_ (_13717_, _13716_, _13715_);
  nand _46212_ (_13718_, _13717_, _06717_);
  nand _46213_ (_13719_, _13718_, _13714_);
  nand _46214_ (_13720_, _13719_, _06751_);
  nand _46215_ (_13721_, _13720_, _13710_);
  nand _46216_ (_13722_, _13721_, _06761_);
  nand _46217_ (_13723_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  nand _46218_ (_13724_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nand _46219_ (_13725_, _13724_, _13723_);
  nand _46220_ (_13726_, _13725_, _06717_);
  nor _46221_ (_13727_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  nor _46222_ (_13728_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nor _46223_ (_13729_, _13728_, _13727_);
  nand _46224_ (_13730_, _13729_, _06716_);
  nand _46225_ (_13731_, _13730_, _13726_);
  nand _46226_ (_13732_, _13731_, _06748_);
  nand _46227_ (_13733_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  nand _46228_ (_13734_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nand _46229_ (_13735_, _13734_, _13733_);
  nand _46230_ (_13736_, _13735_, _06717_);
  nor _46231_ (_13737_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  nor _46232_ (_13738_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nor _46233_ (_13739_, _13738_, _13737_);
  nand _46234_ (_13740_, _13739_, _06716_);
  nand _46235_ (_13741_, _13740_, _13736_);
  nand _46236_ (_13742_, _13741_, _06751_);
  nand _46237_ (_13743_, _13742_, _13732_);
  nand _46238_ (_13744_, _13743_, _06760_);
  nand _46239_ (_13745_, _13744_, _13722_);
  nand _46240_ (_13746_, _13745_, _06780_);
  nand _46241_ (_13747_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  nand _46242_ (_13748_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nand _46243_ (_13749_, _13748_, _13747_);
  nand _46244_ (_13750_, _13749_, _06717_);
  nand _46245_ (_13751_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  nand _46246_ (_13752_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  nand _46247_ (_13753_, _13752_, _13751_);
  nand _46248_ (_13754_, _13753_, _06716_);
  nand _46249_ (_13755_, _13754_, _13750_);
  nand _46250_ (_13756_, _13755_, _06748_);
  nand _46251_ (_13757_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nand _46252_ (_13758_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  nand _46253_ (_13759_, _13758_, _13757_);
  nand _46254_ (_13760_, _13759_, _06717_);
  nand _46255_ (_13761_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  nand _46256_ (_13762_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nand _46257_ (_13763_, _13762_, _13761_);
  nand _46258_ (_13764_, _13763_, _06716_);
  nand _46259_ (_13765_, _13764_, _13760_);
  nand _46260_ (_13766_, _13765_, _06751_);
  nand _46261_ (_13767_, _13766_, _13756_);
  nand _46262_ (_13768_, _13767_, _06761_);
  nor _46263_ (_13769_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nor _46264_ (_13770_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  nor _46265_ (_13771_, _13770_, _13769_);
  nor _46266_ (_13772_, _13771_, _06716_);
  nor _46267_ (_13773_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  nor _46268_ (_13774_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nor _46269_ (_13775_, _13774_, _13773_);
  nor _46270_ (_13776_, _13775_, _06717_);
  nor _46271_ (_13777_, _13776_, _13772_);
  nand _46272_ (_13778_, _13777_, _06748_);
  nor _46273_ (_13779_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nor _46274_ (_13780_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nor _46275_ (_13781_, _13780_, _13779_);
  nand _46276_ (_13782_, _13781_, _06717_);
  nor _46277_ (_13783_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  nor _46278_ (_13784_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  nor _46279_ (_13785_, _13784_, _13783_);
  nand _46280_ (_13786_, _13785_, _06716_);
  nand _46281_ (_13787_, _13786_, _13782_);
  nand _46282_ (_13788_, _13787_, _06751_);
  nand _46283_ (_13789_, _13788_, _13778_);
  nand _46284_ (_13790_, _13789_, _06760_);
  nand _46285_ (_13791_, _13790_, _13768_);
  nand _46286_ (_13792_, _13791_, _06731_);
  nand _46287_ (_13793_, _13792_, _13746_);
  nand _46288_ (_13794_, _13793_, _06734_);
  not _46289_ (_13795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  nand _46290_ (_13796_, _06774_, _13795_);
  nor _46291_ (_13797_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  nor _46292_ (_13798_, _13797_, _06716_);
  nand _46293_ (_13799_, _13798_, _13796_);
  nor _46294_ (_13800_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nor _46295_ (_13801_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nor _46296_ (_13802_, _13801_, _13800_);
  nand _46297_ (_13803_, _13802_, _06716_);
  nand _46298_ (_13804_, _13803_, _13799_);
  nand _46299_ (_13805_, _13804_, _06751_);
  not _46300_ (_13806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  nand _46301_ (_13807_, _06774_, _13806_);
  nor _46302_ (_13808_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nor _46303_ (_13809_, _13808_, _06716_);
  nand _46304_ (_13810_, _13809_, _13807_);
  nor _46305_ (_13811_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nor _46306_ (_13812_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nor _46307_ (_13813_, _13812_, _13811_);
  nand _46308_ (_13814_, _13813_, _06716_);
  nand _46309_ (_13815_, _13814_, _13810_);
  nand _46310_ (_13816_, _13815_, _06748_);
  nand _46311_ (_13817_, _13816_, _13805_);
  nand _46312_ (_13818_, _13817_, _06760_);
  nand _46313_ (_13819_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nand _46314_ (_13820_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  nand _46315_ (_13821_, _13820_, _13819_);
  nand _46316_ (_13822_, _13821_, _06717_);
  nand _46317_ (_13823_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  nand _46318_ (_13824_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nand _46319_ (_13825_, _13824_, _13823_);
  nand _46320_ (_13826_, _13825_, _06716_);
  nand _46321_ (_13827_, _13826_, _13822_);
  nand _46322_ (_13828_, _13827_, _06751_);
  nand _46323_ (_13829_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  nand _46324_ (_13830_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nand _46325_ (_13831_, _13830_, _13829_);
  nand _46326_ (_13832_, _13831_, _06717_);
  nand _46327_ (_13833_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  nand _46328_ (_13834_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  nand _46329_ (_13835_, _13834_, _13833_);
  nand _46330_ (_13836_, _13835_, _06716_);
  nand _46331_ (_13837_, _13836_, _13832_);
  nand _46332_ (_13838_, _13837_, _06748_);
  nand _46333_ (_13839_, _13838_, _13828_);
  nand _46334_ (_13840_, _13839_, _06761_);
  nand _46335_ (_13841_, _13840_, _13818_);
  nand _46336_ (_13842_, _13841_, _06731_);
  nor _46337_ (_13843_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nor _46338_ (_13844_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nor _46339_ (_13845_, _13844_, _13843_);
  nand _46340_ (_13846_, _13845_, _06717_);
  nor _46341_ (_13847_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nor _46342_ (_13848_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  nor _46343_ (_13849_, _13848_, _13847_);
  nand _46344_ (_13850_, _13849_, _06716_);
  nand _46345_ (_13851_, _13850_, _13846_);
  nand _46346_ (_13852_, _13851_, _06751_);
  not _46347_ (_13853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  nand _46348_ (_13854_, _06774_, _13853_);
  not _46349_ (_13855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  nand _46350_ (_13856_, _06771_, _13855_);
  nand _46351_ (_13857_, _13856_, _13854_);
  nand _46352_ (_13858_, _13857_, _06716_);
  nor _46353_ (_13859_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nor _46354_ (_13860_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nor _46355_ (_13861_, _13860_, _13859_);
  nor _46356_ (_13862_, _13861_, _06716_);
  nor _46357_ (_13863_, _13862_, _06751_);
  nand _46358_ (_13864_, _13863_, _13858_);
  nand _46359_ (_13865_, _13864_, _13852_);
  nand _46360_ (_13866_, _13865_, _06760_);
  nand _46361_ (_13867_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  nand _46362_ (_13868_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nand _46363_ (_13869_, _13868_, _13867_);
  nand _46364_ (_13870_, _13869_, _06717_);
  nand _46365_ (_13871_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  nand _46366_ (_13872_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  nand _46367_ (_13873_, _13872_, _13871_);
  nand _46368_ (_13874_, _13873_, _06716_);
  nand _46369_ (_13875_, _13874_, _13870_);
  nand _46370_ (_13876_, _13875_, _06751_);
  nand _46371_ (_13877_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  not _46372_ (_13878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nor _46373_ (_13879_, _06771_, _13878_);
  nor _46374_ (_13880_, _13879_, _06716_);
  nand _46375_ (_13881_, _13880_, _13877_);
  not _46376_ (_13882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  nor _46377_ (_13883_, _06771_, _13882_);
  nand _46378_ (_13884_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  nand _46379_ (_13885_, _13884_, _06716_);
  nor _46380_ (_13887_, _13885_, _13883_);
  nor _46381_ (_13888_, _13887_, _06751_);
  nand _46382_ (_13889_, _13888_, _13881_);
  nand _46383_ (_13890_, _13889_, _13876_);
  nand _46384_ (_13891_, _13890_, _06761_);
  nand _46385_ (_13892_, _13891_, _13866_);
  nand _46386_ (_13893_, _13892_, _06780_);
  nand _46387_ (_13894_, _13893_, _13842_);
  nand _46388_ (_13895_, _13894_, _06733_);
  nand _46389_ (_13896_, _13895_, _13794_);
  nand _46390_ (_13897_, _13896_, _06723_);
  nand _46391_ (_13898_, _13897_, _13700_);
  nand _46392_ (_13899_, _13898_, _25843_);
  nand _46393_ (_13900_, _13899_, _13504_);
  nor _46394_ (_13901_, _13900_, _13105_);
  nand _46395_ (_13902_, _13105_, _24263_);
  nand _46396_ (_13903_, _13902_, _26487_);
  nor _46397_ (_06670_, _13903_, _13901_);
  nand _46398_ (_13904_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nand _46399_ (_13905_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nand _46400_ (_13907_, _13905_, _13904_);
  nand _46401_ (_13908_, _13907_, _06716_);
  nand _46402_ (_13909_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  nand _46403_ (_13910_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  nand _46404_ (_13911_, _13910_, _13909_);
  nand _46405_ (_13912_, _13911_, _06717_);
  nand _46406_ (_13913_, _13912_, _13908_);
  nand _46407_ (_13914_, _13913_, _06748_);
  nand _46408_ (_13915_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nand _46409_ (_13916_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nand _46410_ (_13917_, _13916_, _13915_);
  nand _46411_ (_13918_, _13917_, _06716_);
  nand _46412_ (_13919_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  nand _46413_ (_13920_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  nand _46414_ (_13921_, _13920_, _13919_);
  nand _46415_ (_13922_, _13921_, _06717_);
  nand _46416_ (_13923_, _13922_, _13918_);
  nand _46417_ (_13924_, _13923_, _06751_);
  nand _46418_ (_13925_, _13924_, _13914_);
  nand _46419_ (_13926_, _13925_, _06761_);
  nand _46420_ (_13927_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  nand _46421_ (_13928_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  nand _46422_ (_13929_, _13928_, _13927_);
  nand _46423_ (_13930_, _13929_, _06717_);
  nor _46424_ (_13931_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nor _46425_ (_13932_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nor _46426_ (_13933_, _13932_, _13931_);
  nand _46427_ (_13934_, _13933_, _06716_);
  nand _46428_ (_13935_, _13934_, _13930_);
  nand _46429_ (_13936_, _13935_, _06748_);
  nand _46430_ (_13937_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  nand _46431_ (_13938_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  nand _46432_ (_13939_, _13938_, _13937_);
  nand _46433_ (_13940_, _13939_, _06717_);
  nor _46434_ (_13941_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nor _46435_ (_13942_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  nor _46436_ (_13943_, _13942_, _13941_);
  nand _46437_ (_13944_, _13943_, _06716_);
  nand _46438_ (_13945_, _13944_, _13940_);
  nand _46439_ (_13946_, _13945_, _06751_);
  nand _46440_ (_13947_, _13946_, _13936_);
  nand _46441_ (_13948_, _13947_, _06760_);
  nand _46442_ (_13949_, _13948_, _13926_);
  nand _46443_ (_13950_, _13949_, _06780_);
  nand _46444_ (_13951_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nand _46445_ (_13952_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nand _46446_ (_13953_, _13952_, _13951_);
  nand _46447_ (_13954_, _13953_, _06717_);
  nand _46448_ (_13955_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nand _46449_ (_13956_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  nand _46450_ (_13957_, _13956_, _13955_);
  nand _46451_ (_13958_, _13957_, _06716_);
  nand _46452_ (_13959_, _13958_, _13954_);
  nand _46453_ (_13960_, _13959_, _06748_);
  nand _46454_ (_13961_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  nand _46455_ (_13962_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nand _46456_ (_13963_, _13962_, _13961_);
  nand _46457_ (_13964_, _13963_, _06717_);
  nand _46458_ (_13965_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  nand _46459_ (_13966_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  nand _46460_ (_13967_, _13966_, _13965_);
  nand _46461_ (_13968_, _13967_, _06716_);
  nand _46462_ (_13969_, _13968_, _13964_);
  nand _46463_ (_13970_, _13969_, _06751_);
  nand _46464_ (_13971_, _13970_, _13960_);
  nand _46465_ (_13972_, _13971_, _06761_);
  nor _46466_ (_13973_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nor _46467_ (_13974_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nor _46468_ (_13975_, _13974_, _13973_);
  nand _46469_ (_13976_, _13975_, _06717_);
  nor _46470_ (_13977_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nor _46471_ (_13978_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  nor _46472_ (_13979_, _13978_, _13977_);
  nand _46473_ (_13980_, _13979_, _06716_);
  nand _46474_ (_13981_, _13980_, _13976_);
  nand _46475_ (_13982_, _13981_, _06748_);
  nor _46476_ (_13983_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  nor _46477_ (_13984_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  nor _46478_ (_13985_, _13984_, _13983_);
  nor _46479_ (_13986_, _13985_, _06716_);
  nor _46480_ (_13988_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nor _46481_ (_13989_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nor _46482_ (_13990_, _13989_, _13988_);
  nor _46483_ (_13991_, _13990_, _06717_);
  nor _46484_ (_13992_, _13991_, _13986_);
  nand _46485_ (_13993_, _13992_, _06751_);
  nand _46486_ (_13994_, _13993_, _13982_);
  nand _46487_ (_13995_, _13994_, _06760_);
  nand _46488_ (_13996_, _13995_, _13972_);
  nand _46489_ (_13997_, _13996_, _06731_);
  nand _46490_ (_13998_, _13997_, _13950_);
  nand _46491_ (_13999_, _13998_, _06734_);
  nand _46492_ (_14000_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nand _46493_ (_14001_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand _46494_ (_14002_, _14001_, _14000_);
  nand _46495_ (_14003_, _14002_, _06717_);
  nand _46496_ (_14004_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nand _46497_ (_14005_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand _46498_ (_14006_, _14005_, _14004_);
  nand _46499_ (_14007_, _14006_, _06716_);
  nand _46500_ (_14008_, _14007_, _14003_);
  nand _46501_ (_14009_, _14008_, _06748_);
  nand _46502_ (_14010_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nand _46503_ (_14011_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand _46504_ (_14012_, _14011_, _14010_);
  nand _46505_ (_14013_, _14012_, _06717_);
  nand _46506_ (_14014_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nand _46507_ (_14015_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand _46508_ (_14016_, _14015_, _14014_);
  nand _46509_ (_14017_, _14016_, _06716_);
  nand _46510_ (_14018_, _14017_, _14013_);
  nand _46511_ (_14019_, _14018_, _06751_);
  nand _46512_ (_14020_, _14019_, _14009_);
  nand _46513_ (_14021_, _14020_, _06761_);
  nor _46514_ (_14022_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _46515_ (_14023_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _46516_ (_14024_, _14023_, _14022_);
  nand _46517_ (_14025_, _14024_, _06717_);
  nor _46518_ (_14026_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _46519_ (_14027_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _46520_ (_14028_, _14027_, _14026_);
  nand _46521_ (_14029_, _14028_, _06716_);
  nand _46522_ (_14030_, _14029_, _14025_);
  nand _46523_ (_14031_, _14030_, _06748_);
  nor _46524_ (_14032_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _46525_ (_14033_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor _46526_ (_14034_, _14033_, _14032_);
  nand _46527_ (_14035_, _14034_, _06717_);
  nor _46528_ (_14036_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor _46529_ (_14037_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _46530_ (_14038_, _14037_, _14036_);
  nand _46531_ (_14039_, _14038_, _06716_);
  nand _46532_ (_14040_, _14039_, _14035_);
  nand _46533_ (_14041_, _14040_, _06751_);
  nand _46534_ (_14042_, _14041_, _14031_);
  nand _46535_ (_14043_, _14042_, _06760_);
  nand _46536_ (_14044_, _14043_, _14021_);
  nand _46537_ (_14045_, _14044_, _06780_);
  nand _46538_ (_14046_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nand _46539_ (_14047_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nand _46540_ (_14048_, _14047_, _14046_);
  nand _46541_ (_14049_, _14048_, _06717_);
  nand _46542_ (_14050_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nand _46543_ (_14051_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  nand _46544_ (_14052_, _14051_, _14050_);
  nand _46545_ (_14053_, _14052_, _06716_);
  nand _46546_ (_14054_, _14053_, _14049_);
  nand _46547_ (_14055_, _14054_, _06748_);
  nand _46548_ (_14056_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  nand _46549_ (_14057_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nand _46550_ (_14058_, _14057_, _14056_);
  nand _46551_ (_14059_, _14058_, _06717_);
  nand _46552_ (_14060_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nand _46553_ (_14061_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  nand _46554_ (_14062_, _14061_, _14060_);
  nand _46555_ (_14063_, _14062_, _06716_);
  nand _46556_ (_14064_, _14063_, _14059_);
  nand _46557_ (_14065_, _14064_, _06751_);
  nand _46558_ (_14066_, _14065_, _14055_);
  nand _46559_ (_14067_, _14066_, _06761_);
  nor _46560_ (_14068_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  nor _46561_ (_14069_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nor _46562_ (_14070_, _14069_, _14068_);
  nand _46563_ (_14071_, _14070_, _06717_);
  nor _46564_ (_14072_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nor _46565_ (_14073_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  nor _46566_ (_14074_, _14073_, _14072_);
  nand _46567_ (_14075_, _14074_, _06716_);
  nand _46568_ (_14076_, _14075_, _14071_);
  nand _46569_ (_14077_, _14076_, _06748_);
  nor _46570_ (_14078_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  nor _46571_ (_14079_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nor _46572_ (_14080_, _14079_, _14078_);
  nand _46573_ (_14081_, _14080_, _06717_);
  nor _46574_ (_14082_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nor _46575_ (_14083_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  nor _46576_ (_14084_, _14083_, _14082_);
  nand _46577_ (_14085_, _14084_, _06716_);
  nand _46578_ (_14086_, _14085_, _14081_);
  nand _46579_ (_14087_, _14086_, _06751_);
  nand _46580_ (_14088_, _14087_, _14077_);
  nand _46581_ (_14089_, _14088_, _06760_);
  nand _46582_ (_14090_, _14089_, _14067_);
  nand _46583_ (_14091_, _14090_, _06731_);
  nand _46584_ (_14092_, _14091_, _14045_);
  nand _46585_ (_14093_, _14092_, _06733_);
  nand _46586_ (_14094_, _14093_, _13999_);
  nor _46587_ (_14095_, _14094_, _06723_);
  nand _46588_ (_14096_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  nand _46589_ (_14097_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  nand _46590_ (_14098_, _14097_, _14096_);
  nand _46591_ (_14099_, _14098_, _06717_);
  nand _46592_ (_14100_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nand _46593_ (_14101_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nand _46594_ (_14102_, _14101_, _14100_);
  nand _46595_ (_14103_, _14102_, _06716_);
  nand _46596_ (_14104_, _14103_, _14099_);
  nand _46597_ (_14105_, _14104_, _06748_);
  nand _46598_ (_14106_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  nand _46599_ (_14107_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  nand _46600_ (_14108_, _14107_, _14106_);
  nand _46601_ (_14109_, _14108_, _06717_);
  nand _46602_ (_14110_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  nand _46603_ (_14111_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  nand _46604_ (_14112_, _14111_, _14110_);
  nand _46605_ (_14113_, _14112_, _06716_);
  nand _46606_ (_14114_, _14113_, _14109_);
  nand _46607_ (_14115_, _14114_, _06751_);
  nand _46608_ (_14116_, _14115_, _14105_);
  nand _46609_ (_14117_, _14116_, _06761_);
  nor _46610_ (_14119_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  nor _46611_ (_14120_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  nor _46612_ (_14121_, _14120_, _14119_);
  nand _46613_ (_14122_, _14121_, _06716_);
  nand _46614_ (_14123_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  nand _46615_ (_14124_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nand _46616_ (_14125_, _14124_, _14123_);
  nand _46617_ (_14126_, _14125_, _06717_);
  nand _46618_ (_14127_, _14126_, _14122_);
  nand _46619_ (_14128_, _14127_, _06748_);
  nor _46620_ (_14129_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nor _46621_ (_14130_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nor _46622_ (_14131_, _14130_, _14129_);
  nand _46623_ (_14132_, _14131_, _06716_);
  nand _46624_ (_14133_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  nand _46625_ (_14134_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  nand _46626_ (_14135_, _14134_, _14133_);
  nand _46627_ (_14136_, _14135_, _06717_);
  nand _46628_ (_14137_, _14136_, _14132_);
  nand _46629_ (_14138_, _14137_, _06751_);
  nand _46630_ (_14139_, _14138_, _14128_);
  nand _46631_ (_14140_, _14139_, _06760_);
  nand _46632_ (_14141_, _14140_, _14117_);
  nand _46633_ (_14142_, _14141_, _06780_);
  nand _46634_ (_14143_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  nand _46635_ (_14144_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  nand _46636_ (_14145_, _14144_, _14143_);
  nand _46637_ (_14146_, _14145_, _06717_);
  nand _46638_ (_14147_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  nand _46639_ (_14148_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nand _46640_ (_14149_, _14148_, _14147_);
  nand _46641_ (_14150_, _14149_, _06716_);
  nand _46642_ (_14151_, _14150_, _14146_);
  nand _46643_ (_14152_, _14151_, _06748_);
  nand _46644_ (_14153_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nand _46645_ (_14154_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  nand _46646_ (_14155_, _14154_, _14153_);
  nand _46647_ (_14156_, _14155_, _06717_);
  nand _46648_ (_14157_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  nand _46649_ (_14158_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nand _46650_ (_14159_, _14158_, _14157_);
  nand _46651_ (_14160_, _14159_, _06716_);
  nand _46652_ (_14161_, _14160_, _14156_);
  nand _46653_ (_14162_, _14161_, _06751_);
  nand _46654_ (_14163_, _14162_, _14152_);
  nand _46655_ (_14164_, _14163_, _06761_);
  nor _46656_ (_14165_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nor _46657_ (_14166_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  nor _46658_ (_14167_, _14166_, _14165_);
  nand _46659_ (_14168_, _14167_, _06717_);
  nor _46660_ (_14169_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nor _46661_ (_14170_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nor _46662_ (_14171_, _14170_, _14169_);
  nand _46663_ (_14172_, _14171_, _06716_);
  nand _46664_ (_14173_, _14172_, _14168_);
  nand _46665_ (_14174_, _14173_, _06748_);
  nor _46666_ (_14175_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  nor _46667_ (_14176_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nor _46668_ (_14177_, _14176_, _14175_);
  nand _46669_ (_14178_, _14177_, _06717_);
  nor _46670_ (_14179_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  nor _46671_ (_14180_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  nor _46672_ (_14181_, _14180_, _14179_);
  nand _46673_ (_14182_, _14181_, _06716_);
  nand _46674_ (_14183_, _14182_, _14178_);
  nand _46675_ (_14184_, _14183_, _06751_);
  nand _46676_ (_14185_, _14184_, _14174_);
  nand _46677_ (_14186_, _14185_, _06760_);
  nand _46678_ (_14187_, _14186_, _14164_);
  nand _46679_ (_14188_, _14187_, _06731_);
  nand _46680_ (_14189_, _14188_, _14142_);
  nand _46681_ (_14190_, _14189_, _06734_);
  nor _46682_ (_14191_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  nor _46683_ (_14192_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nor _46684_ (_14193_, _14192_, _14191_);
  nand _46685_ (_14194_, _14193_, _06717_);
  nor _46686_ (_14195_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  nor _46687_ (_14196_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  nor _46688_ (_14197_, _14196_, _14195_);
  nand _46689_ (_14198_, _14197_, _06716_);
  nand _46690_ (_14200_, _14198_, _14194_);
  nand _46691_ (_14201_, _14200_, _06751_);
  nor _46692_ (_14202_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  nor _46693_ (_14203_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  nor _46694_ (_14204_, _14203_, _14202_);
  nand _46695_ (_14205_, _14204_, _06717_);
  nor _46696_ (_14206_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  nor _46697_ (_14207_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nor _46698_ (_14208_, _14207_, _14206_);
  nand _46699_ (_14209_, _14208_, _06716_);
  nand _46700_ (_14210_, _14209_, _14205_);
  nand _46701_ (_14211_, _14210_, _06748_);
  nand _46702_ (_14212_, _14211_, _14201_);
  nand _46703_ (_14213_, _14212_, _06760_);
  nand _46704_ (_14214_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  nand _46705_ (_14215_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nand _46706_ (_14216_, _14215_, _14214_);
  nand _46707_ (_14217_, _14216_, _06717_);
  nand _46708_ (_14218_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nand _46709_ (_14219_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  nand _46710_ (_14221_, _14219_, _14218_);
  nand _46711_ (_14222_, _14221_, _06716_);
  nand _46712_ (_14223_, _14222_, _14217_);
  nand _46713_ (_14224_, _14223_, _06751_);
  nand _46714_ (_14225_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nand _46715_ (_14226_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nand _46716_ (_14227_, _14226_, _14225_);
  nand _46717_ (_14228_, _14227_, _06717_);
  nand _46718_ (_14229_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nand _46719_ (_14230_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  nand _46720_ (_14231_, _14230_, _14229_);
  nand _46721_ (_14232_, _14231_, _06716_);
  nand _46722_ (_14233_, _14232_, _14228_);
  nand _46723_ (_14234_, _14233_, _06748_);
  nand _46724_ (_14235_, _14234_, _14224_);
  nand _46725_ (_14236_, _14235_, _06761_);
  nand _46726_ (_14237_, _14236_, _14213_);
  nand _46727_ (_14238_, _14237_, _06731_);
  nor _46728_ (_14239_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  nor _46729_ (_14240_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  nor _46730_ (_14242_, _14240_, _14239_);
  nand _46731_ (_14243_, _14242_, _06716_);
  nand _46732_ (_14244_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  nand _46733_ (_14245_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nand _46734_ (_14246_, _14245_, _14244_);
  nand _46735_ (_14247_, _14246_, _06717_);
  nand _46736_ (_14248_, _14247_, _14243_);
  nand _46737_ (_14249_, _14248_, _06751_);
  nor _46738_ (_14250_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nor _46739_ (_14251_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  nor _46740_ (_14252_, _14251_, _14250_);
  nand _46741_ (_14253_, _14252_, _06716_);
  nand _46742_ (_14254_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nand _46743_ (_14255_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  nand _46744_ (_14256_, _14255_, _14254_);
  nand _46745_ (_14257_, _14256_, _06717_);
  nand _46746_ (_14258_, _14257_, _14253_);
  nand _46747_ (_14259_, _14258_, _06748_);
  nand _46748_ (_14260_, _14259_, _14249_);
  nand _46749_ (_14261_, _14260_, _06760_);
  nand _46750_ (_14263_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  nand _46751_ (_14264_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  nand _46752_ (_14265_, _14264_, _14263_);
  nand _46753_ (_14266_, _14265_, _06717_);
  nand _46754_ (_14267_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nand _46755_ (_14268_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  nand _46756_ (_14269_, _14268_, _14267_);
  nand _46757_ (_14270_, _14269_, _06716_);
  nand _46758_ (_14271_, _14270_, _14266_);
  nand _46759_ (_14272_, _14271_, _06751_);
  nand _46760_ (_14273_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nand _46761_ (_14274_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  nand _46762_ (_14275_, _14274_, _14273_);
  nand _46763_ (_14276_, _14275_, _06717_);
  nand _46764_ (_14277_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  nand _46765_ (_14278_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nand _46766_ (_14279_, _14278_, _14277_);
  nand _46767_ (_14280_, _14279_, _06716_);
  nand _46768_ (_14281_, _14280_, _14276_);
  nand _46769_ (_14282_, _14281_, _06748_);
  nand _46770_ (_14283_, _14282_, _14272_);
  nand _46771_ (_14284_, _14283_, _06761_);
  nand _46772_ (_14285_, _14284_, _14261_);
  nand _46773_ (_14286_, _14285_, _06780_);
  nand _46774_ (_14287_, _14286_, _14238_);
  nand _46775_ (_14288_, _14287_, _06733_);
  nand _46776_ (_14289_, _14288_, _14190_);
  nor _46777_ (_14290_, _14289_, _13106_);
  nor _46778_ (_14291_, _14290_, _14095_);
  nor _46779_ (_14292_, _14291_, _25929_);
  nand _46780_ (_14293_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nand _46781_ (_14294_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nand _46782_ (_14295_, _14294_, _14293_);
  nand _46783_ (_14296_, _14295_, _06717_);
  nand _46784_ (_14297_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  nand _46785_ (_14298_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  nand _46786_ (_14299_, _14298_, _14297_);
  nand _46787_ (_14300_, _14299_, _06716_);
  nand _46788_ (_14301_, _14300_, _14296_);
  nand _46789_ (_14302_, _14301_, _06748_);
  nand _46790_ (_14303_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nand _46791_ (_14304_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  nand _46792_ (_14305_, _14304_, _14303_);
  nand _46793_ (_14306_, _14305_, _06717_);
  nand _46794_ (_14307_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  nand _46795_ (_14308_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nand _46796_ (_14309_, _14308_, _14307_);
  nand _46797_ (_14310_, _14309_, _06716_);
  nand _46798_ (_14311_, _14310_, _14306_);
  nand _46799_ (_14312_, _14311_, _06751_);
  nand _46800_ (_14313_, _14312_, _14302_);
  nand _46801_ (_14314_, _14313_, _06761_);
  nor _46802_ (_14315_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nor _46803_ (_14316_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nor _46804_ (_14317_, _14316_, _14315_);
  nand _46805_ (_14318_, _14317_, _06717_);
  nor _46806_ (_14319_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  nor _46807_ (_14320_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  nor _46808_ (_14321_, _14320_, _14319_);
  nand _46809_ (_14322_, _14321_, _06716_);
  nand _46810_ (_14323_, _14322_, _14318_);
  nand _46811_ (_14324_, _14323_, _06748_);
  nor _46812_ (_14325_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nor _46813_ (_14326_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nor _46814_ (_14327_, _14326_, _14325_);
  nand _46815_ (_14328_, _14327_, _06717_);
  nor _46816_ (_14329_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  nor _46817_ (_14330_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  nor _46818_ (_14331_, _14330_, _14329_);
  nand _46819_ (_14332_, _14331_, _06716_);
  nand _46820_ (_14333_, _14332_, _14328_);
  nand _46821_ (_14334_, _14333_, _06751_);
  nand _46822_ (_14335_, _14334_, _14324_);
  nand _46823_ (_14336_, _14335_, _06760_);
  nand _46824_ (_14337_, _14336_, _14314_);
  nand _46825_ (_14338_, _14337_, _06731_);
  nand _46826_ (_14339_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  nand _46827_ (_14340_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  nand _46828_ (_14341_, _14340_, _14339_);
  nand _46829_ (_14342_, _14341_, _06717_);
  nand _46830_ (_14343_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  nand _46831_ (_14344_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  nand _46832_ (_14345_, _14344_, _14343_);
  nand _46833_ (_14346_, _14345_, _06716_);
  nand _46834_ (_14347_, _14346_, _14342_);
  nand _46835_ (_14348_, _14347_, _06748_);
  nand _46836_ (_14349_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  nand _46837_ (_14350_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  nand _46838_ (_14351_, _14350_, _14349_);
  nand _46839_ (_14352_, _14351_, _06717_);
  nand _46840_ (_14353_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  nand _46841_ (_14354_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  nand _46842_ (_14355_, _14354_, _14353_);
  nand _46843_ (_14356_, _14355_, _06716_);
  nand _46844_ (_14357_, _14356_, _14352_);
  nand _46845_ (_14358_, _14357_, _06751_);
  nand _46846_ (_14359_, _14358_, _14348_);
  nand _46847_ (_14360_, _14359_, _06761_);
  nor _46848_ (_14361_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  nor _46849_ (_14362_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  nor _46850_ (_14363_, _14362_, _14361_);
  nand _46851_ (_14364_, _14363_, _06716_);
  nand _46852_ (_14365_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  nand _46853_ (_14366_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  nand _46854_ (_14367_, _14366_, _14365_);
  nand _46855_ (_14368_, _14367_, _06717_);
  nand _46856_ (_14369_, _14368_, _14364_);
  nand _46857_ (_14370_, _14369_, _06748_);
  nor _46858_ (_14371_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  nor _46859_ (_14372_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  nor _46860_ (_14373_, _14372_, _14371_);
  nand _46861_ (_14374_, _14373_, _06716_);
  nand _46862_ (_14375_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  nand _46863_ (_14376_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  nand _46864_ (_14377_, _14376_, _14375_);
  nand _46865_ (_14378_, _14377_, _06717_);
  nand _46866_ (_14379_, _14378_, _14374_);
  nand _46867_ (_14380_, _14379_, _06751_);
  nand _46868_ (_14381_, _14380_, _14370_);
  nand _46869_ (_14382_, _14381_, _06760_);
  nand _46870_ (_14383_, _14382_, _14360_);
  nand _46871_ (_14384_, _14383_, _06780_);
  nand _46872_ (_14385_, _14384_, _14338_);
  nand _46873_ (_14386_, _14385_, _06734_);
  nand _46874_ (_14387_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  nand _46875_ (_14388_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nand _46876_ (_14389_, _14388_, _14387_);
  nand _46877_ (_14390_, _14389_, _06717_);
  nand _46878_ (_14391_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  nand _46879_ (_14392_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nand _46880_ (_14394_, _14392_, _14391_);
  nand _46881_ (_14395_, _14394_, _06716_);
  nand _46882_ (_14396_, _14395_, _14390_);
  nand _46883_ (_14397_, _14396_, _06748_);
  nand _46884_ (_14398_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nand _46885_ (_14399_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  nand _46886_ (_14400_, _14399_, _14398_);
  nand _46887_ (_14401_, _14400_, _06717_);
  nand _46888_ (_14402_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  nand _46889_ (_14403_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  nand _46890_ (_14404_, _14403_, _14402_);
  nand _46891_ (_14405_, _14404_, _06716_);
  nand _46892_ (_14406_, _14405_, _14401_);
  nand _46893_ (_14407_, _14406_, _06751_);
  nand _46894_ (_14408_, _14407_, _14397_);
  nand _46895_ (_14409_, _14408_, _06761_);
  nor _46896_ (_14410_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  nor _46897_ (_14411_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  nor _46898_ (_14412_, _14411_, _14410_);
  nand _46899_ (_14413_, _14412_, _06716_);
  nand _46900_ (_14414_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nand _46901_ (_14415_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nand _46902_ (_14416_, _14415_, _14414_);
  nand _46903_ (_14417_, _14416_, _06717_);
  nand _46904_ (_14418_, _14417_, _14413_);
  nand _46905_ (_14419_, _14418_, _06748_);
  nor _46906_ (_14420_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  nor _46907_ (_14421_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nor _46908_ (_14422_, _14421_, _14420_);
  nand _46909_ (_14423_, _14422_, _06716_);
  nand _46910_ (_14424_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nand _46911_ (_14425_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nand _46912_ (_14426_, _14425_, _14424_);
  nand _46913_ (_14427_, _14426_, _06717_);
  nand _46914_ (_14428_, _14427_, _14423_);
  nand _46915_ (_14429_, _14428_, _06751_);
  nand _46916_ (_14430_, _14429_, _14419_);
  nand _46917_ (_14431_, _14430_, _06760_);
  nand _46918_ (_14432_, _14431_, _14409_);
  nand _46919_ (_14433_, _14432_, _06780_);
  nand _46920_ (_14434_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  nand _46921_ (_14435_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nand _46922_ (_14436_, _14435_, _14434_);
  nand _46923_ (_14437_, _14436_, _06717_);
  nand _46924_ (_14438_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nand _46925_ (_14439_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  nand _46926_ (_14440_, _14439_, _14438_);
  nand _46927_ (_14441_, _14440_, _06716_);
  nand _46928_ (_14442_, _14441_, _14437_);
  nand _46929_ (_14443_, _14442_, _06748_);
  nand _46930_ (_14444_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  nand _46931_ (_14445_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nand _46932_ (_14446_, _14445_, _14444_);
  nand _46933_ (_14447_, _14446_, _06717_);
  nand _46934_ (_14448_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nand _46935_ (_14449_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  nand _46936_ (_14450_, _14449_, _14448_);
  nand _46937_ (_14451_, _14450_, _06716_);
  nand _46938_ (_14452_, _14451_, _14447_);
  nand _46939_ (_14453_, _14452_, _06751_);
  nand _46940_ (_14454_, _14453_, _14443_);
  nand _46941_ (_14455_, _14454_, _06761_);
  nor _46942_ (_14456_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  nor _46943_ (_14457_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nor _46944_ (_14458_, _14457_, _14456_);
  nand _46945_ (_14459_, _14458_, _06717_);
  nor _46946_ (_14460_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  nor _46947_ (_14461_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  nor _46948_ (_14462_, _14461_, _14460_);
  nand _46949_ (_14463_, _14462_, _06716_);
  nand _46950_ (_14464_, _14463_, _14459_);
  nand _46951_ (_14465_, _14464_, _06748_);
  nor _46952_ (_14466_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nor _46953_ (_14467_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nor _46954_ (_14468_, _14467_, _14466_);
  nand _46955_ (_14469_, _14468_, _06717_);
  nor _46956_ (_14470_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  nor _46957_ (_14471_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  nor _46958_ (_14472_, _14471_, _14470_);
  nand _46959_ (_14473_, _14472_, _06716_);
  nand _46960_ (_14474_, _14473_, _14469_);
  nand _46961_ (_14475_, _14474_, _06751_);
  nand _46962_ (_14476_, _14475_, _14465_);
  nand _46963_ (_14477_, _14476_, _06760_);
  nand _46964_ (_14478_, _14477_, _14455_);
  nand _46965_ (_14479_, _14478_, _06731_);
  nand _46966_ (_14480_, _14479_, _14433_);
  nand _46967_ (_14481_, _14480_, _06733_);
  nand _46968_ (_14482_, _14481_, _14386_);
  nor _46969_ (_14483_, _14482_, _06723_);
  nand _46970_ (_14484_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  nand _46971_ (_14485_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nand _46972_ (_14486_, _14485_, _14484_);
  nand _46973_ (_14487_, _14486_, _06717_);
  nand _46974_ (_14488_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  nand _46975_ (_14489_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nand _46976_ (_14490_, _14489_, _14488_);
  nand _46977_ (_14491_, _14490_, _06716_);
  nand _46978_ (_14492_, _14491_, _14487_);
  nand _46979_ (_14493_, _14492_, _06748_);
  nand _46980_ (_14494_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  nand _46981_ (_14495_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  nand _46982_ (_14496_, _14495_, _14494_);
  nand _46983_ (_14497_, _14496_, _06717_);
  nand _46984_ (_14498_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  nand _46985_ (_14499_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  nand _46986_ (_14500_, _14499_, _14498_);
  nand _46987_ (_14501_, _14500_, _06716_);
  nand _46988_ (_14502_, _14501_, _14497_);
  nand _46989_ (_14503_, _14502_, _06751_);
  nand _46990_ (_14504_, _14503_, _14493_);
  nand _46991_ (_14505_, _14504_, _06761_);
  nor _46992_ (_14506_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nor _46993_ (_14507_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nor _46994_ (_14508_, _14507_, _14506_);
  nand _46995_ (_14509_, _14508_, _06716_);
  nand _46996_ (_14510_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nand _46997_ (_14511_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  nand _46998_ (_14512_, _14511_, _14510_);
  nand _46999_ (_14513_, _14512_, _06717_);
  nand _47000_ (_14514_, _14513_, _14509_);
  nand _47001_ (_14515_, _14514_, _06748_);
  nor _47002_ (_14516_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nor _47003_ (_14517_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  nor _47004_ (_14518_, _14517_, _14516_);
  nand _47005_ (_14519_, _14518_, _06716_);
  nand _47006_ (_14520_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  nand _47007_ (_14521_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  nand _47008_ (_14522_, _14521_, _14520_);
  nand _47009_ (_14523_, _14522_, _06717_);
  nand _47010_ (_14524_, _14523_, _14519_);
  nand _47011_ (_14525_, _14524_, _06751_);
  nand _47012_ (_14526_, _14525_, _14515_);
  nand _47013_ (_14527_, _14526_, _06760_);
  nand _47014_ (_14528_, _14527_, _14505_);
  nand _47015_ (_14529_, _14528_, _06780_);
  nand _47016_ (_14530_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  nand _47017_ (_14531_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nand _47018_ (_14532_, _14531_, _14530_);
  nand _47019_ (_14533_, _14532_, _06717_);
  nand _47020_ (_14534_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  nand _47021_ (_14535_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  nand _47022_ (_14536_, _14535_, _14534_);
  nand _47023_ (_14537_, _14536_, _06716_);
  nand _47024_ (_14538_, _14537_, _14533_);
  nand _47025_ (_14539_, _14538_, _06748_);
  nand _47026_ (_14540_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nand _47027_ (_14541_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nand _47028_ (_14542_, _14541_, _14540_);
  nand _47029_ (_14543_, _14542_, _06717_);
  nand _47030_ (_14544_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  nand _47031_ (_14545_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  nand _47032_ (_14546_, _14545_, _14544_);
  nand _47033_ (_14547_, _14546_, _06716_);
  nand _47034_ (_14548_, _14547_, _14543_);
  nand _47035_ (_14549_, _14548_, _06751_);
  nand _47036_ (_14550_, _14549_, _14539_);
  nand _47037_ (_14551_, _14550_, _06761_);
  nor _47038_ (_14552_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nor _47039_ (_14553_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  nor _47040_ (_14555_, _14553_, _14552_);
  nand _47041_ (_14556_, _14555_, _06717_);
  nor _47042_ (_14557_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nor _47043_ (_14558_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nor _47044_ (_14559_, _14558_, _14557_);
  nand _47045_ (_14560_, _14559_, _06716_);
  nand _47046_ (_14561_, _14560_, _14556_);
  nand _47047_ (_14562_, _14561_, _06748_);
  nor _47048_ (_14563_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  nor _47049_ (_14564_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  nor _47050_ (_14565_, _14564_, _14563_);
  nand _47051_ (_14566_, _14565_, _06717_);
  nor _47052_ (_14567_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  nor _47053_ (_14568_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nor _47054_ (_14569_, _14568_, _14567_);
  nand _47055_ (_14570_, _14569_, _06716_);
  nand _47056_ (_14571_, _14570_, _14566_);
  nand _47057_ (_14572_, _14571_, _06751_);
  nand _47058_ (_14573_, _14572_, _14562_);
  nand _47059_ (_14574_, _14573_, _06760_);
  nand _47060_ (_14575_, _14574_, _14551_);
  nand _47061_ (_14576_, _14575_, _06731_);
  nand _47062_ (_14577_, _14576_, _14529_);
  nand _47063_ (_14578_, _14577_, _06734_);
  nor _47064_ (_14579_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  nor _47065_ (_14580_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  nor _47066_ (_14581_, _14580_, _14579_);
  nand _47067_ (_14582_, _14581_, _06717_);
  nor _47068_ (_14583_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  nor _47069_ (_14584_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  nor _47070_ (_14585_, _14584_, _14583_);
  nand _47071_ (_14586_, _14585_, _06716_);
  nand _47072_ (_14587_, _14586_, _14582_);
  nand _47073_ (_14588_, _14587_, _06751_);
  nor _47074_ (_14589_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  nor _47075_ (_14590_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  nor _47076_ (_14591_, _14590_, _14589_);
  nand _47077_ (_14592_, _14591_, _06717_);
  nor _47078_ (_14593_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  nor _47079_ (_14594_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  nor _47080_ (_14595_, _14594_, _14593_);
  nand _47081_ (_14596_, _14595_, _06716_);
  nand _47082_ (_14597_, _14596_, _14592_);
  nand _47083_ (_14598_, _14597_, _06748_);
  nand _47084_ (_14599_, _14598_, _14588_);
  nand _47085_ (_14600_, _14599_, _06760_);
  nand _47086_ (_14601_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  nand _47087_ (_14602_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  nand _47088_ (_14603_, _14602_, _14601_);
  nand _47089_ (_14604_, _14603_, _06717_);
  nand _47090_ (_14605_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  nand _47091_ (_14606_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  nand _47092_ (_14607_, _14606_, _14605_);
  nand _47093_ (_14608_, _14607_, _06716_);
  nand _47094_ (_14609_, _14608_, _14604_);
  nand _47095_ (_14610_, _14609_, _06751_);
  nand _47096_ (_14611_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  nand _47097_ (_14612_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  nand _47098_ (_14613_, _14612_, _14611_);
  nand _47099_ (_14614_, _14613_, _06717_);
  nand _47100_ (_14615_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  nand _47101_ (_14616_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  nand _47102_ (_14617_, _14616_, _14615_);
  nand _47103_ (_14618_, _14617_, _06716_);
  nand _47104_ (_14619_, _14618_, _14614_);
  nand _47105_ (_14620_, _14619_, _06748_);
  nand _47106_ (_14621_, _14620_, _14610_);
  nand _47107_ (_14622_, _14621_, _06761_);
  nand _47108_ (_14623_, _14622_, _14600_);
  nand _47109_ (_14624_, _14623_, _06731_);
  nor _47110_ (_14625_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  nor _47111_ (_14626_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nor _47112_ (_14627_, _14626_, _14625_);
  nand _47113_ (_14628_, _14627_, _06716_);
  nand _47114_ (_14629_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nand _47115_ (_14630_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nand _47116_ (_14631_, _14630_, _14629_);
  nand _47117_ (_14632_, _14631_, _06717_);
  nand _47118_ (_14633_, _14632_, _14628_);
  nand _47119_ (_14634_, _14633_, _06751_);
  nor _47120_ (_14635_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  nor _47121_ (_14636_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  nor _47122_ (_14637_, _14636_, _14635_);
  nand _47123_ (_14638_, _14637_, _06716_);
  nand _47124_ (_14639_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  nand _47125_ (_14640_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nand _47126_ (_14641_, _14640_, _14639_);
  nand _47127_ (_14642_, _14641_, _06717_);
  nand _47128_ (_14643_, _14642_, _14638_);
  nand _47129_ (_14644_, _14643_, _06748_);
  nand _47130_ (_14645_, _14644_, _14634_);
  nand _47131_ (_14646_, _14645_, _06760_);
  nand _47132_ (_14647_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  nand _47133_ (_14648_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  nand _47134_ (_14649_, _14648_, _14647_);
  nand _47135_ (_14650_, _14649_, _06717_);
  nand _47136_ (_14651_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  nand _47137_ (_14652_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nand _47138_ (_14653_, _14652_, _14651_);
  nand _47139_ (_14654_, _14653_, _06716_);
  nand _47140_ (_14655_, _14654_, _14650_);
  nand _47141_ (_14656_, _14655_, _06751_);
  nand _47142_ (_14657_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  nand _47143_ (_14658_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nand _47144_ (_14659_, _14658_, _14657_);
  nand _47145_ (_14660_, _14659_, _06717_);
  nand _47146_ (_14661_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nand _47147_ (_14662_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nand _47148_ (_14663_, _14662_, _14661_);
  nand _47149_ (_14664_, _14663_, _06716_);
  nand _47150_ (_14665_, _14664_, _14660_);
  nand _47151_ (_14666_, _14665_, _06748_);
  nand _47152_ (_14667_, _14666_, _14656_);
  nand _47153_ (_14668_, _14667_, _06761_);
  nand _47154_ (_14669_, _14668_, _14646_);
  nand _47155_ (_14670_, _14669_, _06780_);
  nand _47156_ (_14671_, _14670_, _14624_);
  nand _47157_ (_14672_, _14671_, _06733_);
  nand _47158_ (_14673_, _14672_, _14578_);
  nor _47159_ (_14674_, _14673_, _13106_);
  nor _47160_ (_14675_, _14674_, _14483_);
  nor _47161_ (_14676_, _14675_, _25843_);
  nor _47162_ (_14677_, _14676_, _14292_);
  nor _47163_ (_14678_, _14677_, _13105_);
  nand _47164_ (_14679_, _13105_, _24411_);
  nand _47165_ (_14680_, _14679_, _26487_);
  nor _47166_ (_06674_, _14680_, _14678_);
  nand _47167_ (_14681_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  nand _47168_ (_14682_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  nand _47169_ (_14683_, _14682_, _14681_);
  nand _47170_ (_14684_, _14683_, _06717_);
  nand _47171_ (_14685_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nand _47172_ (_14686_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nand _47173_ (_14687_, _14686_, _14685_);
  nand _47174_ (_14688_, _14687_, _06716_);
  nand _47175_ (_14689_, _14688_, _14684_);
  nand _47176_ (_14690_, _14689_, _06748_);
  nand _47177_ (_14691_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nand _47178_ (_14692_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  nand _47179_ (_14693_, _14692_, _14691_);
  nand _47180_ (_14694_, _14693_, _06717_);
  nand _47181_ (_14695_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  nand _47182_ (_14696_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nand _47183_ (_14697_, _14696_, _14695_);
  nand _47184_ (_14698_, _14697_, _06716_);
  nand _47185_ (_14699_, _14698_, _14694_);
  nand _47186_ (_14700_, _14699_, _06751_);
  nand _47187_ (_14701_, _14700_, _14690_);
  nand _47188_ (_14702_, _14701_, _06761_);
  nor _47189_ (_14703_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  nor _47190_ (_14704_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nor _47191_ (_14705_, _14704_, _14703_);
  nand _47192_ (_14706_, _14705_, _06716_);
  nand _47193_ (_14707_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  nand _47194_ (_14708_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  nand _47195_ (_14709_, _14708_, _14707_);
  nand _47196_ (_14710_, _14709_, _06717_);
  nand _47197_ (_14711_, _14710_, _14706_);
  nand _47198_ (_14712_, _14711_, _06748_);
  nor _47199_ (_14713_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  nor _47200_ (_14714_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nor _47201_ (_14715_, _14714_, _14713_);
  nand _47202_ (_14716_, _14715_, _06716_);
  nand _47203_ (_14717_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  nand _47204_ (_14718_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nand _47205_ (_14719_, _14718_, _14717_);
  nand _47206_ (_14720_, _14719_, _06717_);
  nand _47207_ (_14721_, _14720_, _14716_);
  nand _47208_ (_14722_, _14721_, _06751_);
  nand _47209_ (_14723_, _14722_, _14712_);
  nand _47210_ (_14724_, _14723_, _06760_);
  nand _47211_ (_14725_, _14724_, _14702_);
  nand _47212_ (_14726_, _14725_, _06780_);
  nand _47213_ (_14727_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  nand _47214_ (_14728_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nand _47215_ (_14729_, _14728_, _14727_);
  nand _47216_ (_14730_, _14729_, _06717_);
  nand _47217_ (_14731_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nand _47218_ (_14732_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  nand _47219_ (_14733_, _14732_, _14731_);
  nand _47220_ (_14734_, _14733_, _06716_);
  nand _47221_ (_14735_, _14734_, _14730_);
  nand _47222_ (_14736_, _14735_, _06748_);
  nand _47223_ (_14737_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  nand _47224_ (_14738_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  nand _47225_ (_14739_, _14738_, _14737_);
  nand _47226_ (_14740_, _14739_, _06717_);
  nand _47227_ (_14741_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nand _47228_ (_14742_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  nand _47229_ (_14743_, _14742_, _14741_);
  nand _47230_ (_14745_, _14743_, _06716_);
  nand _47231_ (_14746_, _14745_, _14740_);
  nand _47232_ (_14747_, _14746_, _06751_);
  nand _47233_ (_14748_, _14747_, _14736_);
  nand _47234_ (_14749_, _14748_, _06761_);
  nor _47235_ (_14750_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  nor _47236_ (_14751_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nor _47237_ (_14752_, _14751_, _14750_);
  nand _47238_ (_14753_, _14752_, _06717_);
  nor _47239_ (_14754_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nor _47240_ (_14755_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  nor _47241_ (_14756_, _14755_, _14754_);
  nand _47242_ (_14757_, _14756_, _06716_);
  nand _47243_ (_14758_, _14757_, _14753_);
  nand _47244_ (_14759_, _14758_, _06748_);
  nor _47245_ (_14760_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  nor _47246_ (_14761_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nor _47247_ (_14762_, _14761_, _14760_);
  nand _47248_ (_14763_, _14762_, _06717_);
  nor _47249_ (_14764_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  nor _47250_ (_14765_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  nor _47251_ (_14766_, _14765_, _14764_);
  nand _47252_ (_14767_, _14766_, _06716_);
  nand _47253_ (_14768_, _14767_, _14763_);
  nand _47254_ (_14769_, _14768_, _06751_);
  nand _47255_ (_14770_, _14769_, _14759_);
  nand _47256_ (_14771_, _14770_, _06760_);
  nand _47257_ (_14772_, _14771_, _14749_);
  nand _47258_ (_14773_, _14772_, _06731_);
  nand _47259_ (_14774_, _14773_, _14726_);
  nand _47260_ (_14776_, _14774_, _06734_);
  nand _47261_ (_14777_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand _47262_ (_14778_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nand _47263_ (_14779_, _14778_, _14777_);
  nand _47264_ (_14780_, _14779_, _06717_);
  nand _47265_ (_14781_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand _47266_ (_14782_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nand _47267_ (_14783_, _14782_, _14781_);
  nand _47268_ (_14784_, _14783_, _06716_);
  nand _47269_ (_14785_, _14784_, _14780_);
  nand _47270_ (_14786_, _14785_, _06748_);
  nand _47271_ (_14787_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand _47272_ (_14788_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nand _47273_ (_14789_, _14788_, _14787_);
  nand _47274_ (_14790_, _14789_, _06717_);
  nand _47275_ (_14791_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand _47276_ (_14792_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nand _47277_ (_14793_, _14792_, _14791_);
  nand _47278_ (_14794_, _14793_, _06716_);
  nand _47279_ (_14795_, _14794_, _14790_);
  nand _47280_ (_14796_, _14795_, _06751_);
  nand _47281_ (_14797_, _14796_, _14786_);
  nand _47282_ (_14798_, _14797_, _06761_);
  nor _47283_ (_14799_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _47284_ (_14800_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _47285_ (_14801_, _14800_, _14799_);
  nand _47286_ (_14802_, _14801_, _06716_);
  nand _47287_ (_14803_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nand _47288_ (_14804_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand _47289_ (_14805_, _14804_, _14803_);
  nand _47290_ (_14806_, _14805_, _06717_);
  nand _47291_ (_14807_, _14806_, _14802_);
  nand _47292_ (_14808_, _14807_, _06748_);
  nor _47293_ (_14809_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _47294_ (_14810_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor _47295_ (_14811_, _14810_, _14809_);
  nand _47296_ (_14812_, _14811_, _06716_);
  nand _47297_ (_14813_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nand _47298_ (_14814_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand _47299_ (_14815_, _14814_, _14813_);
  nand _47300_ (_14816_, _14815_, _06717_);
  nand _47301_ (_14817_, _14816_, _14812_);
  nand _47302_ (_14818_, _14817_, _06751_);
  nand _47303_ (_14819_, _14818_, _14808_);
  nand _47304_ (_14820_, _14819_, _06760_);
  nand _47305_ (_14821_, _14820_, _14798_);
  nand _47306_ (_14822_, _14821_, _06780_);
  nand _47307_ (_14823_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nand _47308_ (_14824_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nand _47309_ (_14825_, _14824_, _14823_);
  nand _47310_ (_14826_, _14825_, _06717_);
  nand _47311_ (_14827_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  nand _47312_ (_14828_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  nand _47313_ (_14829_, _14828_, _14827_);
  nand _47314_ (_14830_, _14829_, _06716_);
  nand _47315_ (_14831_, _14830_, _14826_);
  nand _47316_ (_14832_, _14831_, _06748_);
  nand _47317_ (_14833_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nand _47318_ (_14834_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  nand _47319_ (_14835_, _14834_, _14833_);
  nand _47320_ (_14836_, _14835_, _06717_);
  nand _47321_ (_14837_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  nand _47322_ (_14838_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nand _47323_ (_14839_, _14838_, _14837_);
  nand _47324_ (_14840_, _14839_, _06716_);
  nand _47325_ (_14841_, _14840_, _14836_);
  nand _47326_ (_14842_, _14841_, _06751_);
  nand _47327_ (_14843_, _14842_, _14832_);
  nand _47328_ (_14844_, _14843_, _06761_);
  not _47329_ (_14845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nand _47330_ (_14846_, _06774_, _14845_);
  nor _47331_ (_14847_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nor _47332_ (_14848_, _14847_, _06716_);
  nand _47333_ (_14849_, _14848_, _14846_);
  nor _47334_ (_14850_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  nor _47335_ (_14851_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  nor _47336_ (_14852_, _14851_, _14850_);
  nand _47337_ (_14853_, _14852_, _06716_);
  nand _47338_ (_14854_, _14853_, _14849_);
  nand _47339_ (_14855_, _14854_, _06748_);
  nor _47340_ (_14856_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nor _47341_ (_14857_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  nor _47342_ (_14858_, _14857_, _14856_);
  nand _47343_ (_14859_, _14858_, _06717_);
  nor _47344_ (_14860_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nor _47345_ (_14861_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nor _47346_ (_14862_, _14861_, _14860_);
  nand _47347_ (_14863_, _14862_, _06716_);
  nand _47348_ (_14864_, _14863_, _14859_);
  nand _47349_ (_14865_, _14864_, _06751_);
  nand _47350_ (_14866_, _14865_, _14855_);
  nand _47351_ (_14867_, _14866_, _06760_);
  nand _47352_ (_14868_, _14867_, _14844_);
  nand _47353_ (_14869_, _14868_, _06731_);
  nand _47354_ (_14870_, _14869_, _14822_);
  nand _47355_ (_14871_, _14870_, _06733_);
  nand _47356_ (_14872_, _14871_, _14776_);
  nor _47357_ (_14873_, _14872_, _06723_);
  nand _47358_ (_14874_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nand _47359_ (_14875_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  nand _47360_ (_14876_, _14875_, _14874_);
  nand _47361_ (_14877_, _14876_, _06717_);
  nand _47362_ (_14878_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  nand _47363_ (_14879_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nand _47364_ (_14880_, _14879_, _14878_);
  nand _47365_ (_14881_, _14880_, _06716_);
  nand _47366_ (_14882_, _14881_, _14877_);
  nand _47367_ (_14883_, _14882_, _06748_);
  nand _47368_ (_14884_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nand _47369_ (_14885_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  nand _47370_ (_14886_, _14885_, _14884_);
  nand _47371_ (_14887_, _14886_, _06717_);
  nand _47372_ (_14888_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  nand _47373_ (_14889_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nand _47374_ (_14890_, _14889_, _14888_);
  nand _47375_ (_14891_, _14890_, _06716_);
  nand _47376_ (_14892_, _14891_, _14887_);
  nand _47377_ (_14893_, _14892_, _06751_);
  nand _47378_ (_14894_, _14893_, _14883_);
  nand _47379_ (_14895_, _14894_, _06761_);
  nor _47380_ (_14896_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nor _47381_ (_14897_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  nor _47382_ (_14898_, _14897_, _14896_);
  nand _47383_ (_14899_, _14898_, _06717_);
  nor _47384_ (_14900_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nor _47385_ (_14901_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nor _47386_ (_14902_, _14901_, _14900_);
  nand _47387_ (_14903_, _14902_, _06716_);
  nand _47388_ (_14904_, _14903_, _14899_);
  nand _47389_ (_14905_, _14904_, _06748_);
  not _47390_ (_14906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nand _47391_ (_14907_, _06774_, _14906_);
  nor _47392_ (_14908_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  nor _47393_ (_14909_, _14908_, _06716_);
  nand _47394_ (_14910_, _14909_, _14907_);
  nor _47395_ (_14911_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nor _47396_ (_14912_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  nor _47397_ (_14913_, _14912_, _14911_);
  nand _47398_ (_14914_, _14913_, _06716_);
  nand _47399_ (_14915_, _14914_, _14910_);
  nand _47400_ (_14916_, _14915_, _06751_);
  nand _47401_ (_14917_, _14916_, _14905_);
  nand _47402_ (_14918_, _14917_, _06760_);
  nand _47403_ (_14919_, _14918_, _14895_);
  nand _47404_ (_14920_, _14919_, _06780_);
  nand _47405_ (_14921_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  nand _47406_ (_14922_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  nand _47407_ (_14923_, _14922_, _14921_);
  nand _47408_ (_14924_, _14923_, _06717_);
  nand _47409_ (_14925_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nand _47410_ (_14927_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nand _47411_ (_14928_, _14927_, _14925_);
  nand _47412_ (_14929_, _14928_, _06716_);
  nand _47413_ (_14930_, _14929_, _14924_);
  nand _47414_ (_14931_, _14930_, _06748_);
  nand _47415_ (_14932_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  nand _47416_ (_14933_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  nand _47417_ (_14934_, _14933_, _14932_);
  nand _47418_ (_14935_, _14934_, _06717_);
  nand _47419_ (_14936_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nand _47420_ (_14937_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nand _47421_ (_14938_, _14937_, _14936_);
  nand _47422_ (_14939_, _14938_, _06716_);
  nand _47423_ (_14940_, _14939_, _14935_);
  nand _47424_ (_14941_, _14940_, _06751_);
  nand _47425_ (_14942_, _14941_, _14931_);
  nand _47426_ (_14943_, _14942_, _06761_);
  not _47427_ (_14944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  nand _47428_ (_14945_, _06774_, _14944_);
  nor _47429_ (_14946_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  nor _47430_ (_14947_, _14946_, _06716_);
  nand _47431_ (_14948_, _14947_, _14945_);
  nor _47432_ (_14949_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  nor _47433_ (_14950_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nor _47434_ (_14951_, _14950_, _14949_);
  nand _47435_ (_14952_, _14951_, _06716_);
  nand _47436_ (_14953_, _14952_, _14948_);
  nand _47437_ (_14954_, _14953_, _06748_);
  nor _47438_ (_14955_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nor _47439_ (_14956_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  nor _47440_ (_14957_, _14956_, _14955_);
  nand _47441_ (_14958_, _14957_, _06717_);
  nor _47442_ (_14959_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  nor _47443_ (_14960_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nor _47444_ (_14961_, _14960_, _14959_);
  nand _47445_ (_14962_, _14961_, _06716_);
  nand _47446_ (_14963_, _14962_, _14958_);
  nand _47447_ (_14964_, _14963_, _06751_);
  nand _47448_ (_14965_, _14964_, _14954_);
  nand _47449_ (_14966_, _14965_, _06760_);
  nand _47450_ (_14967_, _14966_, _14943_);
  nand _47451_ (_14968_, _14967_, _06731_);
  nand _47452_ (_14969_, _14968_, _14920_);
  nand _47453_ (_14970_, _14969_, _06733_);
  nand _47454_ (_14971_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  nand _47455_ (_14972_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  nand _47456_ (_14973_, _14972_, _14971_);
  nand _47457_ (_14974_, _14973_, _06716_);
  nand _47458_ (_14975_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nand _47459_ (_14976_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  nand _47460_ (_14977_, _14976_, _14975_);
  nand _47461_ (_14978_, _14977_, _06717_);
  nand _47462_ (_14979_, _14978_, _14974_);
  nand _47463_ (_14980_, _14979_, _06748_);
  nand _47464_ (_14981_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  nand _47465_ (_14982_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  nand _47466_ (_14983_, _14982_, _14981_);
  nand _47467_ (_14984_, _14983_, _06716_);
  nand _47468_ (_14985_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nand _47469_ (_14986_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  nand _47470_ (_14988_, _14986_, _14985_);
  nand _47471_ (_14989_, _14988_, _06717_);
  nand _47472_ (_14990_, _14989_, _14984_);
  nand _47473_ (_14991_, _14990_, _06751_);
  nand _47474_ (_14992_, _14991_, _14980_);
  nand _47475_ (_14993_, _14992_, _06761_);
  nand _47476_ (_14994_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  nand _47477_ (_14995_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  nand _47478_ (_14996_, _14995_, _14994_);
  nand _47479_ (_14997_, _14996_, _06717_);
  nor _47480_ (_14998_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nor _47481_ (_14999_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  nor _47482_ (_15000_, _14999_, _14998_);
  nand _47483_ (_15001_, _15000_, _06716_);
  nand _47484_ (_15002_, _15001_, _14997_);
  nand _47485_ (_15003_, _15002_, _06748_);
  nand _47486_ (_15004_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nand _47487_ (_15005_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nand _47488_ (_15006_, _15005_, _15004_);
  nand _47489_ (_15007_, _15006_, _06717_);
  nor _47490_ (_15008_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  nor _47491_ (_15009_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nor _47492_ (_15010_, _15009_, _15008_);
  nand _47493_ (_15011_, _15010_, _06716_);
  nand _47494_ (_15012_, _15011_, _15007_);
  nand _47495_ (_15013_, _15012_, _06751_);
  nand _47496_ (_15014_, _15013_, _15003_);
  nand _47497_ (_15015_, _15014_, _06760_);
  nand _47498_ (_15016_, _15015_, _14993_);
  nand _47499_ (_15017_, _15016_, _06780_);
  nand _47500_ (_15018_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  nand _47501_ (_15019_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  nand _47502_ (_15020_, _15019_, _15018_);
  nand _47503_ (_15021_, _15020_, _06717_);
  nand _47504_ (_15022_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  nand _47505_ (_15023_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nand _47506_ (_15024_, _15023_, _15022_);
  nand _47507_ (_15025_, _15024_, _06716_);
  nand _47508_ (_15026_, _15025_, _15021_);
  nand _47509_ (_15027_, _15026_, _06748_);
  nand _47510_ (_15028_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nand _47511_ (_15029_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nand _47512_ (_15030_, _15029_, _15028_);
  nand _47513_ (_15031_, _15030_, _06717_);
  nand _47514_ (_15032_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  nand _47515_ (_15033_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  nand _47516_ (_15034_, _15033_, _15032_);
  nand _47517_ (_15035_, _15034_, _06716_);
  nand _47518_ (_15036_, _15035_, _15031_);
  nand _47519_ (_15037_, _15036_, _06751_);
  nand _47520_ (_15038_, _15037_, _15027_);
  nand _47521_ (_15039_, _15038_, _06761_);
  nor _47522_ (_15040_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  nor _47523_ (_15041_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nor _47524_ (_15042_, _15041_, _15040_);
  nand _47525_ (_15043_, _15042_, _06717_);
  nor _47526_ (_15044_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  nor _47527_ (_15045_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  nor _47528_ (_15046_, _15045_, _15044_);
  nand _47529_ (_15047_, _15046_, _06716_);
  nand _47530_ (_15048_, _15047_, _15043_);
  nand _47531_ (_15049_, _15048_, _06748_);
  nor _47532_ (_15050_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nor _47533_ (_15051_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nor _47534_ (_15052_, _15051_, _15050_);
  nor _47535_ (_15053_, _15052_, _06716_);
  nor _47536_ (_15054_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nor _47537_ (_15055_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  nor _47538_ (_15056_, _15055_, _15054_);
  nor _47539_ (_15057_, _15056_, _06717_);
  nor _47540_ (_15058_, _15057_, _15053_);
  nand _47541_ (_15059_, _15058_, _06751_);
  nand _47542_ (_15060_, _15059_, _15049_);
  nand _47543_ (_15061_, _15060_, _06760_);
  nand _47544_ (_15062_, _15061_, _15039_);
  nand _47545_ (_15063_, _15062_, _06731_);
  nand _47546_ (_15064_, _15063_, _15017_);
  nand _47547_ (_15065_, _15064_, _06734_);
  nand _47548_ (_15066_, _15065_, _14970_);
  nor _47549_ (_15067_, _15066_, _13106_);
  nor _47550_ (_15068_, _15067_, _14873_);
  nor _47551_ (_15069_, _15068_, _25929_);
  nand _47552_ (_15070_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  nand _47553_ (_15071_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  nand _47554_ (_15072_, _15071_, _15070_);
  nand _47555_ (_15073_, _15072_, _06717_);
  nand _47556_ (_15074_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nand _47557_ (_15075_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nand _47558_ (_15076_, _15075_, _15074_);
  nand _47559_ (_15077_, _15076_, _06716_);
  nand _47560_ (_15078_, _15077_, _15073_);
  nand _47561_ (_15079_, _15078_, _06748_);
  nand _47562_ (_15080_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  nand _47563_ (_15081_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nand _47564_ (_15082_, _15081_, _15080_);
  nand _47565_ (_15083_, _15082_, _06717_);
  nand _47566_ (_15084_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nand _47567_ (_15085_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  nand _47568_ (_15086_, _15085_, _15084_);
  nand _47569_ (_15087_, _15086_, _06716_);
  nand _47570_ (_15088_, _15087_, _15083_);
  nand _47571_ (_15089_, _15088_, _06751_);
  nand _47572_ (_15090_, _15089_, _15079_);
  nand _47573_ (_15091_, _15090_, _06761_);
  nor _47574_ (_15092_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  nor _47575_ (_15093_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  nor _47576_ (_15094_, _15093_, _15092_);
  nand _47577_ (_15095_, _15094_, _06717_);
  nor _47578_ (_15096_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  nor _47579_ (_15097_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nor _47580_ (_15099_, _15097_, _15096_);
  nand _47581_ (_15100_, _15099_, _06716_);
  nand _47582_ (_15101_, _15100_, _15095_);
  nand _47583_ (_15102_, _15101_, _06748_);
  nor _47584_ (_15103_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nor _47585_ (_15104_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  nor _47586_ (_15105_, _15104_, _15103_);
  nand _47587_ (_15106_, _15105_, _06717_);
  nor _47588_ (_15107_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nor _47589_ (_15108_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  nor _47590_ (_15109_, _15108_, _15107_);
  nand _47591_ (_15110_, _15109_, _06716_);
  nand _47592_ (_15111_, _15110_, _15106_);
  nand _47593_ (_15112_, _15111_, _06751_);
  nand _47594_ (_15113_, _15112_, _15102_);
  nand _47595_ (_15114_, _15113_, _06760_);
  nand _47596_ (_15115_, _15114_, _15091_);
  nand _47597_ (_15116_, _15115_, _06731_);
  nand _47598_ (_15117_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nand _47599_ (_15118_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nand _47600_ (_15119_, _15118_, _15117_);
  nand _47601_ (_15120_, _15119_, _06717_);
  nand _47602_ (_15121_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  nand _47603_ (_15122_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  nand _47604_ (_15123_, _15122_, _15121_);
  nand _47605_ (_15124_, _15123_, _06716_);
  nand _47606_ (_15125_, _15124_, _15120_);
  nand _47607_ (_15126_, _15125_, _06748_);
  nand _47608_ (_15127_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  nand _47609_ (_15128_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nand _47610_ (_15129_, _15128_, _15127_);
  nand _47611_ (_15130_, _15129_, _06717_);
  nand _47612_ (_15131_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nand _47613_ (_15132_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nand _47614_ (_15133_, _15132_, _15131_);
  nand _47615_ (_15134_, _15133_, _06716_);
  nand _47616_ (_15135_, _15134_, _15130_);
  nand _47617_ (_15136_, _15135_, _06751_);
  nand _47618_ (_15137_, _15136_, _15126_);
  nand _47619_ (_15138_, _15137_, _06761_);
  nor _47620_ (_15139_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  nor _47621_ (_15140_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  nor _47622_ (_15141_, _15140_, _15139_);
  nand _47623_ (_15142_, _15141_, _06716_);
  nand _47624_ (_15143_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  nand _47625_ (_15144_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nand _47626_ (_15145_, _15144_, _15143_);
  nand _47627_ (_15146_, _15145_, _06717_);
  nand _47628_ (_15147_, _15146_, _15142_);
  nand _47629_ (_15148_, _15147_, _06748_);
  nor _47630_ (_15149_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nor _47631_ (_15150_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nor _47632_ (_15151_, _15150_, _15149_);
  nand _47633_ (_15152_, _15151_, _06716_);
  nand _47634_ (_15153_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nand _47635_ (_15154_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  nand _47636_ (_15155_, _15154_, _15153_);
  nand _47637_ (_15156_, _15155_, _06717_);
  nand _47638_ (_15157_, _15156_, _15152_);
  nand _47639_ (_15158_, _15157_, _06751_);
  nand _47640_ (_15159_, _15158_, _15148_);
  nand _47641_ (_15160_, _15159_, _06760_);
  nand _47642_ (_15161_, _15160_, _15138_);
  nand _47643_ (_15162_, _15161_, _06780_);
  nand _47644_ (_15163_, _15162_, _15116_);
  nand _47645_ (_15164_, _15163_, _06734_);
  nand _47646_ (_15165_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nand _47647_ (_15166_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  nand _47648_ (_15167_, _15166_, _15165_);
  nand _47649_ (_15168_, _15167_, _06717_);
  nand _47650_ (_15169_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  nand _47651_ (_15170_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nand _47652_ (_15171_, _15170_, _15169_);
  nand _47653_ (_15172_, _15171_, _06716_);
  nand _47654_ (_15173_, _15172_, _15168_);
  nand _47655_ (_15174_, _15173_, _06748_);
  nand _47656_ (_15175_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  nand _47657_ (_15176_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  nand _47658_ (_15177_, _15176_, _15175_);
  nand _47659_ (_15178_, _15177_, _06717_);
  nand _47660_ (_15179_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nand _47661_ (_15180_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  nand _47662_ (_15181_, _15180_, _15179_);
  nand _47663_ (_15182_, _15181_, _06716_);
  nand _47664_ (_15183_, _15182_, _15178_);
  nand _47665_ (_15184_, _15183_, _06751_);
  nand _47666_ (_15185_, _15184_, _15174_);
  nand _47667_ (_15186_, _15185_, _06761_);
  nor _47668_ (_15187_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  nor _47669_ (_15188_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nor _47670_ (_15189_, _15188_, _15187_);
  nand _47671_ (_15190_, _15189_, _06716_);
  nand _47672_ (_15191_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nand _47673_ (_15192_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nand _47674_ (_15193_, _15192_, _15191_);
  nand _47675_ (_15194_, _15193_, _06717_);
  nand _47676_ (_15195_, _15194_, _15190_);
  nand _47677_ (_15196_, _15195_, _06748_);
  nor _47678_ (_15197_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  nor _47679_ (_15198_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nor _47680_ (_15199_, _15198_, _15197_);
  nand _47681_ (_15200_, _15199_, _06716_);
  nand _47682_ (_15201_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  nand _47683_ (_15202_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  nand _47684_ (_15203_, _15202_, _15201_);
  nand _47685_ (_15204_, _15203_, _06717_);
  nand _47686_ (_15205_, _15204_, _15200_);
  nand _47687_ (_15206_, _15205_, _06751_);
  nand _47688_ (_15207_, _15206_, _15196_);
  nand _47689_ (_15208_, _15207_, _06760_);
  nand _47690_ (_15209_, _15208_, _15186_);
  nand _47691_ (_15210_, _15209_, _06780_);
  nand _47692_ (_15211_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  nand _47693_ (_15212_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nand _47694_ (_15213_, _15212_, _15211_);
  nand _47695_ (_15214_, _15213_, _06717_);
  nand _47696_ (_15215_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  nand _47697_ (_15216_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  nand _47698_ (_15217_, _15216_, _15215_);
  nand _47699_ (_15218_, _15217_, _06716_);
  nand _47700_ (_15219_, _15218_, _15214_);
  nand _47701_ (_15220_, _15219_, _06748_);
  nand _47702_ (_15221_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  nand _47703_ (_15222_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  nand _47704_ (_15223_, _15222_, _15221_);
  nand _47705_ (_15224_, _15223_, _06717_);
  nand _47706_ (_15225_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nand _47707_ (_15226_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nand _47708_ (_15227_, _15226_, _15225_);
  nand _47709_ (_15228_, _15227_, _06716_);
  nand _47710_ (_15229_, _15228_, _15224_);
  nand _47711_ (_15230_, _15229_, _06751_);
  nand _47712_ (_15231_, _15230_, _15220_);
  nand _47713_ (_15232_, _15231_, _06761_);
  nor _47714_ (_15233_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  nor _47715_ (_15234_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nor _47716_ (_15235_, _15234_, _15233_);
  nand _47717_ (_15236_, _15235_, _06717_);
  nor _47718_ (_15237_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nor _47719_ (_15238_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  nor _47720_ (_15239_, _15238_, _15237_);
  nand _47721_ (_15240_, _15239_, _06716_);
  nand _47722_ (_15241_, _15240_, _15236_);
  nand _47723_ (_15242_, _15241_, _06748_);
  nor _47724_ (_15243_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  nor _47725_ (_15244_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  nor _47726_ (_15245_, _15244_, _15243_);
  nand _47727_ (_15246_, _15245_, _06717_);
  nor _47728_ (_15247_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  nor _47729_ (_15248_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nor _47730_ (_15249_, _15248_, _15247_);
  nand _47731_ (_15250_, _15249_, _06716_);
  nand _47732_ (_15251_, _15250_, _15246_);
  nand _47733_ (_15252_, _15251_, _06751_);
  nand _47734_ (_15253_, _15252_, _15242_);
  nand _47735_ (_15254_, _15253_, _06760_);
  nand _47736_ (_15255_, _15254_, _15232_);
  nand _47737_ (_15256_, _15255_, _06731_);
  nand _47738_ (_15257_, _15256_, _15210_);
  nand _47739_ (_15258_, _15257_, _06733_);
  nand _47740_ (_15259_, _15258_, _15164_);
  nor _47741_ (_15260_, _15259_, _06723_);
  nand _47742_ (_15261_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nand _47743_ (_15262_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nand _47744_ (_15263_, _15262_, _15261_);
  nand _47745_ (_15264_, _15263_, _06717_);
  nand _47746_ (_15265_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  nand _47747_ (_15266_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nand _47748_ (_15267_, _15266_, _15265_);
  nand _47749_ (_15268_, _15267_, _06716_);
  nand _47750_ (_15269_, _15268_, _15264_);
  nand _47751_ (_15270_, _15269_, _06748_);
  nand _47752_ (_15271_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  nand _47753_ (_15272_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  nand _47754_ (_15273_, _15272_, _15271_);
  nand _47755_ (_15274_, _15273_, _06717_);
  nand _47756_ (_15275_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  nand _47757_ (_15276_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nand _47758_ (_15277_, _15276_, _15275_);
  nand _47759_ (_15278_, _15277_, _06716_);
  nand _47760_ (_15279_, _15278_, _15274_);
  nand _47761_ (_15280_, _15279_, _06751_);
  nand _47762_ (_15281_, _15280_, _15270_);
  nand _47763_ (_15282_, _15281_, _06761_);
  nor _47764_ (_15283_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  nor _47765_ (_15284_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  nor _47766_ (_15285_, _15284_, _15283_);
  nand _47767_ (_15286_, _15285_, _06716_);
  nand _47768_ (_15287_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  nand _47769_ (_15288_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nand _47770_ (_15289_, _15288_, _15287_);
  nand _47771_ (_15290_, _15289_, _06717_);
  nand _47772_ (_15291_, _15290_, _15286_);
  nand _47773_ (_15292_, _15291_, _06748_);
  nor _47774_ (_15293_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  nor _47775_ (_15294_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  nor _47776_ (_15295_, _15294_, _15293_);
  nand _47777_ (_15296_, _15295_, _06716_);
  nand _47778_ (_15297_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nand _47779_ (_15298_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nand _47780_ (_15299_, _15298_, _15297_);
  nand _47781_ (_15300_, _15299_, _06717_);
  nand _47782_ (_15301_, _15300_, _15296_);
  nand _47783_ (_15302_, _15301_, _06751_);
  nand _47784_ (_15303_, _15302_, _15292_);
  nand _47785_ (_15304_, _15303_, _06760_);
  nand _47786_ (_15305_, _15304_, _15282_);
  nand _47787_ (_15306_, _15305_, _06780_);
  nand _47788_ (_15307_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nand _47789_ (_15308_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nand _47790_ (_15310_, _15308_, _15307_);
  nand _47791_ (_15311_, _15310_, _06717_);
  nand _47792_ (_15312_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  nand _47793_ (_15313_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  nand _47794_ (_15314_, _15313_, _15312_);
  nand _47795_ (_15315_, _15314_, _06716_);
  nand _47796_ (_15316_, _15315_, _15311_);
  nand _47797_ (_15317_, _15316_, _06748_);
  nand _47798_ (_15318_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nand _47799_ (_15319_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  nand _47800_ (_15320_, _15319_, _15318_);
  nand _47801_ (_15321_, _15320_, _06717_);
  nand _47802_ (_15322_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nand _47803_ (_15323_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nand _47804_ (_15324_, _15323_, _15322_);
  nand _47805_ (_15325_, _15324_, _06716_);
  nand _47806_ (_15326_, _15325_, _15321_);
  nand _47807_ (_15327_, _15326_, _06751_);
  nand _47808_ (_15328_, _15327_, _15317_);
  nand _47809_ (_15329_, _15328_, _06761_);
  nor _47810_ (_15330_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  nor _47811_ (_15331_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  nor _47812_ (_15332_, _15331_, _15330_);
  nand _47813_ (_15333_, _15332_, _06717_);
  nor _47814_ (_15334_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  nor _47815_ (_15335_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nor _47816_ (_15336_, _15335_, _15334_);
  nand _47817_ (_15337_, _15336_, _06716_);
  nand _47818_ (_15338_, _15337_, _15333_);
  nand _47819_ (_15339_, _15338_, _06748_);
  nor _47820_ (_15341_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nor _47821_ (_15342_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nor _47822_ (_15343_, _15342_, _15341_);
  nand _47823_ (_15344_, _15343_, _06717_);
  nor _47824_ (_15345_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  nor _47825_ (_15346_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  nor _47826_ (_15347_, _15346_, _15345_);
  nand _47827_ (_15348_, _15347_, _06716_);
  nand _47828_ (_15349_, _15348_, _15344_);
  nand _47829_ (_15350_, _15349_, _06751_);
  nand _47830_ (_15351_, _15350_, _15339_);
  nand _47831_ (_15352_, _15351_, _06760_);
  nand _47832_ (_15353_, _15352_, _15329_);
  nand _47833_ (_15354_, _15353_, _06731_);
  nand _47834_ (_15355_, _15354_, _15306_);
  nand _47835_ (_15356_, _15355_, _06734_);
  nor _47836_ (_15357_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  nor _47837_ (_15358_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nor _47838_ (_15359_, _15358_, _15357_);
  nand _47839_ (_15360_, _15359_, _06717_);
  nor _47840_ (_15362_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  nor _47841_ (_15363_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  nor _47842_ (_15364_, _15363_, _15362_);
  nand _47843_ (_15365_, _15364_, _06716_);
  nand _47844_ (_15366_, _15365_, _15360_);
  nand _47845_ (_15367_, _15366_, _06751_);
  nor _47846_ (_15368_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  nor _47847_ (_15369_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  nor _47848_ (_15370_, _15369_, _15368_);
  nand _47849_ (_15371_, _15370_, _06717_);
  nor _47850_ (_15372_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nor _47851_ (_15373_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nor _47852_ (_15374_, _15373_, _15372_);
  nand _47853_ (_15375_, _15374_, _06716_);
  nand _47854_ (_15376_, _15375_, _15371_);
  nand _47855_ (_15377_, _15376_, _06748_);
  nand _47856_ (_15378_, _15377_, _15367_);
  nand _47857_ (_15379_, _15378_, _06760_);
  nand _47858_ (_15380_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  nand _47859_ (_15381_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  nand _47860_ (_15383_, _15381_, _15380_);
  nand _47861_ (_15384_, _15383_, _06717_);
  nand _47862_ (_15385_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nand _47863_ (_15386_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nand _47864_ (_15387_, _15386_, _15385_);
  nand _47865_ (_15388_, _15387_, _06716_);
  nand _47866_ (_15389_, _15388_, _15384_);
  nand _47867_ (_15390_, _15389_, _06751_);
  nand _47868_ (_15391_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nand _47869_ (_15392_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  nand _47870_ (_15393_, _15392_, _15391_);
  nand _47871_ (_15394_, _15393_, _06717_);
  nand _47872_ (_15395_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nand _47873_ (_15396_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nand _47874_ (_15397_, _15396_, _15395_);
  nand _47875_ (_15398_, _15397_, _06716_);
  nand _47876_ (_15399_, _15398_, _15394_);
  nand _47877_ (_15400_, _15399_, _06748_);
  nand _47878_ (_15401_, _15400_, _15390_);
  nand _47879_ (_15402_, _15401_, _06761_);
  nand _47880_ (_15404_, _15402_, _15379_);
  nand _47881_ (_15405_, _15404_, _06731_);
  nor _47882_ (_15406_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  nor _47883_ (_15407_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  nor _47884_ (_15408_, _15407_, _15406_);
  nand _47885_ (_15409_, _15408_, _06716_);
  nand _47886_ (_15410_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  nand _47887_ (_15411_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nand _47888_ (_15412_, _15411_, _15410_);
  nand _47889_ (_15413_, _15412_, _06717_);
  nand _47890_ (_15414_, _15413_, _15409_);
  nand _47891_ (_15415_, _15414_, _06751_);
  nor _47892_ (_15416_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nor _47893_ (_15417_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nor _47894_ (_15418_, _15417_, _15416_);
  nand _47895_ (_15419_, _15418_, _06716_);
  nand _47896_ (_15420_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nand _47897_ (_15421_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  nand _47898_ (_15422_, _15421_, _15420_);
  nand _47899_ (_15423_, _15422_, _06717_);
  nand _47900_ (_15424_, _15423_, _15419_);
  nand _47901_ (_15425_, _15424_, _06748_);
  nand _47902_ (_15426_, _15425_, _15415_);
  nand _47903_ (_15427_, _15426_, _06760_);
  nand _47904_ (_15428_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  nand _47905_ (_15429_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  nand _47906_ (_15430_, _15429_, _15428_);
  nand _47907_ (_15431_, _15430_, _06717_);
  nand _47908_ (_15432_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nand _47909_ (_15433_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  nand _47910_ (_15434_, _15433_, _15432_);
  nand _47911_ (_15435_, _15434_, _06716_);
  nand _47912_ (_15436_, _15435_, _15431_);
  nand _47913_ (_15437_, _15436_, _06751_);
  nand _47914_ (_15438_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nand _47915_ (_15439_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  nand _47916_ (_15440_, _15439_, _15438_);
  nand _47917_ (_15441_, _15440_, _06717_);
  nand _47918_ (_15442_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  nand _47919_ (_15443_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nand _47920_ (_15444_, _15443_, _15442_);
  nand _47921_ (_15445_, _15444_, _06716_);
  nand _47922_ (_15446_, _15445_, _15441_);
  nand _47923_ (_15447_, _15446_, _06748_);
  nand _47924_ (_15448_, _15447_, _15437_);
  nand _47925_ (_15449_, _15448_, _06761_);
  nand _47926_ (_15450_, _15449_, _15427_);
  nand _47927_ (_15451_, _15450_, _06780_);
  nand _47928_ (_15452_, _15451_, _15405_);
  nand _47929_ (_15453_, _15452_, _06733_);
  nand _47930_ (_15455_, _15453_, _15356_);
  nor _47931_ (_15456_, _15455_, _13106_);
  nor _47932_ (_15457_, _15456_, _15260_);
  nor _47933_ (_15458_, _15457_, _25843_);
  nor _47934_ (_15459_, _15458_, _15069_);
  nor _47935_ (_15460_, _15459_, _13105_);
  nand _47936_ (_15461_, _13105_, _24382_);
  nand _47937_ (_15462_, _15461_, _26487_);
  nor _47938_ (_06676_, _15462_, _15460_);
  nand _47939_ (_15463_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nand _47940_ (_15464_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nand _47941_ (_15465_, _15464_, _15463_);
  nand _47942_ (_15466_, _15465_, _06717_);
  nand _47943_ (_15467_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  nand _47944_ (_15468_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  nand _47945_ (_15469_, _15468_, _15467_);
  nand _47946_ (_15470_, _15469_, _06716_);
  nand _47947_ (_15471_, _15470_, _15466_);
  nand _47948_ (_15472_, _15471_, _06748_);
  nand _47949_ (_15473_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nand _47950_ (_15474_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  nand _47951_ (_15475_, _15474_, _15473_);
  nand _47952_ (_15476_, _15475_, _06717_);
  nand _47953_ (_15477_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  nand _47954_ (_15478_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nand _47955_ (_15479_, _15478_, _15477_);
  nand _47956_ (_15480_, _15479_, _06716_);
  nand _47957_ (_15481_, _15480_, _15476_);
  nand _47958_ (_15482_, _15481_, _06751_);
  nand _47959_ (_15483_, _15482_, _15472_);
  nand _47960_ (_15484_, _15483_, _06761_);
  nor _47961_ (_15485_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  nor _47962_ (_15486_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  nor _47963_ (_15487_, _15486_, _15485_);
  nand _47964_ (_15488_, _15487_, _06717_);
  nor _47965_ (_15489_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  nor _47966_ (_15490_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  nor _47967_ (_15491_, _15490_, _15489_);
  nand _47968_ (_15492_, _15491_, _06716_);
  nand _47969_ (_15493_, _15492_, _15488_);
  nand _47970_ (_15494_, _15493_, _06748_);
  nor _47971_ (_15495_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nor _47972_ (_15496_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nor _47973_ (_15497_, _15496_, _15495_);
  nand _47974_ (_15498_, _15497_, _06717_);
  nor _47975_ (_15499_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nor _47976_ (_15500_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  nor _47977_ (_15501_, _15500_, _15499_);
  nand _47978_ (_15502_, _15501_, _06716_);
  nand _47979_ (_15503_, _15502_, _15498_);
  nand _47980_ (_15504_, _15503_, _06751_);
  nand _47981_ (_15505_, _15504_, _15494_);
  nand _47982_ (_15506_, _15505_, _06760_);
  nand _47983_ (_15507_, _15506_, _15484_);
  nand _47984_ (_15508_, _15507_, _06731_);
  nand _47985_ (_15509_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nand _47986_ (_15510_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  nand _47987_ (_15511_, _15510_, _15509_);
  nand _47988_ (_15512_, _15511_, _06717_);
  nand _47989_ (_15513_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  nand _47990_ (_15514_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nand _47991_ (_15515_, _15514_, _15513_);
  nand _47992_ (_15516_, _15515_, _06716_);
  nand _47993_ (_15517_, _15516_, _15512_);
  nand _47994_ (_15518_, _15517_, _06748_);
  nand _47995_ (_15519_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  nand _47996_ (_15520_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  nand _47997_ (_15521_, _15520_, _15519_);
  nand _47998_ (_15522_, _15521_, _06717_);
  nand _47999_ (_15523_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nand _48000_ (_15525_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  nand _48001_ (_15526_, _15525_, _15523_);
  nand _48002_ (_15527_, _15526_, _06716_);
  nand _48003_ (_15528_, _15527_, _15522_);
  nand _48004_ (_15529_, _15528_, _06751_);
  nand _48005_ (_15530_, _15529_, _15518_);
  nand _48006_ (_15531_, _15530_, _06761_);
  nor _48007_ (_15532_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nor _48008_ (_15533_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nor _48009_ (_15534_, _15533_, _15532_);
  nand _48010_ (_15535_, _15534_, _06716_);
  nand _48011_ (_15536_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nand _48012_ (_15537_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  nand _48013_ (_15538_, _15537_, _15536_);
  nand _48014_ (_15539_, _15538_, _06717_);
  nand _48015_ (_15540_, _15539_, _15535_);
  nand _48016_ (_15541_, _15540_, _06748_);
  nor _48017_ (_15542_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  nor _48018_ (_15543_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  nor _48019_ (_15544_, _15543_, _15542_);
  nand _48020_ (_15546_, _15544_, _06716_);
  nand _48021_ (_15547_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  nand _48022_ (_15548_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nand _48023_ (_15549_, _15548_, _15547_);
  nand _48024_ (_15550_, _15549_, _06717_);
  nand _48025_ (_15551_, _15550_, _15546_);
  nand _48026_ (_15552_, _15551_, _06751_);
  nand _48027_ (_15553_, _15552_, _15541_);
  nand _48028_ (_15554_, _15553_, _06760_);
  nand _48029_ (_15555_, _15554_, _15531_);
  nand _48030_ (_15556_, _15555_, _06780_);
  nand _48031_ (_15557_, _15556_, _15508_);
  nand _48032_ (_15558_, _15557_, _06734_);
  nand _48033_ (_15559_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand _48034_ (_15560_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand _48035_ (_15561_, _15560_, _15559_);
  nand _48036_ (_15562_, _15561_, _06717_);
  nand _48037_ (_15563_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nand _48038_ (_15564_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nand _48039_ (_15565_, _15564_, _15563_);
  nand _48040_ (_15567_, _15565_, _06716_);
  nand _48041_ (_15568_, _15567_, _15562_);
  nand _48042_ (_15569_, _15568_, _06748_);
  nand _48043_ (_15570_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand _48044_ (_15571_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand _48045_ (_15572_, _15571_, _15570_);
  nand _48046_ (_15573_, _15572_, _06717_);
  nand _48047_ (_15574_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nand _48048_ (_15575_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nand _48049_ (_15576_, _15575_, _15574_);
  nand _48050_ (_15577_, _15576_, _06716_);
  nand _48051_ (_15578_, _15577_, _15573_);
  nand _48052_ (_15579_, _15578_, _06751_);
  nand _48053_ (_15580_, _15579_, _15569_);
  nand _48054_ (_15581_, _15580_, _06761_);
  nor _48055_ (_15582_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor _48056_ (_15583_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _48057_ (_15584_, _15583_, _15582_);
  nand _48058_ (_15585_, _15584_, _06716_);
  nand _48059_ (_15586_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand _48060_ (_15587_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand _48061_ (_15588_, _15587_, _15586_);
  nand _48062_ (_15589_, _15588_, _06717_);
  nand _48063_ (_15590_, _15589_, _15585_);
  nand _48064_ (_15591_, _15590_, _06748_);
  nor _48065_ (_15592_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _48066_ (_15593_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor _48067_ (_15594_, _15593_, _15592_);
  nand _48068_ (_15595_, _15594_, _06716_);
  nand _48069_ (_15596_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand _48070_ (_15597_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand _48071_ (_15598_, _15597_, _15596_);
  nand _48072_ (_15599_, _15598_, _06717_);
  nand _48073_ (_15600_, _15599_, _15595_);
  nand _48074_ (_15601_, _15600_, _06751_);
  nand _48075_ (_15602_, _15601_, _15591_);
  nand _48076_ (_15603_, _15602_, _06760_);
  nand _48077_ (_15604_, _15603_, _15581_);
  nand _48078_ (_15605_, _15604_, _06780_);
  nand _48079_ (_15606_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nand _48080_ (_15607_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nand _48081_ (_15608_, _15607_, _15606_);
  nand _48082_ (_15609_, _15608_, _06717_);
  nand _48083_ (_15610_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nand _48084_ (_15611_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  nand _48085_ (_15612_, _15611_, _15610_);
  nand _48086_ (_15613_, _15612_, _06716_);
  nand _48087_ (_15614_, _15613_, _15609_);
  nand _48088_ (_15615_, _15614_, _06748_);
  nand _48089_ (_15616_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  nand _48090_ (_15617_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  nand _48091_ (_15618_, _15617_, _15616_);
  nand _48092_ (_15619_, _15618_, _06717_);
  nand _48093_ (_15620_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  nand _48094_ (_15621_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nand _48095_ (_15622_, _15621_, _15620_);
  nand _48096_ (_15623_, _15622_, _06716_);
  nand _48097_ (_15624_, _15623_, _15619_);
  nand _48098_ (_15625_, _15624_, _06751_);
  nand _48099_ (_15626_, _15625_, _15615_);
  nand _48100_ (_15627_, _15626_, _06761_);
  nor _48101_ (_15628_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nor _48102_ (_15629_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  nor _48103_ (_15630_, _15629_, _15628_);
  nand _48104_ (_15631_, _15630_, _06717_);
  nor _48105_ (_15632_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  nor _48106_ (_15633_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  nor _48107_ (_15634_, _15633_, _15632_);
  nand _48108_ (_15635_, _15634_, _06716_);
  nand _48109_ (_15636_, _15635_, _15631_);
  nand _48110_ (_15637_, _15636_, _06748_);
  nor _48111_ (_15638_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nor _48112_ (_15639_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  nor _48113_ (_15640_, _15639_, _15638_);
  nand _48114_ (_15641_, _15640_, _06717_);
  nor _48115_ (_15642_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nor _48116_ (_15643_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  nor _48117_ (_15644_, _15643_, _15642_);
  nand _48118_ (_15645_, _15644_, _06716_);
  nand _48119_ (_15646_, _15645_, _15641_);
  nand _48120_ (_15647_, _15646_, _06751_);
  nand _48121_ (_15648_, _15647_, _15637_);
  nand _48122_ (_15649_, _15648_, _06760_);
  nand _48123_ (_15650_, _15649_, _15627_);
  nand _48124_ (_15651_, _15650_, _06731_);
  nand _48125_ (_15652_, _15651_, _15605_);
  nand _48126_ (_15653_, _15652_, _06733_);
  nand _48127_ (_15654_, _15653_, _15558_);
  nor _48128_ (_15655_, _15654_, _06723_);
  nand _48129_ (_15656_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nand _48130_ (_15657_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nand _48131_ (_15658_, _15657_, _15656_);
  nand _48132_ (_15659_, _15658_, _06717_);
  nand _48133_ (_15660_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  nand _48134_ (_15661_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nand _48135_ (_15662_, _15661_, _15660_);
  nand _48136_ (_15663_, _15662_, _06716_);
  nand _48137_ (_15664_, _15663_, _15659_);
  nand _48138_ (_15665_, _15664_, _06748_);
  nand _48139_ (_15666_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nand _48140_ (_15667_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  nand _48141_ (_15668_, _15667_, _15666_);
  nand _48142_ (_15669_, _15668_, _06717_);
  nand _48143_ (_15670_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  nand _48144_ (_15671_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nand _48145_ (_15672_, _15671_, _15670_);
  nand _48146_ (_15673_, _15672_, _06716_);
  nand _48147_ (_15674_, _15673_, _15669_);
  nand _48148_ (_15675_, _15674_, _06751_);
  nand _48149_ (_15676_, _15675_, _15665_);
  nand _48150_ (_15677_, _15676_, _06761_);
  nor _48151_ (_15678_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  nor _48152_ (_15679_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  nor _48153_ (_15680_, _15679_, _15678_);
  nand _48154_ (_15681_, _15680_, _06716_);
  nand _48155_ (_15682_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  nand _48156_ (_15683_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nand _48157_ (_15684_, _15683_, _15682_);
  nand _48158_ (_15685_, _15684_, _06717_);
  nand _48159_ (_15686_, _15685_, _15681_);
  nand _48160_ (_15687_, _15686_, _06748_);
  nor _48161_ (_15688_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nor _48162_ (_15689_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  nor _48163_ (_15690_, _15689_, _15688_);
  nand _48164_ (_15691_, _15690_, _06716_);
  nand _48165_ (_15692_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nand _48166_ (_15693_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  nand _48167_ (_15694_, _15693_, _15692_);
  nand _48168_ (_15695_, _15694_, _06717_);
  nand _48169_ (_15696_, _15695_, _15691_);
  nand _48170_ (_15697_, _15696_, _06751_);
  nand _48171_ (_15698_, _15697_, _15687_);
  nand _48172_ (_15699_, _15698_, _06760_);
  nand _48173_ (_15700_, _15699_, _15677_);
  nand _48174_ (_15701_, _15700_, _06780_);
  nand _48175_ (_15702_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  nand _48176_ (_15703_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  nand _48177_ (_15704_, _15703_, _15702_);
  nand _48178_ (_15705_, _15704_, _06717_);
  nand _48179_ (_15706_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  nand _48180_ (_15707_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nand _48181_ (_15708_, _15707_, _15706_);
  nand _48182_ (_15709_, _15708_, _06716_);
  nand _48183_ (_15710_, _15709_, _15705_);
  nand _48184_ (_15711_, _15710_, _06748_);
  nand _48185_ (_15712_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nand _48186_ (_15713_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  nand _48187_ (_15714_, _15713_, _15712_);
  nand _48188_ (_15715_, _15714_, _06717_);
  nand _48189_ (_15716_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nand _48190_ (_15717_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nand _48191_ (_15718_, _15717_, _15716_);
  nand _48192_ (_15719_, _15718_, _06716_);
  nand _48193_ (_15720_, _15719_, _15715_);
  nand _48194_ (_15721_, _15720_, _06751_);
  nand _48195_ (_15722_, _15721_, _15711_);
  nand _48196_ (_15723_, _15722_, _06761_);
  nor _48197_ (_15724_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  nor _48198_ (_15725_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nor _48199_ (_15726_, _15725_, _15724_);
  nand _48200_ (_15727_, _15726_, _06717_);
  nor _48201_ (_15728_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nor _48202_ (_15729_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  nor _48203_ (_15730_, _15729_, _15728_);
  nand _48204_ (_15731_, _15730_, _06716_);
  nand _48205_ (_15732_, _15731_, _15727_);
  nand _48206_ (_15733_, _15732_, _06748_);
  nor _48207_ (_15734_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  nor _48208_ (_15735_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nor _48209_ (_15736_, _15735_, _15734_);
  nand _48210_ (_15737_, _15736_, _06717_);
  nor _48211_ (_15738_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  nor _48212_ (_15739_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  nor _48213_ (_15740_, _15739_, _15738_);
  nand _48214_ (_15741_, _15740_, _06716_);
  nand _48215_ (_15742_, _15741_, _15737_);
  nand _48216_ (_15743_, _15742_, _06751_);
  nand _48217_ (_15744_, _15743_, _15733_);
  nand _48218_ (_15745_, _15744_, _06760_);
  nand _48219_ (_15746_, _15745_, _15723_);
  nand _48220_ (_15747_, _15746_, _06731_);
  nand _48221_ (_15748_, _15747_, _15701_);
  nand _48222_ (_15749_, _15748_, _06734_);
  nor _48223_ (_15750_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nor _48224_ (_15751_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  nor _48225_ (_15752_, _15751_, _15750_);
  nand _48226_ (_15753_, _15752_, _06717_);
  nor _48227_ (_15754_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  nor _48228_ (_15755_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nor _48229_ (_15756_, _15755_, _15754_);
  nand _48230_ (_15757_, _15756_, _06716_);
  nand _48231_ (_15758_, _15757_, _15753_);
  nand _48232_ (_15759_, _15758_, _06751_);
  nor _48233_ (_15760_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nor _48234_ (_15761_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  nor _48235_ (_15762_, _15761_, _15760_);
  nand _48236_ (_15763_, _15762_, _06717_);
  nor _48237_ (_15764_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  nor _48238_ (_15765_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nor _48239_ (_15766_, _15765_, _15764_);
  nand _48240_ (_15767_, _15766_, _06716_);
  nand _48241_ (_15768_, _15767_, _15763_);
  nand _48242_ (_15769_, _15768_, _06748_);
  nand _48243_ (_15770_, _15769_, _15759_);
  nand _48244_ (_15771_, _15770_, _06760_);
  nand _48245_ (_15772_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  nand _48246_ (_15773_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nand _48247_ (_15774_, _15773_, _15772_);
  nand _48248_ (_15775_, _15774_, _06717_);
  nand _48249_ (_15776_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  nand _48250_ (_15777_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  nand _48251_ (_15778_, _15777_, _15776_);
  nand _48252_ (_15779_, _15778_, _06716_);
  nand _48253_ (_15780_, _15779_, _15775_);
  nand _48254_ (_15781_, _15780_, _06751_);
  nand _48255_ (_15782_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nand _48256_ (_15783_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nand _48257_ (_15784_, _15783_, _15782_);
  nand _48258_ (_15785_, _15784_, _06717_);
  nand _48259_ (_15786_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nand _48260_ (_15787_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  nand _48261_ (_15788_, _15787_, _15786_);
  nand _48262_ (_15789_, _15788_, _06716_);
  nand _48263_ (_15790_, _15789_, _15785_);
  nand _48264_ (_15791_, _15790_, _06748_);
  nand _48265_ (_15792_, _15791_, _15781_);
  nand _48266_ (_15793_, _15792_, _06761_);
  nand _48267_ (_15794_, _15793_, _15771_);
  nand _48268_ (_15795_, _15794_, _06731_);
  nor _48269_ (_15796_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  nor _48270_ (_15797_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  nor _48271_ (_15798_, _15797_, _15796_);
  nand _48272_ (_15799_, _15798_, _06716_);
  nand _48273_ (_15800_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  nand _48274_ (_15801_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  nand _48275_ (_15802_, _15801_, _15800_);
  nand _48276_ (_15803_, _15802_, _06717_);
  nand _48277_ (_15804_, _15803_, _15799_);
  nand _48278_ (_15805_, _15804_, _06751_);
  nor _48279_ (_15806_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nor _48280_ (_15807_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nor _48281_ (_15808_, _15807_, _15806_);
  nand _48282_ (_15809_, _15808_, _06716_);
  nand _48283_ (_15810_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  nand _48284_ (_15811_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  nand _48285_ (_15812_, _15811_, _15810_);
  nand _48286_ (_15813_, _15812_, _06717_);
  nand _48287_ (_15814_, _15813_, _15809_);
  nand _48288_ (_15815_, _15814_, _06748_);
  nand _48289_ (_15816_, _15815_, _15805_);
  nand _48290_ (_15817_, _15816_, _06760_);
  nand _48291_ (_15818_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  nand _48292_ (_15819_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  nand _48293_ (_15820_, _15819_, _15818_);
  nand _48294_ (_15821_, _15820_, _06717_);
  nand _48295_ (_15822_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nand _48296_ (_15823_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nand _48297_ (_15824_, _15823_, _15822_);
  nand _48298_ (_15825_, _15824_, _06716_);
  nand _48299_ (_15826_, _15825_, _15821_);
  nand _48300_ (_15827_, _15826_, _06751_);
  nand _48301_ (_15828_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nand _48302_ (_15829_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  nand _48303_ (_15830_, _15829_, _15828_);
  nand _48304_ (_15831_, _15830_, _06717_);
  nand _48305_ (_15832_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  nand _48306_ (_15833_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nand _48307_ (_15834_, _15833_, _15832_);
  nand _48308_ (_15835_, _15834_, _06716_);
  nand _48309_ (_15836_, _15835_, _15831_);
  nand _48310_ (_15837_, _15836_, _06748_);
  nand _48311_ (_15838_, _15837_, _15827_);
  nand _48312_ (_15839_, _15838_, _06761_);
  nand _48313_ (_15840_, _15839_, _15817_);
  nand _48314_ (_15841_, _15840_, _06780_);
  nand _48315_ (_15842_, _15841_, _15795_);
  nand _48316_ (_15843_, _15842_, _06733_);
  nand _48317_ (_15844_, _15843_, _15749_);
  nor _48318_ (_15845_, _15844_, _13106_);
  nor _48319_ (_15846_, _15845_, _15655_);
  nor _48320_ (_15847_, _15846_, _25929_);
  nand _48321_ (_15848_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  nand _48322_ (_15849_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nand _48323_ (_15850_, _15849_, _15848_);
  nand _48324_ (_15851_, _15850_, _06717_);
  nand _48325_ (_15852_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nand _48326_ (_15853_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  nand _48327_ (_15854_, _15853_, _15852_);
  nand _48328_ (_15855_, _15854_, _06716_);
  nand _48329_ (_15856_, _15855_, _15851_);
  nand _48330_ (_15858_, _15856_, _06748_);
  nand _48331_ (_15859_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nand _48332_ (_15860_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  nand _48333_ (_15861_, _15860_, _15859_);
  nand _48334_ (_15862_, _15861_, _06717_);
  nand _48335_ (_15863_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  nand _48336_ (_15864_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  nand _48337_ (_15865_, _15864_, _15863_);
  nand _48338_ (_15866_, _15865_, _06716_);
  nand _48339_ (_15867_, _15866_, _15862_);
  nand _48340_ (_15868_, _15867_, _06751_);
  nand _48341_ (_15869_, _15868_, _15858_);
  nand _48342_ (_15870_, _15869_, _06761_);
  nor _48343_ (_15871_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  nor _48344_ (_15872_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nor _48345_ (_15873_, _15872_, _15871_);
  nand _48346_ (_15874_, _15873_, _06716_);
  nand _48347_ (_15875_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  nand _48348_ (_15876_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nand _48349_ (_15877_, _15876_, _15875_);
  nand _48350_ (_15878_, _15877_, _06717_);
  nand _48351_ (_15879_, _15878_, _15874_);
  nand _48352_ (_15880_, _15879_, _06748_);
  nor _48353_ (_15881_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  nor _48354_ (_15882_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nor _48355_ (_15883_, _15882_, _15881_);
  nand _48356_ (_15884_, _15883_, _06716_);
  nand _48357_ (_15885_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  nand _48358_ (_15886_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nand _48359_ (_15887_, _15886_, _15885_);
  nand _48360_ (_15888_, _15887_, _06717_);
  nand _48361_ (_15889_, _15888_, _15884_);
  nand _48362_ (_15890_, _15889_, _06751_);
  nand _48363_ (_15891_, _15890_, _15880_);
  nand _48364_ (_15892_, _15891_, _06760_);
  nand _48365_ (_15893_, _15892_, _15870_);
  nand _48366_ (_15894_, _15893_, _06780_);
  nand _48367_ (_15895_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  nand _48368_ (_15896_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  nand _48369_ (_15897_, _15896_, _15895_);
  nand _48370_ (_15898_, _15897_, _06717_);
  nand _48371_ (_15899_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  nand _48372_ (_15900_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  nand _48373_ (_15901_, _15900_, _15899_);
  nand _48374_ (_15902_, _15901_, _06716_);
  nand _48375_ (_15903_, _15902_, _15898_);
  nand _48376_ (_15904_, _15903_, _06748_);
  nand _48377_ (_15905_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nand _48378_ (_15906_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nand _48379_ (_15907_, _15906_, _15905_);
  nand _48380_ (_15908_, _15907_, _06717_);
  nand _48381_ (_15909_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  nand _48382_ (_15910_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  nand _48383_ (_15911_, _15910_, _15909_);
  nand _48384_ (_15912_, _15911_, _06716_);
  nand _48385_ (_15913_, _15912_, _15908_);
  nand _48386_ (_15914_, _15913_, _06751_);
  nand _48387_ (_15915_, _15914_, _15904_);
  nand _48388_ (_15916_, _15915_, _06761_);
  nor _48389_ (_15917_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nor _48390_ (_15918_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nor _48391_ (_15919_, _15918_, _15917_);
  nand _48392_ (_15920_, _15919_, _06717_);
  nor _48393_ (_15921_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  nor _48394_ (_15922_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  nor _48395_ (_15923_, _15922_, _15921_);
  nand _48396_ (_15924_, _15923_, _06716_);
  nand _48397_ (_15925_, _15924_, _15920_);
  nand _48398_ (_15926_, _15925_, _06748_);
  nor _48399_ (_15927_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nor _48400_ (_15928_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nor _48401_ (_15929_, _15928_, _15927_);
  nand _48402_ (_15930_, _15929_, _06717_);
  nor _48403_ (_15931_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  nor _48404_ (_15932_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  nor _48405_ (_15933_, _15932_, _15931_);
  nand _48406_ (_15934_, _15933_, _06716_);
  nand _48407_ (_15935_, _15934_, _15930_);
  nand _48408_ (_15936_, _15935_, _06751_);
  nand _48409_ (_15937_, _15936_, _15926_);
  nand _48410_ (_15939_, _15937_, _06760_);
  nand _48411_ (_15940_, _15939_, _15916_);
  nand _48412_ (_15941_, _15940_, _06731_);
  nand _48413_ (_15942_, _15941_, _15894_);
  nand _48414_ (_15943_, _15942_, _06733_);
  nand _48415_ (_15944_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nand _48416_ (_15945_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  nand _48417_ (_15946_, _15945_, _15944_);
  nand _48418_ (_15947_, _15946_, _06717_);
  nand _48419_ (_15948_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  nand _48420_ (_15949_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nand _48421_ (_15950_, _15949_, _15948_);
  nand _48422_ (_15951_, _15950_, _06716_);
  nand _48423_ (_15952_, _15951_, _15947_);
  nand _48424_ (_15953_, _15952_, _06748_);
  nand _48425_ (_15954_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  nand _48426_ (_15955_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  nand _48427_ (_15956_, _15955_, _15954_);
  nand _48428_ (_15957_, _15956_, _06717_);
  nand _48429_ (_15958_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nand _48430_ (_15960_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  nand _48431_ (_15961_, _15960_, _15958_);
  nand _48432_ (_15962_, _15961_, _06716_);
  nand _48433_ (_15963_, _15962_, _15957_);
  nand _48434_ (_15964_, _15963_, _06751_);
  nand _48435_ (_15965_, _15964_, _15953_);
  nand _48436_ (_15966_, _15965_, _06761_);
  nor _48437_ (_15967_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  nor _48438_ (_15968_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  nor _48439_ (_15969_, _15968_, _15967_);
  nand _48440_ (_15970_, _15969_, _06717_);
  nor _48441_ (_15971_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  nor _48442_ (_15972_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nor _48443_ (_15973_, _15972_, _15971_);
  nand _48444_ (_15974_, _15973_, _06716_);
  nand _48445_ (_15975_, _15974_, _15970_);
  nand _48446_ (_15976_, _15975_, _06748_);
  nor _48447_ (_15977_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  nor _48448_ (_15978_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nor _48449_ (_15979_, _15978_, _15977_);
  nand _48450_ (_15980_, _15979_, _06717_);
  nor _48451_ (_15981_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  nor _48452_ (_15982_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  nor _48453_ (_15983_, _15982_, _15981_);
  nand _48454_ (_15984_, _15983_, _06716_);
  nand _48455_ (_15985_, _15984_, _15980_);
  nand _48456_ (_15986_, _15985_, _06751_);
  nand _48457_ (_15987_, _15986_, _15976_);
  nand _48458_ (_15988_, _15987_, _06760_);
  nand _48459_ (_15989_, _15988_, _15966_);
  nand _48460_ (_15991_, _15989_, _06731_);
  nand _48461_ (_15992_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nand _48462_ (_15993_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  nand _48463_ (_15994_, _15993_, _15992_);
  nand _48464_ (_15995_, _15994_, _06717_);
  nand _48465_ (_15996_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  nand _48466_ (_15997_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nand _48467_ (_15998_, _15997_, _15996_);
  nand _48468_ (_15999_, _15998_, _06716_);
  nand _48469_ (_16000_, _15999_, _15995_);
  nand _48470_ (_16001_, _16000_, _06748_);
  nand _48471_ (_16002_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nand _48472_ (_16003_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  nand _48473_ (_16004_, _16003_, _16002_);
  nand _48474_ (_16005_, _16004_, _06717_);
  nand _48475_ (_16006_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  nand _48476_ (_16007_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  nand _48477_ (_16008_, _16007_, _16006_);
  nand _48478_ (_16009_, _16008_, _06716_);
  nand _48479_ (_16010_, _16009_, _16005_);
  nand _48480_ (_16011_, _16010_, _06751_);
  nand _48481_ (_16012_, _16011_, _16001_);
  nand _48482_ (_16013_, _16012_, _06761_);
  nor _48483_ (_16014_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  nor _48484_ (_16015_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  nor _48485_ (_16016_, _16015_, _16014_);
  nand _48486_ (_16017_, _16016_, _06716_);
  nand _48487_ (_16018_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nand _48488_ (_16019_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nand _48489_ (_16020_, _16019_, _16018_);
  nand _48490_ (_16021_, _16020_, _06717_);
  nand _48491_ (_16022_, _16021_, _16017_);
  nand _48492_ (_16023_, _16022_, _06748_);
  nor _48493_ (_16024_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  nor _48494_ (_16025_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  nor _48495_ (_16026_, _16025_, _16024_);
  nand _48496_ (_16027_, _16026_, _06716_);
  nand _48497_ (_16028_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nand _48498_ (_16029_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nand _48499_ (_16030_, _16029_, _16028_);
  nand _48500_ (_16031_, _16030_, _06717_);
  nand _48501_ (_16032_, _16031_, _16027_);
  nand _48502_ (_16033_, _16032_, _06751_);
  nand _48503_ (_16034_, _16033_, _16023_);
  nand _48504_ (_16035_, _16034_, _06760_);
  nand _48505_ (_16036_, _16035_, _16013_);
  nand _48506_ (_16037_, _16036_, _06780_);
  nand _48507_ (_16038_, _16037_, _15991_);
  nand _48508_ (_16039_, _16038_, _06734_);
  nand _48509_ (_16040_, _16039_, _15943_);
  nor _48510_ (_16041_, _16040_, _06723_);
  nand _48511_ (_16042_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nand _48512_ (_16043_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  nand _48513_ (_16044_, _16043_, _16042_);
  nand _48514_ (_16045_, _16044_, _06716_);
  nand _48515_ (_16046_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  nand _48516_ (_16047_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  nand _48517_ (_16048_, _16047_, _16046_);
  nand _48518_ (_16049_, _16048_, _06717_);
  nand _48519_ (_16050_, _16049_, _16045_);
  nand _48520_ (_16051_, _16050_, _06748_);
  nand _48521_ (_16052_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  nand _48522_ (_16053_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  nand _48523_ (_16054_, _16053_, _16052_);
  nand _48524_ (_16055_, _16054_, _06716_);
  nand _48525_ (_16056_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nand _48526_ (_16057_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  nand _48527_ (_16058_, _16057_, _16056_);
  nand _48528_ (_16059_, _16058_, _06717_);
  nand _48529_ (_16060_, _16059_, _16055_);
  nand _48530_ (_16062_, _16060_, _06751_);
  nand _48531_ (_16063_, _16062_, _16051_);
  nand _48532_ (_16064_, _16063_, _06761_);
  nand _48533_ (_16065_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  nand _48534_ (_16066_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nand _48535_ (_16067_, _16066_, _16065_);
  nand _48536_ (_16068_, _16067_, _06717_);
  nor _48537_ (_16069_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  nor _48538_ (_16070_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nor _48539_ (_16071_, _16070_, _16069_);
  nand _48540_ (_16072_, _16071_, _06716_);
  nand _48541_ (_16073_, _16072_, _16068_);
  nand _48542_ (_16074_, _16073_, _06748_);
  nand _48543_ (_16075_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  nand _48544_ (_16076_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nand _48545_ (_16077_, _16076_, _16075_);
  nand _48546_ (_16078_, _16077_, _06717_);
  nor _48547_ (_16079_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  nor _48548_ (_16080_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nor _48549_ (_16081_, _16080_, _16079_);
  nand _48550_ (_16082_, _16081_, _06716_);
  nand _48551_ (_16083_, _16082_, _16078_);
  nand _48552_ (_16084_, _16083_, _06751_);
  nand _48553_ (_16085_, _16084_, _16074_);
  nand _48554_ (_16086_, _16085_, _06760_);
  nand _48555_ (_16087_, _16086_, _16064_);
  nand _48556_ (_16088_, _16087_, _06780_);
  nand _48557_ (_16089_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  nand _48558_ (_16090_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  nand _48559_ (_16091_, _16090_, _16089_);
  nand _48560_ (_16093_, _16091_, _06717_);
  nand _48561_ (_16094_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  nand _48562_ (_16095_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nand _48563_ (_16096_, _16095_, _16094_);
  nand _48564_ (_16097_, _16096_, _06716_);
  nand _48565_ (_16098_, _16097_, _16093_);
  nand _48566_ (_16099_, _16098_, _06748_);
  nand _48567_ (_16100_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  nand _48568_ (_16101_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nand _48569_ (_16102_, _16101_, _16100_);
  nand _48570_ (_16103_, _16102_, _06717_);
  nand _48571_ (_16104_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nand _48572_ (_16105_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  nand _48573_ (_16106_, _16105_, _16104_);
  nand _48574_ (_16107_, _16106_, _06716_);
  nand _48575_ (_16108_, _16107_, _16103_);
  nand _48576_ (_16109_, _16108_, _06751_);
  nand _48577_ (_16110_, _16109_, _16099_);
  nand _48578_ (_16111_, _16110_, _06761_);
  nor _48579_ (_16112_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  nor _48580_ (_16113_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  nor _48581_ (_16114_, _16113_, _16112_);
  nand _48582_ (_16115_, _16114_, _06717_);
  nor _48583_ (_16116_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  nor _48584_ (_16117_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nor _48585_ (_16118_, _16117_, _16116_);
  nand _48586_ (_16119_, _16118_, _06716_);
  nand _48587_ (_16120_, _16119_, _16115_);
  nand _48588_ (_16121_, _16120_, _06748_);
  nor _48589_ (_16122_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nor _48590_ (_16123_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  nor _48591_ (_16124_, _16123_, _16122_);
  nor _48592_ (_16125_, _16124_, _06716_);
  nor _48593_ (_16126_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  nor _48594_ (_16127_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nor _48595_ (_16128_, _16127_, _16126_);
  nor _48596_ (_16129_, _16128_, _06717_);
  nor _48597_ (_16130_, _16129_, _16125_);
  nand _48598_ (_16131_, _16130_, _06751_);
  nand _48599_ (_16132_, _16131_, _16121_);
  nand _48600_ (_16133_, _16132_, _06760_);
  nand _48601_ (_16134_, _16133_, _16111_);
  nand _48602_ (_16135_, _16134_, _06731_);
  nand _48603_ (_16136_, _16135_, _16088_);
  nand _48604_ (_16137_, _16136_, _06734_);
  nand _48605_ (_16138_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  nand _48606_ (_16139_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nand _48607_ (_16140_, _16139_, _16138_);
  nand _48608_ (_16141_, _16140_, _06717_);
  nand _48609_ (_16142_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  nand _48610_ (_16143_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  nand _48611_ (_16144_, _16143_, _16142_);
  nand _48612_ (_16145_, _16144_, _06716_);
  nand _48613_ (_16146_, _16145_, _16141_);
  nand _48614_ (_16147_, _16146_, _06748_);
  nand _48615_ (_16148_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  nand _48616_ (_16149_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nand _48617_ (_16150_, _16149_, _16148_);
  nand _48618_ (_16151_, _16150_, _06717_);
  nand _48619_ (_16152_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nand _48620_ (_16153_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  nand _48621_ (_16154_, _16153_, _16152_);
  nand _48622_ (_16155_, _16154_, _06716_);
  nand _48623_ (_16156_, _16155_, _16151_);
  nand _48624_ (_16157_, _16156_, _06751_);
  nand _48625_ (_16158_, _16157_, _16147_);
  nand _48626_ (_16159_, _16158_, _06761_);
  nor _48627_ (_16160_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  nor _48628_ (_16161_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  nor _48629_ (_16162_, _16161_, _16160_);
  nand _48630_ (_16164_, _16162_, _06717_);
  nor _48631_ (_16165_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  nor _48632_ (_16166_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nor _48633_ (_16167_, _16166_, _16165_);
  nand _48634_ (_16168_, _16167_, _06716_);
  nand _48635_ (_16169_, _16168_, _16164_);
  nand _48636_ (_16170_, _16169_, _06748_);
  nor _48637_ (_16171_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nor _48638_ (_16172_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  nor _48639_ (_16173_, _16172_, _16171_);
  nand _48640_ (_16174_, _16173_, _06717_);
  nor _48641_ (_16175_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nor _48642_ (_16176_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  nor _48643_ (_16177_, _16176_, _16175_);
  nand _48644_ (_16178_, _16177_, _06716_);
  nand _48645_ (_16179_, _16178_, _16174_);
  nand _48646_ (_16180_, _16179_, _06751_);
  nand _48647_ (_16181_, _16180_, _16170_);
  nand _48648_ (_16182_, _16181_, _06760_);
  nand _48649_ (_16183_, _16182_, _16159_);
  nand _48650_ (_16184_, _16183_, _06731_);
  nand _48651_ (_16185_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nand _48652_ (_16186_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  nand _48653_ (_16187_, _16186_, _16185_);
  nand _48654_ (_16188_, _16187_, _06717_);
  nand _48655_ (_16189_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  nand _48656_ (_16190_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  nand _48657_ (_16191_, _16190_, _16189_);
  nand _48658_ (_16192_, _16191_, _06716_);
  nand _48659_ (_16193_, _16192_, _16188_);
  nand _48660_ (_16194_, _16193_, _06748_);
  nand _48661_ (_16195_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nand _48662_ (_16196_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nand _48663_ (_16197_, _16196_, _16195_);
  nand _48664_ (_16198_, _16197_, _06717_);
  nand _48665_ (_16199_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  nand _48666_ (_16200_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  nand _48667_ (_16201_, _16200_, _16199_);
  nand _48668_ (_16202_, _16201_, _06716_);
  nand _48669_ (_16203_, _16202_, _16198_);
  nand _48670_ (_16204_, _16203_, _06751_);
  nand _48671_ (_16205_, _16204_, _16194_);
  nand _48672_ (_16206_, _16205_, _06761_);
  nor _48673_ (_16207_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nor _48674_ (_16208_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nor _48675_ (_16209_, _16208_, _16207_);
  nand _48676_ (_16210_, _16209_, _06717_);
  nor _48677_ (_16211_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  nor _48678_ (_16212_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  nor _48679_ (_16213_, _16212_, _16211_);
  nand _48680_ (_16214_, _16213_, _06716_);
  nand _48681_ (_16215_, _16214_, _16210_);
  nand _48682_ (_16216_, _16215_, _06748_);
  nor _48683_ (_16217_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  nor _48684_ (_16218_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  nor _48685_ (_16219_, _16218_, _16217_);
  nand _48686_ (_16220_, _16219_, _06717_);
  nor _48687_ (_16221_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nor _48688_ (_16222_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nor _48689_ (_16223_, _16222_, _16221_);
  nand _48690_ (_16224_, _16223_, _06716_);
  nand _48691_ (_16225_, _16224_, _16220_);
  nand _48692_ (_16226_, _16225_, _06751_);
  nand _48693_ (_16227_, _16226_, _16216_);
  nand _48694_ (_16228_, _16227_, _06760_);
  nand _48695_ (_16229_, _16228_, _16206_);
  nand _48696_ (_16230_, _16229_, _06780_);
  nand _48697_ (_16231_, _16230_, _16184_);
  nand _48698_ (_16232_, _16231_, _06733_);
  nand _48699_ (_16233_, _16232_, _16137_);
  nor _48700_ (_16234_, _16233_, _13106_);
  nor _48701_ (_16235_, _16234_, _16041_);
  nor _48702_ (_16236_, _16235_, _25843_);
  nor _48703_ (_16237_, _16236_, _15847_);
  nor _48704_ (_16238_, _16237_, _13105_);
  nand _48705_ (_16239_, _13105_, _24324_);
  nand _48706_ (_16240_, _16239_, _26487_);
  nor _48707_ (_06696_, _16240_, _16238_);
  nand _48708_ (_16241_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nand _48709_ (_16242_, _03867_, _24927_);
  nand _48710_ (_06699_, _16242_, _16241_);
  nand _48711_ (_16243_, _11827_, _24789_);
  nand _48712_ (_16244_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  nand _48713_ (_06702_, _16244_, _16243_);
  nand _48714_ (_16245_, _11827_, _25150_);
  nand _48715_ (_16246_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  nand _48716_ (_06707_, _16246_, _16245_);
  nand _48717_ (_16247_, _11931_, _25099_);
  nand _48718_ (_16248_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  nand _48719_ (_06710_, _16248_, _16247_);
  nand _48720_ (_16249_, _04308_, _28096_);
  nand _48721_ (_16250_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nand _48722_ (_06722_, _16250_, _16249_);
  nand _48723_ (_16251_, _11931_, _25203_);
  nand _48724_ (_16252_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  nand _48725_ (_06725_, _16252_, _16251_);
  nand _48726_ (_16253_, _13080_, _28096_);
  nand _48727_ (_16254_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  nand _48728_ (_06727_, _16254_, _16253_);
  nand _48729_ (_16255_, _03858_, _25203_);
  nand _48730_ (_16256_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  nand _48731_ (_06729_, _16256_, _16255_);
  nand _48732_ (_16257_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nand _48733_ (_16258_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nand _48734_ (_16259_, _16258_, _16257_);
  nand _48735_ (_16260_, _16259_, _06717_);
  nand _48736_ (_16261_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  nand _48737_ (_16262_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  nand _48738_ (_16263_, _16262_, _16261_);
  nand _48739_ (_16264_, _16263_, _06716_);
  nand _48740_ (_16266_, _16264_, _16260_);
  nand _48741_ (_16267_, _16266_, _06748_);
  nand _48742_ (_16268_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nand _48743_ (_16269_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nand _48744_ (_16270_, _16269_, _16268_);
  nand _48745_ (_16271_, _16270_, _06717_);
  nand _48746_ (_16272_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nand _48747_ (_16273_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  nand _48748_ (_16274_, _16273_, _16272_);
  nand _48749_ (_16275_, _16274_, _06716_);
  nand _48750_ (_16276_, _16275_, _16271_);
  nand _48751_ (_16277_, _16276_, _06751_);
  nand _48752_ (_16278_, _16277_, _16267_);
  nand _48753_ (_16279_, _16278_, _06761_);
  nor _48754_ (_16280_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  nor _48755_ (_16281_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nor _48756_ (_16282_, _16281_, _16280_);
  nand _48757_ (_16283_, _16282_, _06717_);
  nor _48758_ (_16284_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  nor _48759_ (_16285_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  nor _48760_ (_16286_, _16285_, _16284_);
  nand _48761_ (_16287_, _16286_, _06716_);
  nand _48762_ (_16288_, _16287_, _16283_);
  nand _48763_ (_16289_, _16288_, _06748_);
  nor _48764_ (_16290_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nor _48765_ (_16291_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nor _48766_ (_16292_, _16291_, _16290_);
  nand _48767_ (_16293_, _16292_, _06717_);
  nor _48768_ (_16294_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nor _48769_ (_16295_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  nor _48770_ (_16296_, _16295_, _16294_);
  nand _48771_ (_16297_, _16296_, _06716_);
  nand _48772_ (_16298_, _16297_, _16293_);
  nand _48773_ (_16299_, _16298_, _06751_);
  nand _48774_ (_16300_, _16299_, _16289_);
  nand _48775_ (_16301_, _16300_, _06760_);
  nand _48776_ (_16302_, _16301_, _16279_);
  nand _48777_ (_16303_, _16302_, _06731_);
  nand _48778_ (_16304_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  nand _48779_ (_16305_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  nand _48780_ (_16307_, _16305_, _16304_);
  nand _48781_ (_16308_, _16307_, _06717_);
  nand _48782_ (_16309_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nand _48783_ (_16310_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nand _48784_ (_16311_, _16310_, _16309_);
  nand _48785_ (_16312_, _16311_, _06716_);
  nand _48786_ (_16313_, _16312_, _16308_);
  nand _48787_ (_16314_, _16313_, _06748_);
  nand _48788_ (_16315_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  nand _48789_ (_16316_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  nand _48790_ (_16317_, _16316_, _16315_);
  nand _48791_ (_16318_, _16317_, _06717_);
  nand _48792_ (_16319_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nand _48793_ (_16320_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nand _48794_ (_16321_, _16320_, _16319_);
  nand _48795_ (_16322_, _16321_, _06716_);
  nand _48796_ (_16323_, _16322_, _16318_);
  nand _48797_ (_16324_, _16323_, _06751_);
  nand _48798_ (_16325_, _16324_, _16314_);
  nand _48799_ (_16326_, _16325_, _06761_);
  nor _48800_ (_16328_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  nor _48801_ (_16329_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  nor _48802_ (_16330_, _16329_, _16328_);
  nand _48803_ (_16331_, _16330_, _06716_);
  nand _48804_ (_16332_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  nand _48805_ (_16333_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nand _48806_ (_16334_, _16333_, _16332_);
  nand _48807_ (_16335_, _16334_, _06717_);
  nand _48808_ (_16336_, _16335_, _16331_);
  nand _48809_ (_16337_, _16336_, _06748_);
  nor _48810_ (_16338_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  nor _48811_ (_16339_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  nor _48812_ (_16340_, _16339_, _16338_);
  nand _48813_ (_16341_, _16340_, _06716_);
  nand _48814_ (_16342_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  nand _48815_ (_16343_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nand _48816_ (_16344_, _16343_, _16342_);
  nand _48817_ (_16345_, _16344_, _06717_);
  nand _48818_ (_16346_, _16345_, _16341_);
  nand _48819_ (_16347_, _16346_, _06751_);
  nand _48820_ (_16348_, _16347_, _16337_);
  nand _48821_ (_16349_, _16348_, _06760_);
  nand _48822_ (_16350_, _16349_, _16326_);
  nand _48823_ (_16351_, _16350_, _06780_);
  nand _48824_ (_16352_, _16351_, _16303_);
  nand _48825_ (_16353_, _16352_, _06734_);
  nand _48826_ (_16354_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nand _48827_ (_16355_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand _48828_ (_16356_, _16355_, _16354_);
  nand _48829_ (_16357_, _16356_, _06717_);
  nand _48830_ (_16358_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nand _48831_ (_16359_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand _48832_ (_16360_, _16359_, _16358_);
  nand _48833_ (_16361_, _16360_, _06716_);
  nand _48834_ (_16362_, _16361_, _16357_);
  nand _48835_ (_16363_, _16362_, _06748_);
  nand _48836_ (_16364_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nand _48837_ (_16365_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nand _48838_ (_16366_, _16365_, _16364_);
  nand _48839_ (_16367_, _16366_, _06717_);
  nand _48840_ (_16368_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nand _48841_ (_16369_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nand _48842_ (_16370_, _16369_, _16368_);
  nand _48843_ (_16371_, _16370_, _06716_);
  nand _48844_ (_16372_, _16371_, _16367_);
  nand _48845_ (_16373_, _16372_, _06751_);
  nand _48846_ (_16374_, _16373_, _16363_);
  nand _48847_ (_16375_, _16374_, _06761_);
  nor _48848_ (_16376_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _48849_ (_16377_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _48850_ (_16378_, _16377_, _16376_);
  nand _48851_ (_16379_, _16378_, _06716_);
  nand _48852_ (_16380_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nand _48853_ (_16381_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nand _48854_ (_16382_, _16381_, _16380_);
  nand _48855_ (_16383_, _16382_, _06717_);
  nand _48856_ (_16384_, _16383_, _16379_);
  nand _48857_ (_16385_, _16384_, _06748_);
  nor _48858_ (_16386_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _48859_ (_16387_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor _48860_ (_16388_, _16387_, _16386_);
  nand _48861_ (_16389_, _16388_, _06716_);
  nand _48862_ (_16390_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nand _48863_ (_16391_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nand _48864_ (_16392_, _16391_, _16390_);
  nand _48865_ (_16393_, _16392_, _06717_);
  nand _48866_ (_16394_, _16393_, _16389_);
  nand _48867_ (_16395_, _16394_, _06751_);
  nand _48868_ (_16396_, _16395_, _16385_);
  nand _48869_ (_16397_, _16396_, _06760_);
  nand _48870_ (_16398_, _16397_, _16375_);
  nand _48871_ (_16399_, _16398_, _06780_);
  nand _48872_ (_16400_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nand _48873_ (_16401_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  nand _48874_ (_16402_, _16401_, _16400_);
  nand _48875_ (_16403_, _16402_, _06717_);
  nand _48876_ (_16404_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  nand _48877_ (_16405_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nand _48878_ (_16406_, _16405_, _16404_);
  nand _48879_ (_16407_, _16406_, _06716_);
  nand _48880_ (_16408_, _16407_, _16403_);
  nand _48881_ (_16409_, _16408_, _06748_);
  nand _48882_ (_16410_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nand _48883_ (_16411_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nand _48884_ (_16412_, _16411_, _16410_);
  nand _48885_ (_16413_, _16412_, _06717_);
  nand _48886_ (_16414_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nand _48887_ (_16415_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  nand _48888_ (_16416_, _16415_, _16414_);
  nand _48889_ (_16417_, _16416_, _06716_);
  nand _48890_ (_16418_, _16417_, _16413_);
  nand _48891_ (_16419_, _16418_, _06751_);
  nand _48892_ (_16420_, _16419_, _16409_);
  nand _48893_ (_16421_, _16420_, _06761_);
  nor _48894_ (_16422_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  nor _48895_ (_16423_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nor _48896_ (_16424_, _16423_, _16422_);
  nand _48897_ (_16425_, _16424_, _06717_);
  nor _48898_ (_16426_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  nor _48899_ (_16427_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  nor _48900_ (_16428_, _16427_, _16426_);
  nand _48901_ (_16429_, _16428_, _06716_);
  nand _48902_ (_16430_, _16429_, _16425_);
  nand _48903_ (_16431_, _16430_, _06748_);
  nor _48904_ (_16432_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nor _48905_ (_16433_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  nor _48906_ (_16434_, _16433_, _16432_);
  nand _48907_ (_16435_, _16434_, _06717_);
  nor _48908_ (_16436_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  nor _48909_ (_16437_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  nor _48910_ (_16438_, _16437_, _16436_);
  nand _48911_ (_16439_, _16438_, _06716_);
  nand _48912_ (_16440_, _16439_, _16435_);
  nand _48913_ (_16441_, _16440_, _06751_);
  nand _48914_ (_16442_, _16441_, _16431_);
  nand _48915_ (_16443_, _16442_, _06760_);
  nand _48916_ (_16444_, _16443_, _16421_);
  nand _48917_ (_16445_, _16444_, _06731_);
  nand _48918_ (_16446_, _16445_, _16399_);
  nand _48919_ (_16447_, _16446_, _06733_);
  nand _48920_ (_16448_, _16447_, _16353_);
  nor _48921_ (_16449_, _16448_, _06723_);
  nand _48922_ (_16450_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nand _48923_ (_16451_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nand _48924_ (_16452_, _16451_, _16450_);
  nand _48925_ (_16453_, _16452_, _06717_);
  nand _48926_ (_16454_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  nand _48927_ (_16455_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  nand _48928_ (_16456_, _16455_, _16454_);
  nand _48929_ (_16457_, _16456_, _06716_);
  nand _48930_ (_16458_, _16457_, _16453_);
  nand _48931_ (_16459_, _16458_, _06748_);
  nand _48932_ (_16460_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  nand _48933_ (_16461_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nand _48934_ (_16462_, _16461_, _16460_);
  nand _48935_ (_16463_, _16462_, _06717_);
  nand _48936_ (_16464_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nand _48937_ (_16465_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  nand _48938_ (_16466_, _16465_, _16464_);
  nand _48939_ (_16467_, _16466_, _06716_);
  nand _48940_ (_16468_, _16467_, _16463_);
  nand _48941_ (_16469_, _16468_, _06751_);
  nand _48942_ (_16470_, _16469_, _16459_);
  nand _48943_ (_16471_, _16470_, _06761_);
  nor _48944_ (_16472_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nor _48945_ (_16473_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  nor _48946_ (_16474_, _16473_, _16472_);
  nand _48947_ (_16475_, _16474_, _06716_);
  nand _48948_ (_16476_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nand _48949_ (_16477_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  nand _48950_ (_16478_, _16477_, _16476_);
  nand _48951_ (_16479_, _16478_, _06717_);
  nand _48952_ (_16480_, _16479_, _16475_);
  nand _48953_ (_16481_, _16480_, _06748_);
  nor _48954_ (_16482_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  nor _48955_ (_16483_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nor _48956_ (_16484_, _16483_, _16482_);
  nand _48957_ (_16485_, _16484_, _06716_);
  nand _48958_ (_16486_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nand _48959_ (_16487_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nand _48960_ (_16488_, _16487_, _16486_);
  nand _48961_ (_16489_, _16488_, _06717_);
  nand _48962_ (_16490_, _16489_, _16485_);
  nand _48963_ (_16491_, _16490_, _06751_);
  nand _48964_ (_16492_, _16491_, _16481_);
  nand _48965_ (_16493_, _16492_, _06760_);
  nand _48966_ (_16494_, _16493_, _16471_);
  nand _48967_ (_16495_, _16494_, _06780_);
  nand _48968_ (_16496_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  nand _48969_ (_16497_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nand _48970_ (_16498_, _16497_, _16496_);
  nand _48971_ (_16499_, _16498_, _06717_);
  nand _48972_ (_16500_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  nand _48973_ (_16501_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  nand _48974_ (_16502_, _16501_, _16500_);
  nand _48975_ (_16503_, _16502_, _06716_);
  nand _48976_ (_16504_, _16503_, _16499_);
  nand _48977_ (_16505_, _16504_, _06748_);
  nand _48978_ (_16506_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nand _48979_ (_16507_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nand _48980_ (_16508_, _16507_, _16506_);
  nand _48981_ (_16509_, _16508_, _06717_);
  nand _48982_ (_16510_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  nand _48983_ (_16511_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  nand _48984_ (_16512_, _16511_, _16510_);
  nand _48985_ (_16513_, _16512_, _06716_);
  nand _48986_ (_16514_, _16513_, _16509_);
  nand _48987_ (_16515_, _16514_, _06751_);
  nand _48988_ (_16516_, _16515_, _16505_);
  nand _48989_ (_16517_, _16516_, _06761_);
  nor _48990_ (_16518_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nor _48991_ (_16519_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  nor _48992_ (_16520_, _16519_, _16518_);
  nand _48993_ (_16521_, _16520_, _06717_);
  nor _48994_ (_16522_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nor _48995_ (_16523_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nor _48996_ (_16524_, _16523_, _16522_);
  nand _48997_ (_16525_, _16524_, _06716_);
  nand _48998_ (_16526_, _16525_, _16521_);
  nand _48999_ (_16527_, _16526_, _06748_);
  nor _49000_ (_16528_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  nor _49001_ (_16529_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nor _49002_ (_16530_, _16529_, _16528_);
  nand _49003_ (_16531_, _16530_, _06717_);
  nor _49004_ (_16532_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nor _49005_ (_16533_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  nor _49006_ (_16534_, _16533_, _16532_);
  nand _49007_ (_16535_, _16534_, _06716_);
  nand _49008_ (_16536_, _16535_, _16531_);
  nand _49009_ (_16537_, _16536_, _06751_);
  nand _49010_ (_16538_, _16537_, _16527_);
  nand _49011_ (_16539_, _16538_, _06760_);
  nand _49012_ (_16540_, _16539_, _16517_);
  nand _49013_ (_16541_, _16540_, _06731_);
  nand _49014_ (_16542_, _16541_, _16495_);
  nand _49015_ (_16543_, _16542_, _06734_);
  nor _49016_ (_16544_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nor _49017_ (_16545_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  nor _49018_ (_16546_, _16545_, _16544_);
  nand _49019_ (_16547_, _16546_, _06717_);
  nor _49020_ (_16548_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  nor _49021_ (_16549_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nor _49022_ (_16550_, _16549_, _16548_);
  nand _49023_ (_16551_, _16550_, _06716_);
  nand _49024_ (_16552_, _16551_, _16547_);
  nand _49025_ (_16553_, _16552_, _06751_);
  nor _49026_ (_16554_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  nor _49027_ (_16555_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  nor _49028_ (_16556_, _16555_, _16554_);
  nand _49029_ (_16557_, _16556_, _06717_);
  nor _49030_ (_16558_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  nor _49031_ (_16559_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nor _49032_ (_16560_, _16559_, _16558_);
  nand _49033_ (_16561_, _16560_, _06716_);
  nand _49034_ (_16562_, _16561_, _16557_);
  nand _49035_ (_16563_, _16562_, _06748_);
  nand _49036_ (_16564_, _16563_, _16553_);
  nand _49037_ (_16565_, _16564_, _06760_);
  nand _49038_ (_16566_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  nand _49039_ (_16567_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nand _49040_ (_16568_, _16567_, _16566_);
  nand _49041_ (_16569_, _16568_, _06717_);
  nand _49042_ (_16570_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nand _49043_ (_16571_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  nand _49044_ (_16572_, _16571_, _16570_);
  nand _49045_ (_16573_, _16572_, _06716_);
  nand _49046_ (_16574_, _16573_, _16569_);
  nand _49047_ (_16575_, _16574_, _06751_);
  nand _49048_ (_16576_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  nand _49049_ (_16577_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  nand _49050_ (_16579_, _16577_, _16576_);
  nand _49051_ (_16580_, _16579_, _06717_);
  nand _49052_ (_16581_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nand _49053_ (_16582_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nand _49054_ (_16583_, _16582_, _16581_);
  nand _49055_ (_16584_, _16583_, _06716_);
  nand _49056_ (_16585_, _16584_, _16580_);
  nand _49057_ (_16586_, _16585_, _06748_);
  nand _49058_ (_16587_, _16586_, _16575_);
  nand _49059_ (_16588_, _16587_, _06761_);
  nand _49060_ (_16589_, _16588_, _16565_);
  nand _49061_ (_16590_, _16589_, _06731_);
  nor _49062_ (_16591_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  nor _49063_ (_16592_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nor _49064_ (_16593_, _16592_, _16591_);
  nand _49065_ (_16594_, _16593_, _06716_);
  nand _49066_ (_16595_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  nand _49067_ (_16596_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nand _49068_ (_16597_, _16596_, _16595_);
  nand _49069_ (_16598_, _16597_, _06717_);
  nand _49070_ (_16599_, _16598_, _16594_);
  nand _49071_ (_16600_, _16599_, _06751_);
  nor _49072_ (_16601_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nor _49073_ (_16602_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nor _49074_ (_16603_, _16602_, _16601_);
  nand _49075_ (_16604_, _16603_, _06716_);
  nand _49076_ (_16605_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nand _49077_ (_16606_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  nand _49078_ (_16607_, _16606_, _16605_);
  nand _49079_ (_16608_, _16607_, _06717_);
  nand _49080_ (_16609_, _16608_, _16604_);
  nand _49081_ (_16610_, _16609_, _06748_);
  nand _49082_ (_16611_, _16610_, _16600_);
  nand _49083_ (_16612_, _16611_, _06760_);
  nand _49084_ (_16613_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  nand _49085_ (_16614_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  nand _49086_ (_16615_, _16614_, _16613_);
  nand _49087_ (_16616_, _16615_, _06717_);
  nand _49088_ (_16617_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nand _49089_ (_16618_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  nand _49090_ (_16619_, _16618_, _16617_);
  nand _49091_ (_16620_, _16619_, _06716_);
  nand _49092_ (_16621_, _16620_, _16616_);
  nand _49093_ (_16622_, _16621_, _06751_);
  nand _49094_ (_16623_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  nand _49095_ (_16624_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  nand _49096_ (_16625_, _16624_, _16623_);
  nand _49097_ (_16626_, _16625_, _06717_);
  nand _49098_ (_16627_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  nand _49099_ (_16628_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nand _49100_ (_16629_, _16628_, _16627_);
  nand _49101_ (_16630_, _16629_, _06716_);
  nand _49102_ (_16631_, _16630_, _16626_);
  nand _49103_ (_16632_, _16631_, _06748_);
  nand _49104_ (_16633_, _16632_, _16622_);
  nand _49105_ (_16634_, _16633_, _06761_);
  nand _49106_ (_16635_, _16634_, _16612_);
  nand _49107_ (_16636_, _16635_, _06780_);
  nand _49108_ (_16637_, _16636_, _16590_);
  nand _49109_ (_16638_, _16637_, _06733_);
  nand _49110_ (_16639_, _16638_, _16543_);
  nor _49111_ (_16640_, _16639_, _13106_);
  nor _49112_ (_16641_, _16640_, _16449_);
  nor _49113_ (_16642_, _16641_, _25929_);
  nand _49114_ (_16643_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nand _49115_ (_16644_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  nand _49116_ (_16645_, _16644_, _16643_);
  nand _49117_ (_16646_, _16645_, _06717_);
  nand _49118_ (_16647_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  nand _49119_ (_16648_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  nand _49120_ (_16649_, _16648_, _16647_);
  nand _49121_ (_16650_, _16649_, _06716_);
  nand _49122_ (_16651_, _16650_, _16646_);
  nand _49123_ (_16652_, _16651_, _06748_);
  nand _49124_ (_16653_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  nand _49125_ (_16654_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nand _49126_ (_16655_, _16654_, _16653_);
  nand _49127_ (_16656_, _16655_, _06717_);
  nand _49128_ (_16657_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nand _49129_ (_16658_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  nand _49130_ (_16659_, _16658_, _16657_);
  nand _49131_ (_16660_, _16659_, _06716_);
  nand _49132_ (_16661_, _16660_, _16656_);
  nand _49133_ (_16662_, _16661_, _06751_);
  nand _49134_ (_16663_, _16662_, _16652_);
  nand _49135_ (_16664_, _16663_, _06761_);
  nor _49136_ (_16665_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  nor _49137_ (_16666_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  nor _49138_ (_16667_, _16666_, _16665_);
  nand _49139_ (_16668_, _16667_, _06716_);
  nand _49140_ (_16669_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nand _49141_ (_16670_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nand _49142_ (_16671_, _16670_, _16669_);
  nand _49143_ (_16672_, _16671_, _06717_);
  nand _49144_ (_16673_, _16672_, _16668_);
  nand _49145_ (_16674_, _16673_, _06748_);
  nor _49146_ (_16675_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  nor _49147_ (_16676_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor _49148_ (_16677_, _16676_, _16675_);
  nand _49149_ (_16678_, _16677_, _06716_);
  nand _49150_ (_16679_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nand _49151_ (_16680_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nand _49152_ (_16681_, _16680_, _16679_);
  nand _49153_ (_16682_, _16681_, _06717_);
  nand _49154_ (_16683_, _16682_, _16678_);
  nand _49155_ (_16684_, _16683_, _06751_);
  nand _49156_ (_16685_, _16684_, _16674_);
  nand _49157_ (_16686_, _16685_, _06760_);
  nand _49158_ (_16687_, _16686_, _16664_);
  nand _49159_ (_16688_, _16687_, _06780_);
  nand _49160_ (_16689_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  nand _49161_ (_16690_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  nand _49162_ (_16691_, _16690_, _16689_);
  nand _49163_ (_16692_, _16691_, _06717_);
  nand _49164_ (_16693_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nand _49165_ (_16694_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nand _49166_ (_16695_, _16694_, _16693_);
  nand _49167_ (_16696_, _16695_, _06716_);
  nand _49168_ (_16697_, _16696_, _16692_);
  nand _49169_ (_16698_, _16697_, _06748_);
  nand _49170_ (_16700_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  nand _49171_ (_16701_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  nand _49172_ (_16702_, _16701_, _16700_);
  nand _49173_ (_16703_, _16702_, _06717_);
  nand _49174_ (_16704_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nand _49175_ (_16705_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  nand _49176_ (_16706_, _16705_, _16704_);
  nand _49177_ (_16707_, _16706_, _06716_);
  nand _49178_ (_16708_, _16707_, _16703_);
  nand _49179_ (_16709_, _16708_, _06751_);
  nand _49180_ (_16710_, _16709_, _16698_);
  nand _49181_ (_16711_, _16710_, _06761_);
  nor _49182_ (_16712_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  nor _49183_ (_16713_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  nor _49184_ (_16714_, _16713_, _16712_);
  nand _49185_ (_16715_, _16714_, _06717_);
  nor _49186_ (_16716_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nor _49187_ (_16717_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  nor _49188_ (_16718_, _16717_, _16716_);
  nand _49189_ (_16719_, _16718_, _06716_);
  nand _49190_ (_16720_, _16719_, _16715_);
  nand _49191_ (_16721_, _16720_, _06748_);
  nor _49192_ (_16722_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  nor _49193_ (_16723_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nor _49194_ (_16724_, _16723_, _16722_);
  nand _49195_ (_16725_, _16724_, _06717_);
  nor _49196_ (_16726_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  nor _49197_ (_16727_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  nor _49198_ (_16728_, _16727_, _16726_);
  nand _49199_ (_16729_, _16728_, _06716_);
  nand _49200_ (_16730_, _16729_, _16725_);
  nand _49201_ (_16731_, _16730_, _06751_);
  nand _49202_ (_16732_, _16731_, _16721_);
  nand _49203_ (_16733_, _16732_, _06760_);
  nand _49204_ (_16734_, _16733_, _16711_);
  nand _49205_ (_16735_, _16734_, _06731_);
  nand _49206_ (_16736_, _16735_, _16688_);
  nand _49207_ (_16737_, _16736_, _06733_);
  nand _49208_ (_16738_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  nand _49209_ (_16739_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  nand _49210_ (_16740_, _16739_, _16738_);
  nand _49211_ (_16741_, _16740_, _06717_);
  nand _49212_ (_16742_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  nand _49213_ (_16743_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  nand _49214_ (_16744_, _16743_, _16742_);
  nand _49215_ (_16745_, _16744_, _06716_);
  nand _49216_ (_16746_, _16745_, _16741_);
  nand _49217_ (_16747_, _16746_, _06748_);
  nand _49218_ (_16748_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nand _49219_ (_16749_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nand _49220_ (_16750_, _16749_, _16748_);
  nand _49221_ (_16751_, _16750_, _06717_);
  nand _49222_ (_16752_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  nand _49223_ (_16753_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  nand _49224_ (_16754_, _16753_, _16752_);
  nand _49225_ (_16755_, _16754_, _06716_);
  nand _49226_ (_16756_, _16755_, _16751_);
  nand _49227_ (_16757_, _16756_, _06751_);
  nand _49228_ (_16758_, _16757_, _16747_);
  nand _49229_ (_16759_, _16758_, _06761_);
  nor _49230_ (_16760_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nor _49231_ (_16761_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  nor _49232_ (_16762_, _16761_, _16760_);
  nand _49233_ (_16763_, _16762_, _06717_);
  nor _49234_ (_16764_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nor _49235_ (_16765_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nor _49236_ (_16766_, _16765_, _16764_);
  nand _49237_ (_16767_, _16766_, _06716_);
  nand _49238_ (_16768_, _16767_, _16763_);
  nand _49239_ (_16769_, _16768_, _06748_);
  nor _49240_ (_16770_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  nor _49241_ (_16771_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  nor _49242_ (_16772_, _16771_, _16770_);
  nand _49243_ (_16773_, _16772_, _06717_);
  nor _49244_ (_16774_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  nor _49245_ (_16775_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nor _49246_ (_16776_, _16775_, _16774_);
  nand _49247_ (_16777_, _16776_, _06716_);
  nand _49248_ (_16778_, _16777_, _16773_);
  nand _49249_ (_16779_, _16778_, _06751_);
  nand _49250_ (_16781_, _16779_, _16769_);
  nand _49251_ (_16782_, _16781_, _06760_);
  nand _49252_ (_16783_, _16782_, _16759_);
  nand _49253_ (_16784_, _16783_, _06731_);
  nand _49254_ (_16785_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nand _49255_ (_16786_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  nand _49256_ (_16787_, _16786_, _16785_);
  nand _49257_ (_16788_, _16787_, _06717_);
  nand _49258_ (_16789_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  nand _49259_ (_16790_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nand _49260_ (_16791_, _16790_, _16789_);
  nand _49261_ (_16792_, _16791_, _06716_);
  nand _49262_ (_16793_, _16792_, _16788_);
  nand _49263_ (_16794_, _16793_, _06748_);
  nand _49264_ (_16795_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nand _49265_ (_16796_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  nand _49266_ (_16797_, _16796_, _16795_);
  nand _49267_ (_16798_, _16797_, _06717_);
  nand _49268_ (_16799_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  nand _49269_ (_16800_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  nand _49270_ (_16801_, _16800_, _16799_);
  nand _49271_ (_16802_, _16801_, _06716_);
  nand _49272_ (_16803_, _16802_, _16798_);
  nand _49273_ (_16804_, _16803_, _06751_);
  nand _49274_ (_16805_, _16804_, _16794_);
  nand _49275_ (_16806_, _16805_, _06761_);
  nor _49276_ (_16807_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  nor _49277_ (_16808_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  nor _49278_ (_16809_, _16808_, _16807_);
  nand _49279_ (_16810_, _16809_, _06716_);
  nand _49280_ (_16811_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nand _49281_ (_16812_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  nand _49282_ (_16813_, _16812_, _16811_);
  nand _49283_ (_16814_, _16813_, _06717_);
  nand _49284_ (_16815_, _16814_, _16810_);
  nand _49285_ (_16816_, _16815_, _06748_);
  nor _49286_ (_16817_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  nor _49287_ (_16818_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nor _49288_ (_16819_, _16818_, _16817_);
  nand _49289_ (_16820_, _16819_, _06716_);
  nand _49290_ (_16821_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nand _49291_ (_16822_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nand _49292_ (_16823_, _16822_, _16821_);
  nand _49293_ (_16824_, _16823_, _06717_);
  nand _49294_ (_16825_, _16824_, _16820_);
  nand _49295_ (_16826_, _16825_, _06751_);
  nand _49296_ (_16827_, _16826_, _16816_);
  nand _49297_ (_16828_, _16827_, _06760_);
  nand _49298_ (_16829_, _16828_, _16806_);
  nand _49299_ (_16830_, _16829_, _06780_);
  nand _49300_ (_16831_, _16830_, _16784_);
  nand _49301_ (_16832_, _16831_, _06734_);
  nand _49302_ (_16833_, _16832_, _16737_);
  nor _49303_ (_16834_, _16833_, _06723_);
  nand _49304_ (_16835_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nand _49305_ (_16836_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nand _49306_ (_16837_, _16836_, _16835_);
  nand _49307_ (_16838_, _16837_, _06716_);
  nand _49308_ (_16839_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  nand _49309_ (_16840_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nand _49310_ (_16842_, _16840_, _16839_);
  nand _49311_ (_16843_, _16842_, _06717_);
  nand _49312_ (_16844_, _16843_, _16838_);
  nand _49313_ (_16845_, _16844_, _06748_);
  nand _49314_ (_16846_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nand _49315_ (_16847_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  nand _49316_ (_16848_, _16847_, _16846_);
  nand _49317_ (_16849_, _16848_, _06716_);
  nand _49318_ (_16850_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  nand _49319_ (_16851_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  nand _49320_ (_16852_, _16851_, _16850_);
  nand _49321_ (_16853_, _16852_, _06717_);
  nand _49322_ (_16854_, _16853_, _16849_);
  nand _49323_ (_16855_, _16854_, _06751_);
  nand _49324_ (_16856_, _16855_, _16845_);
  nand _49325_ (_16857_, _16856_, _06761_);
  nand _49326_ (_16858_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nand _49327_ (_16859_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nand _49328_ (_16860_, _16859_, _16858_);
  nand _49329_ (_16861_, _16860_, _06717_);
  nor _49330_ (_16862_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  nor _49331_ (_16863_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nor _49332_ (_16864_, _16863_, _16862_);
  nand _49333_ (_16865_, _16864_, _06716_);
  nand _49334_ (_16866_, _16865_, _16861_);
  nand _49335_ (_16867_, _16866_, _06748_);
  nand _49336_ (_16868_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  nand _49337_ (_16869_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nand _49338_ (_16870_, _16869_, _16868_);
  nand _49339_ (_16871_, _16870_, _06717_);
  nor _49340_ (_16872_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  nor _49341_ (_16873_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  nor _49342_ (_16874_, _16873_, _16872_);
  nand _49343_ (_16875_, _16874_, _06716_);
  nand _49344_ (_16876_, _16875_, _16871_);
  nand _49345_ (_16877_, _16876_, _06751_);
  nand _49346_ (_16878_, _16877_, _16867_);
  nand _49347_ (_16879_, _16878_, _06760_);
  nand _49348_ (_16880_, _16879_, _16857_);
  nand _49349_ (_16881_, _16880_, _06780_);
  nand _49350_ (_16882_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nand _49351_ (_16883_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  nand _49352_ (_16884_, _16883_, _16882_);
  nand _49353_ (_16885_, _16884_, _06717_);
  nand _49354_ (_16886_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nand _49355_ (_16887_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  nand _49356_ (_16888_, _16887_, _16886_);
  nand _49357_ (_16889_, _16888_, _06716_);
  nand _49358_ (_16890_, _16889_, _16885_);
  nand _49359_ (_16891_, _16890_, _06748_);
  nand _49360_ (_16892_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  nand _49361_ (_16893_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  nand _49362_ (_16894_, _16893_, _16892_);
  nand _49363_ (_16895_, _16894_, _06717_);
  nand _49364_ (_16896_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  nand _49365_ (_16897_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nand _49366_ (_16898_, _16897_, _16896_);
  nand _49367_ (_16899_, _16898_, _06716_);
  nand _49368_ (_16900_, _16899_, _16895_);
  nand _49369_ (_16901_, _16900_, _06751_);
  nand _49370_ (_16903_, _16901_, _16891_);
  nand _49371_ (_16904_, _16903_, _06761_);
  nor _49372_ (_16905_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nor _49373_ (_16906_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  nor _49374_ (_16907_, _16906_, _16905_);
  nand _49375_ (_16908_, _16907_, _06717_);
  nor _49376_ (_16909_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nor _49377_ (_16910_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  nor _49378_ (_16911_, _16910_, _16909_);
  nand _49379_ (_16912_, _16911_, _06716_);
  nand _49380_ (_16913_, _16912_, _16908_);
  nand _49381_ (_16914_, _16913_, _06748_);
  nor _49382_ (_16915_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nor _49383_ (_16916_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  nor _49384_ (_16917_, _16916_, _16915_);
  nor _49385_ (_16918_, _16917_, _06716_);
  nor _49386_ (_16919_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  nor _49387_ (_16920_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nor _49388_ (_16921_, _16920_, _16919_);
  nor _49389_ (_16922_, _16921_, _06717_);
  nor _49390_ (_16924_, _16922_, _16918_);
  nand _49391_ (_16925_, _16924_, _06751_);
  nand _49392_ (_16926_, _16925_, _16914_);
  nand _49393_ (_16927_, _16926_, _06760_);
  nand _49394_ (_16928_, _16927_, _16904_);
  nand _49395_ (_16929_, _16928_, _06731_);
  nand _49396_ (_16930_, _16929_, _16881_);
  nand _49397_ (_16931_, _16930_, _06734_);
  nand _49398_ (_16932_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nand _49399_ (_16933_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  nand _49400_ (_16934_, _16933_, _16932_);
  nand _49401_ (_16935_, _16934_, _06717_);
  nand _49402_ (_16936_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  nand _49403_ (_16937_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nand _49404_ (_16938_, _16937_, _16936_);
  nand _49405_ (_16939_, _16938_, _06716_);
  nand _49406_ (_16940_, _16939_, _16935_);
  nand _49407_ (_16941_, _16940_, _06748_);
  nand _49408_ (_16942_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nand _49409_ (_16943_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  nand _49410_ (_16944_, _16943_, _16942_);
  nand _49411_ (_16945_, _16944_, _06717_);
  nand _49412_ (_16946_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nand _49413_ (_16947_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nand _49414_ (_16948_, _16947_, _16946_);
  nand _49415_ (_16949_, _16948_, _06716_);
  nand _49416_ (_16950_, _16949_, _16945_);
  nand _49417_ (_16951_, _16950_, _06751_);
  nand _49418_ (_16952_, _16951_, _16941_);
  nand _49419_ (_16953_, _16952_, _06761_);
  nor _49420_ (_16954_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  nor _49421_ (_16955_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nor _49422_ (_16956_, _16955_, _16954_);
  nand _49423_ (_16957_, _16956_, _06717_);
  nor _49424_ (_16958_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  nor _49425_ (_16959_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  nor _49426_ (_16960_, _16959_, _16958_);
  nand _49427_ (_16961_, _16960_, _06716_);
  nand _49428_ (_16962_, _16961_, _16957_);
  nand _49429_ (_16963_, _16962_, _06748_);
  nor _49430_ (_16964_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  nor _49431_ (_16965_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nor _49432_ (_16966_, _16965_, _16964_);
  nand _49433_ (_16967_, _16966_, _06717_);
  nor _49434_ (_16968_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  nor _49435_ (_16969_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  nor _49436_ (_16970_, _16969_, _16968_);
  nand _49437_ (_16971_, _16970_, _06716_);
  nand _49438_ (_16972_, _16971_, _16967_);
  nand _49439_ (_16973_, _16972_, _06751_);
  nand _49440_ (_16974_, _16973_, _16963_);
  nand _49441_ (_16975_, _16974_, _06760_);
  nand _49442_ (_16976_, _16975_, _16953_);
  nand _49443_ (_16977_, _16976_, _06731_);
  nand _49444_ (_16978_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  nand _49445_ (_16979_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  nand _49446_ (_16980_, _16979_, _16978_);
  nand _49447_ (_16981_, _16980_, _06717_);
  nand _49448_ (_16982_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nand _49449_ (_16983_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nand _49450_ (_16984_, _16983_, _16982_);
  nand _49451_ (_16985_, _16984_, _06716_);
  nand _49452_ (_16986_, _16985_, _16981_);
  nand _49453_ (_16987_, _16986_, _06748_);
  nand _49454_ (_16988_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  nand _49455_ (_16989_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  nand _49456_ (_16990_, _16989_, _16988_);
  nand _49457_ (_16991_, _16990_, _06717_);
  nand _49458_ (_16992_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nand _49459_ (_16993_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  nand _49460_ (_16994_, _16993_, _16992_);
  nand _49461_ (_16995_, _16994_, _06716_);
  nand _49462_ (_16996_, _16995_, _16991_);
  nand _49463_ (_16997_, _16996_, _06751_);
  nand _49464_ (_16998_, _16997_, _16987_);
  nand _49465_ (_16999_, _16998_, _06761_);
  nor _49466_ (_17000_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  nor _49467_ (_17001_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  nor _49468_ (_17002_, _17001_, _17000_);
  nand _49469_ (_17003_, _17002_, _06717_);
  nor _49470_ (_17004_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nor _49471_ (_17005_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  nor _49472_ (_17006_, _17005_, _17004_);
  nand _49473_ (_17007_, _17006_, _06716_);
  nand _49474_ (_17008_, _17007_, _17003_);
  nand _49475_ (_17009_, _17008_, _06748_);
  nor _49476_ (_17010_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  nor _49477_ (_17011_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  nor _49478_ (_17012_, _17011_, _17010_);
  nand _49479_ (_17013_, _17012_, _06717_);
  nor _49480_ (_17014_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  nor _49481_ (_17015_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nor _49482_ (_17016_, _17015_, _17014_);
  nand _49483_ (_17017_, _17016_, _06716_);
  nand _49484_ (_17018_, _17017_, _17013_);
  nand _49485_ (_17019_, _17018_, _06751_);
  nand _49486_ (_17020_, _17019_, _17009_);
  nand _49487_ (_17021_, _17020_, _06760_);
  nand _49488_ (_17022_, _17021_, _16999_);
  nand _49489_ (_17023_, _17022_, _06780_);
  nand _49490_ (_17024_, _17023_, _16977_);
  nand _49491_ (_17025_, _17024_, _06733_);
  nand _49492_ (_17026_, _17025_, _16931_);
  nor _49493_ (_17027_, _17026_, _13106_);
  nor _49494_ (_17028_, _17027_, _16834_);
  nor _49495_ (_17029_, _17028_, _25843_);
  nor _49496_ (_17030_, _17029_, _16642_);
  nor _49497_ (_17031_, _17030_, _13105_);
  not _49498_ (_17032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nand _49499_ (_17033_, _13105_, _17032_);
  nand _49500_ (_17034_, _17033_, _26487_);
  nor _49501_ (_06736_, _17034_, _17031_);
  nand _49502_ (_17035_, _11783_, _24789_);
  nand _49503_ (_17036_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  nand _49504_ (_06742_, _17036_, _17035_);
  nand _49505_ (_17037_, _12260_, _24789_);
  nand _49506_ (_17038_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nand _49507_ (_06746_, _17038_, _17037_);
  nand _49508_ (_17039_, _11738_, _25099_);
  nand _49509_ (_17040_, _11741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  nand _49510_ (_06750_, _17040_, _17039_);
  nand _49511_ (_17041_, _12260_, _25150_);
  nand _49512_ (_17042_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nand _49513_ (_06752_, _17042_, _17041_);
  nand _49514_ (_17043_, _11862_, _25150_);
  nand _49515_ (_17044_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  nand _49516_ (_06754_, _17044_, _17043_);
  nand _49517_ (_17045_, _03894_, _25099_);
  nand _49518_ (_17046_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  nand _49519_ (_06757_, _17046_, _17045_);
  nor _49520_ (_17047_, _07942_, _25680_);
  not _49521_ (_17048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  not _49522_ (_17049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _49523_ (_17050_, _07960_, _17049_);
  not _49524_ (_17051_, _17050_);
  nor _49525_ (_17052_, _17051_, _17048_);
  nand _49526_ (_17053_, _17052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  not _49527_ (_17054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  not _49528_ (_17055_, _17052_);
  nand _49529_ (_17056_, _17055_, _17054_);
  nand _49530_ (_17057_, _17056_, _17053_);
  nor _49531_ (_17058_, _07664_, _05826_);
  nor _49532_ (_17059_, _17058_, _07948_);
  not _49533_ (_17060_, _17059_);
  nor _49534_ (_17061_, _17060_, _17057_);
  nand _49535_ (_17062_, _17060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  not _49536_ (_17063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _49537_ (_17064_, _07980_, _07945_);
  nor _49538_ (_17065_, _17064_, _17063_);
  nand _49539_ (_17066_, _17065_, _07983_);
  nand _49540_ (_17067_, _17066_, _17062_);
  nor _49541_ (_17068_, _17067_, _17061_);
  nand _49542_ (_17069_, _17068_, _07942_);
  nand _49543_ (_17070_, _17069_, _26487_);
  nor _49544_ (_06762_, _17070_, _17047_);
  nor _49545_ (_17071_, _04175_, _25194_);
  nor _49546_ (_17072_, _07562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _49547_ (_17073_, _17072_, _07564_);
  nor _49548_ (_17074_, _07637_, _04181_);
  nor _49549_ (_17075_, _17074_, _17073_);
  nor _49550_ (_17076_, _17075_, _01644_);
  nor _49551_ (_17077_, _01642_, _01589_);
  nor _49552_ (_17078_, _17077_, _17076_);
  nand _49553_ (_17079_, _17078_, _04175_);
  nand _49554_ (_17080_, _17079_, _26487_);
  nor _49555_ (_06782_, _17080_, _17071_);
  nand _49556_ (_17081_, _11931_, _24927_);
  nand _49557_ (_17082_, _11933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  nand _49558_ (_06785_, _17082_, _17081_);
  nand _49559_ (_17083_, _11973_, _25203_);
  nand _49560_ (_17084_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nand _49561_ (_06789_, _17084_, _17083_);
  nor _49562_ (_17085_, _04173_, _25089_);
  nor _49563_ (_17086_, _01635_, _04183_);
  not _49564_ (_17087_, _01635_);
  nor _49565_ (_17088_, _17087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _49566_ (_17089_, _17088_, _17086_);
  nor _49567_ (_17090_, _17089_, _01616_);
  not _49568_ (_17091_, _01606_);
  nand _49569_ (_17092_, _17091_, _04183_);
  nor _49570_ (_17093_, _07530_, _07747_);
  nand _49571_ (_17094_, _17093_, _17092_);
  not _49572_ (_17095_, _01598_);
  nand _49573_ (_17096_, _17095_, _04183_);
  nor _49574_ (_17097_, _07537_, _04208_);
  nand _49575_ (_17098_, _17097_, _17096_);
  nand _49576_ (_17099_, _17098_, _17094_);
  nor _49577_ (_17100_, _17099_, _17090_);
  nand _49578_ (_17101_, _17100_, _04173_);
  nand _49579_ (_17102_, _17101_, _04175_);
  nor _49580_ (_17103_, _17102_, _17085_);
  nor _49581_ (_17104_, _04175_, _04183_);
  nor _49582_ (_17105_, _17104_, _17103_);
  nor _49583_ (_06791_, _17105_, rst);
  nand _49584_ (_17106_, _11783_, _28096_);
  nand _49585_ (_17107_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  nand _49586_ (_06799_, _17107_, _17106_);
  nand _49587_ (_17108_, _12976_, _25099_);
  nand _49588_ (_17109_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nand _49589_ (_06803_, _17109_, _17108_);
  nand _49590_ (_17110_, _11772_, _28096_);
  nand _49591_ (_17111_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  nand _49592_ (_06805_, _17111_, _17110_);
  nor _49593_ (_17112_, _05824_, _25139_);
  not _49594_ (_17113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nand _49595_ (_17114_, _05824_, _17113_);
  nand _49596_ (_17115_, _17114_, _26487_);
  nor _49597_ (_06806_, _17115_, _17112_);
  nand _49598_ (_17116_, _12038_, _24830_);
  nand _49599_ (_17117_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nand _49600_ (_06811_, _17117_, _17116_);
  nand _49601_ (_17118_, _11783_, _25099_);
  nand _49602_ (_17119_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  nand _49603_ (_06812_, _17119_, _17118_);
  nand _49604_ (_17120_, _11772_, _25150_);
  nand _49605_ (_17121_, _11776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  nand _49606_ (_06813_, _17121_, _17120_);
  nand _49607_ (_17122_, _12976_, _24830_);
  nand _49608_ (_17123_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  nand _49609_ (_06815_, _17123_, _17122_);
  nand _49610_ (_17124_, _11783_, _25203_);
  nand _49611_ (_17125_, _11785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nand _49612_ (_06817_, _17125_, _17124_);
  nor _49613_ (_06819_, _00536_, _27980_);
  nand _49614_ (_17126_, _12038_, _24789_);
  nand _49615_ (_17127_, _12040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  nand _49616_ (_06824_, _17127_, _17126_);
  nand _49617_ (_17128_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  nand _49618_ (_17129_, _10084_, _25150_);
  nand _49619_ (_06831_, _17129_, _17128_);
  nand _49620_ (_17130_, _11973_, _24789_);
  nand _49621_ (_17131_, _11975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nand _49622_ (_06832_, _17131_, _17130_);
  nand _49623_ (_17132_, _13056_, _24830_);
  nand _49624_ (_17133_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nand _49625_ (_06841_, _17133_, _17132_);
  nand _49626_ (_17134_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  nand _49627_ (_17135_, _10084_, _24927_);
  nand _49628_ (_06866_, _17135_, _17134_);
  nor _49629_ (_17136_, _07818_, _00954_);
  nand _49630_ (_17137_, _17136_, _24789_);
  not _49631_ (_17138_, _17136_);
  nand _49632_ (_17139_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nand _49633_ (_06870_, _17139_, _17137_);
  nand _49634_ (_17140_, _17136_, _25150_);
  nand _49635_ (_17141_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nand _49636_ (_06874_, _17141_, _17140_);
  nand _49637_ (_17142_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  nand _49638_ (_17143_, _10084_, _25039_);
  nand _49639_ (_06884_, _17143_, _17142_);
  nand _49640_ (_17144_, _12260_, _24927_);
  nand _49641_ (_17145_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  nand _49642_ (_06887_, _17145_, _17144_);
  nand _49643_ (_17146_, _11862_, _24830_);
  nand _49644_ (_17147_, _11864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nand _49645_ (_06890_, _17147_, _17146_);
  nand _49646_ (_17148_, _12260_, _25203_);
  nand _49647_ (_17149_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  nand _49648_ (_06901_, _17149_, _17148_);
  nand _49649_ (_17150_, _13056_, _25203_);
  nand _49650_ (_17151_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  nand _49651_ (_06903_, _17151_, _17150_);
  nand _49652_ (_17152_, _13056_, _28096_);
  nand _49653_ (_17153_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nand _49654_ (_06908_, _17153_, _17152_);
  nand _49655_ (_17154_, _12260_, _25039_);
  nand _49656_ (_17155_, _12262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  nand _49657_ (_06911_, _17155_, _17154_);
  nand _49658_ (_17156_, _12235_, _28096_);
  nand _49659_ (_17157_, _12237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  nand _49660_ (_06918_, _17157_, _17156_);
  nand _49661_ (_17158_, _13056_, _25099_);
  nand _49662_ (_17159_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  nand _49663_ (_06927_, _17159_, _17158_);
  nand _49664_ (_17160_, _08168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  nand _49665_ (_17161_, _08167_, _24830_);
  nand _49666_ (_06933_, _17161_, _17160_);
  nand _49667_ (_17162_, _11919_, _24830_);
  nand _49668_ (_17163_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  nand _49669_ (_06940_, _17163_, _17162_);
  nand _49670_ (_17164_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  nand _49671_ (_17165_, _10084_, _24789_);
  nand _49672_ (_06942_, _17165_, _17164_);
  nand _49673_ (_17166_, _17136_, _25099_);
  nand _49674_ (_17167_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  nand _49675_ (_06949_, _17167_, _17166_);
  nand _49676_ (_17168_, _17136_, _24830_);
  nand _49677_ (_17169_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  nand _49678_ (_06954_, _17169_, _17168_);
  nand _49679_ (_17170_, _03442_, _24789_);
  nand _49680_ (_17171_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  nand _49681_ (_06956_, _17171_, _17170_);
  nand _49682_ (_17172_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  nand _49683_ (_17173_, _12698_, _24927_);
  nand _49684_ (_06961_, _17173_, _17172_);
  nand _49685_ (_17174_, _00979_, _25203_);
  nand _49686_ (_17175_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  nand _49687_ (_06963_, _17175_, _17174_);
  nand _49688_ (_17176_, _00479_, _24789_);
  nand _49689_ (_17177_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  nand _49690_ (_06965_, _17177_, _17176_);
  nand _49691_ (_17178_, _08354_, _24830_);
  nand _49692_ (_17179_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  nand _49693_ (_06987_, _17179_, _17178_);
  nand _49694_ (_17180_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  nand _49695_ (_17181_, _12698_, _25099_);
  nand _49696_ (_06991_, _17181_, _17180_);
  nand _49697_ (_17182_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  nand _49698_ (_17183_, _12671_, _25150_);
  nand _49699_ (_06996_, _17183_, _17182_);
  nand _49700_ (_17184_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  nand _49701_ (_17185_, _12671_, _24830_);
  nand _49702_ (_07002_, _17185_, _17184_);
  nand _49703_ (_17186_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  nand _49704_ (_17187_, _12642_, _24927_);
  nand _49705_ (_07008_, _17187_, _17186_);
  nand _49706_ (_17188_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  nand _49707_ (_17189_, _12642_, _25099_);
  nand _49708_ (_07016_, _17189_, _17188_);
  nand _49709_ (_17190_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  nand _49710_ (_17191_, _08212_, _24789_);
  nand _49711_ (_07018_, _17191_, _17190_);
  nand _49712_ (_17192_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nand _49713_ (_17193_, _12618_, _25150_);
  nand _49714_ (_07021_, _17193_, _17192_);
  nand _49715_ (_17194_, _28059_, _24927_);
  nand _49716_ (_17195_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  nand _49717_ (_07024_, _17195_, _17194_);
  nand _49718_ (_17196_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  nand _49719_ (_17197_, _08212_, _25150_);
  nand _49720_ (_07026_, _17197_, _17196_);
  nand _49721_ (_17198_, _17136_, _25039_);
  nand _49722_ (_17199_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nand _49723_ (_07028_, _17199_, _17198_);
  nand _49724_ (_17200_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  nand _49725_ (_17201_, _12618_, _25203_);
  nand _49726_ (_07031_, _17201_, _17200_);
  nand _49727_ (_17202_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nand _49728_ (_17203_, _12590_, _25039_);
  nand _49729_ (_07041_, _17203_, _17202_);
  nand _49730_ (_17204_, _17136_, _25203_);
  nand _49731_ (_17205_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nand _49732_ (_07043_, _17205_, _17204_);
  nand _49733_ (_17206_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nand _49734_ (_17207_, _12590_, _25099_);
  nand _49735_ (_07047_, _17207_, _17206_);
  nand _49736_ (_17208_, _17136_, _28096_);
  nand _49737_ (_17209_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  nand _49738_ (_07049_, _17209_, _17208_);
  nand _49739_ (_17210_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  nand _49740_ (_17211_, _12566_, _25150_);
  nand _49741_ (_07052_, _17211_, _17210_);
  nand _49742_ (_17212_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  nand _49743_ (_17213_, _12566_, _25099_);
  nand _49744_ (_07061_, _17213_, _17212_);
  nand _49745_ (_17214_, _12413_, _25150_);
  nand _49746_ (_17215_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nand _49747_ (_07067_, _17215_, _17214_);
  nand _49748_ (_17216_, _12413_, _25039_);
  nand _49749_ (_17217_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  nand _49750_ (_07070_, _17217_, _17216_);
  nand _49751_ (_17218_, _12522_, _25150_);
  nand _49752_ (_17219_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nand _49753_ (_07074_, _17219_, _17218_);
  nor _49754_ (_17220_, _07818_, _00393_);
  nand _49755_ (_17221_, _17220_, _28096_);
  not _49756_ (_17222_, _17220_);
  nand _49757_ (_17223_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  nand _49758_ (_07078_, _17223_, _17221_);
  nand _49759_ (_17224_, _12522_, _25039_);
  nand _49760_ (_17225_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  nand _49761_ (_07081_, _17225_, _17224_);
  nand _49762_ (_17226_, _12522_, _24830_);
  nand _49763_ (_17227_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nand _49764_ (_07085_, _17227_, _17226_);
  nand _49765_ (_17228_, _12498_, _24789_);
  nand _49766_ (_17229_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nand _49767_ (_07087_, _17229_, _17228_);
  nand _49768_ (_17230_, _12498_, _24927_);
  nand _49769_ (_17231_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  nand _49770_ (_07089_, _17231_, _17230_);
  nand _49771_ (_17232_, _17220_, _25099_);
  nand _49772_ (_17233_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nand _49773_ (_07092_, _17233_, _17232_);
  nand _49774_ (_17234_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nand _49775_ (_17235_, _10084_, _28096_);
  nand _49776_ (_07094_, _17235_, _17234_);
  nand _49777_ (_17236_, _12498_, _25099_);
  nand _49778_ (_17237_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  nand _49779_ (_07099_, _17237_, _17236_);
  nand _49780_ (_17238_, _12483_, _25150_);
  nand _49781_ (_17239_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  nand _49782_ (_07120_, _17239_, _17238_);
  nand _49783_ (_17240_, _10085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  nand _49784_ (_17241_, _10084_, _25099_);
  nand _49785_ (_07125_, _17241_, _17240_);
  nand _49786_ (_17242_, _12483_, _28096_);
  nand _49787_ (_17243_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nand _49788_ (_07128_, _17243_, _17242_);
  nand _49789_ (_17244_, _07819_, _24789_);
  nand _49790_ (_17245_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  nand _49791_ (_07131_, _17245_, _17244_);
  nand _49792_ (_17246_, _17220_, _25203_);
  nand _49793_ (_17247_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  nand _49794_ (_07133_, _17247_, _17246_);
  nand _49795_ (_17248_, _12465_, _28096_);
  nand _49796_ (_17249_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  nand _49797_ (_07137_, _17249_, _17248_);
  nand _49798_ (_17250_, _05848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  nand _49799_ (_17251_, _05847_, _24830_);
  nand _49800_ (_07140_, _17251_, _17250_);
  nand _49801_ (_17252_, _17220_, _24927_);
  nand _49802_ (_17253_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  nand _49803_ (_07143_, _17253_, _17252_);
  nand _49804_ (_17254_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nand _49805_ (_17255_, _12671_, _28096_);
  nand _49806_ (_07147_, _17255_, _17254_);
  nand _49807_ (_17256_, _17220_, _25039_);
  nand _49808_ (_17257_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  nand _49809_ (_07149_, _17257_, _17256_);
  nand _49810_ (_17258_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  nand _49811_ (_17259_, _12642_, _24789_);
  nand _49812_ (_07151_, _17259_, _17258_);
  nand _49813_ (_17260_, _12643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nand _49814_ (_17261_, _12642_, _25203_);
  nand _49815_ (_07154_, _17261_, _17260_);
  nand _49816_ (_17262_, _11919_, _28096_);
  nand _49817_ (_17263_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  nand _49818_ (_07158_, _17263_, _17262_);
  nand _49819_ (_17264_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nand _49820_ (_17265_, _08212_, _24830_);
  nand _49821_ (_28311_, _17265_, _17264_);
  nand _49822_ (_17266_, _11919_, _25039_);
  nand _49823_ (_17267_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  nand _49824_ (_07161_, _17267_, _17266_);
  nand _49825_ (_17268_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  nand _49826_ (_17269_, _12618_, _24830_);
  nand _49827_ (_07165_, _17269_, _17268_);
  nand _49828_ (_17270_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  nand _49829_ (_17271_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  nand _49830_ (_17273_, _17271_, _17270_);
  nand _49831_ (_17274_, _17273_, _06717_);
  nand _49832_ (_17275_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  nand _49833_ (_17276_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  nand _49834_ (_17277_, _17276_, _17275_);
  nand _49835_ (_17278_, _17277_, _06716_);
  nand _49836_ (_17279_, _17278_, _17274_);
  nand _49837_ (_17280_, _17279_, _06748_);
  nand _49838_ (_17281_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  nand _49839_ (_17282_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  nand _49840_ (_17284_, _17282_, _17281_);
  nand _49841_ (_17285_, _17284_, _06717_);
  nand _49842_ (_17286_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  nand _49843_ (_17287_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  nand _49844_ (_17288_, _17287_, _17286_);
  nand _49845_ (_17289_, _17288_, _06716_);
  nand _49846_ (_17290_, _17289_, _17285_);
  nand _49847_ (_17291_, _17290_, _06751_);
  nand _49848_ (_17292_, _17291_, _17280_);
  nand _49849_ (_17293_, _17292_, _06761_);
  nor _49850_ (_17294_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  nor _49851_ (_17295_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  nor _49852_ (_17296_, _17295_, _17294_);
  nand _49853_ (_17297_, _17296_, _06716_);
  nand _49854_ (_17298_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  nand _49855_ (_17299_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  nand _49856_ (_17300_, _17299_, _17298_);
  nand _49857_ (_17301_, _17300_, _06717_);
  nand _49858_ (_17302_, _17301_, _17297_);
  nand _49859_ (_17303_, _17302_, _06748_);
  nor _49860_ (_17304_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  nor _49861_ (_17305_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  nor _49862_ (_17306_, _17305_, _17304_);
  nand _49863_ (_17307_, _17306_, _06716_);
  nand _49864_ (_17308_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  nand _49865_ (_17309_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  nand _49866_ (_17310_, _17309_, _17308_);
  nand _49867_ (_17311_, _17310_, _06717_);
  nand _49868_ (_17312_, _17311_, _17307_);
  nand _49869_ (_17313_, _17312_, _06751_);
  nand _49870_ (_17314_, _17313_, _17303_);
  nand _49871_ (_17315_, _17314_, _06760_);
  nand _49872_ (_17316_, _17315_, _17293_);
  nand _49873_ (_17317_, _17316_, _06780_);
  nand _49874_ (_17318_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  nand _49875_ (_17319_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  nand _49876_ (_17320_, _17319_, _17318_);
  nand _49877_ (_17321_, _17320_, _06717_);
  nand _49878_ (_17322_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  nand _49879_ (_17323_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  nand _49880_ (_17324_, _17323_, _17322_);
  nand _49881_ (_17325_, _17324_, _06716_);
  nand _49882_ (_17326_, _17325_, _17321_);
  nand _49883_ (_17327_, _17326_, _06748_);
  nand _49884_ (_17328_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  nand _49885_ (_17329_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  nand _49886_ (_17330_, _17329_, _17328_);
  nand _49887_ (_17331_, _17330_, _06717_);
  nand _49888_ (_17332_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  nand _49889_ (_17333_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  nand _49890_ (_17334_, _17333_, _17332_);
  nand _49891_ (_17335_, _17334_, _06716_);
  nand _49892_ (_17336_, _17335_, _17331_);
  nand _49893_ (_17337_, _17336_, _06751_);
  nand _49894_ (_17338_, _17337_, _17327_);
  nand _49895_ (_17339_, _17338_, _06761_);
  nor _49896_ (_17340_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  nor _49897_ (_17341_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  nor _49898_ (_17342_, _17341_, _17340_);
  nand _49899_ (_17343_, _17342_, _06717_);
  nor _49900_ (_17345_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  nor _49901_ (_17346_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  nor _49902_ (_17347_, _17346_, _17345_);
  nand _49903_ (_17348_, _17347_, _06716_);
  nand _49904_ (_17349_, _17348_, _17343_);
  nand _49905_ (_17350_, _17349_, _06748_);
  nor _49906_ (_17351_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  nor _49907_ (_17352_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  nor _49908_ (_17353_, _17352_, _17351_);
  nand _49909_ (_17354_, _17353_, _06717_);
  nor _49910_ (_17355_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  nor _49911_ (_17356_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nor _49912_ (_17357_, _17356_, _17355_);
  nand _49913_ (_17358_, _17357_, _06716_);
  nand _49914_ (_17359_, _17358_, _17354_);
  nand _49915_ (_17360_, _17359_, _06751_);
  nand _49916_ (_17361_, _17360_, _17350_);
  nand _49917_ (_17362_, _17361_, _06760_);
  nand _49918_ (_17363_, _17362_, _17339_);
  nand _49919_ (_17364_, _17363_, _06731_);
  nand _49920_ (_17365_, _17364_, _17317_);
  nand _49921_ (_17366_, _17365_, _06734_);
  nand _49922_ (_17367_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand _49923_ (_17368_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand _49924_ (_17369_, _17368_, _17367_);
  nand _49925_ (_17370_, _17369_, _06717_);
  nand _49926_ (_17371_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nand _49927_ (_17372_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nand _49928_ (_17373_, _17372_, _17371_);
  nand _49929_ (_17374_, _17373_, _06716_);
  nand _49930_ (_17375_, _17374_, _17370_);
  nand _49931_ (_17376_, _17375_, _06748_);
  nand _49932_ (_17377_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand _49933_ (_17378_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand _49934_ (_17379_, _17378_, _17377_);
  nand _49935_ (_17380_, _17379_, _06717_);
  nand _49936_ (_17381_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nand _49937_ (_17382_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nand _49938_ (_17383_, _17382_, _17381_);
  nand _49939_ (_17384_, _17383_, _06716_);
  nand _49940_ (_17385_, _17384_, _17380_);
  nand _49941_ (_17386_, _17385_, _06751_);
  nand _49942_ (_17387_, _17386_, _17376_);
  nand _49943_ (_17388_, _17387_, _06761_);
  nor _49944_ (_17389_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor _49945_ (_17390_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _49946_ (_17391_, _17390_, _17389_);
  nand _49947_ (_17392_, _17391_, _06716_);
  nand _49948_ (_17393_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand _49949_ (_17394_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand _49950_ (_17395_, _17394_, _17393_);
  nand _49951_ (_17396_, _17395_, _06717_);
  nand _49952_ (_17397_, _17396_, _17392_);
  nand _49953_ (_17398_, _17397_, _06748_);
  nor _49954_ (_17399_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nor _49955_ (_17400_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor _49956_ (_17401_, _17400_, _17399_);
  nand _49957_ (_17402_, _17401_, _06716_);
  nand _49958_ (_17403_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand _49959_ (_17404_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand _49960_ (_17405_, _17404_, _17403_);
  nand _49961_ (_17406_, _17405_, _06717_);
  nand _49962_ (_17407_, _17406_, _17402_);
  nand _49963_ (_17408_, _17407_, _06751_);
  nand _49964_ (_17409_, _17408_, _17398_);
  nand _49965_ (_17410_, _17409_, _06760_);
  nand _49966_ (_17411_, _17410_, _17388_);
  nand _49967_ (_17412_, _17411_, _06780_);
  nand _49968_ (_17413_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  nand _49969_ (_17414_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  nand _49970_ (_17415_, _17414_, _17413_);
  nand _49971_ (_17416_, _17415_, _06717_);
  nand _49972_ (_17417_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  nand _49973_ (_17418_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  nand _49974_ (_17419_, _17418_, _17417_);
  nand _49975_ (_17420_, _17419_, _06716_);
  nand _49976_ (_17421_, _17420_, _17416_);
  nand _49977_ (_17422_, _17421_, _06748_);
  nand _49978_ (_17423_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  nand _49979_ (_17424_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  nand _49980_ (_17425_, _17424_, _17423_);
  nand _49981_ (_17426_, _17425_, _06717_);
  nand _49982_ (_17427_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  nand _49983_ (_17428_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  nand _49984_ (_17429_, _17428_, _17427_);
  nand _49985_ (_17430_, _17429_, _06716_);
  nand _49986_ (_17431_, _17430_, _17426_);
  nand _49987_ (_17432_, _17431_, _06751_);
  nand _49988_ (_17433_, _17432_, _17422_);
  nand _49989_ (_17434_, _17433_, _06761_);
  not _49990_ (_17435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  nand _49991_ (_17436_, _06774_, _17435_);
  nor _49992_ (_17437_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  nor _49993_ (_17438_, _17437_, _06716_);
  nand _49994_ (_17439_, _17438_, _17436_);
  nor _49995_ (_17440_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  nor _49996_ (_17441_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  nor _49997_ (_17442_, _17441_, _17440_);
  nand _49998_ (_17443_, _17442_, _06716_);
  nand _49999_ (_17444_, _17443_, _17439_);
  nand _50000_ (_17445_, _17444_, _06748_);
  nor _50001_ (_17446_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  nor _50002_ (_17447_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  nor _50003_ (_17448_, _17447_, _17446_);
  nand _50004_ (_17449_, _17448_, _06717_);
  nor _50005_ (_17450_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nor _50006_ (_17451_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  nor _50007_ (_17452_, _17451_, _17450_);
  nand _50008_ (_17453_, _17452_, _06716_);
  nand _50009_ (_17454_, _17453_, _17449_);
  nand _50010_ (_17455_, _17454_, _06751_);
  nand _50011_ (_17456_, _17455_, _17445_);
  nand _50012_ (_17457_, _17456_, _06760_);
  nand _50013_ (_17458_, _17457_, _17434_);
  nand _50014_ (_17459_, _17458_, _06731_);
  nand _50015_ (_17460_, _17459_, _17412_);
  nand _50016_ (_17461_, _17460_, _06733_);
  nand _50017_ (_17462_, _17461_, _17366_);
  nor _50018_ (_17463_, _17462_, _06723_);
  nand _50019_ (_17464_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  nand _50020_ (_17465_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  nand _50021_ (_17466_, _17465_, _17464_);
  nand _50022_ (_17467_, _17466_, _06717_);
  nand _50023_ (_17468_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  nand _50024_ (_17469_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  nand _50025_ (_17470_, _17469_, _17468_);
  nand _50026_ (_17471_, _17470_, _06716_);
  nand _50027_ (_17472_, _17471_, _17467_);
  nand _50028_ (_17473_, _17472_, _06748_);
  nand _50029_ (_17474_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  nand _50030_ (_17476_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  nand _50031_ (_17477_, _17476_, _17474_);
  nand _50032_ (_17478_, _17477_, _06717_);
  nand _50033_ (_17479_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  nand _50034_ (_17480_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  nand _50035_ (_17481_, _17480_, _17479_);
  nand _50036_ (_17482_, _17481_, _06716_);
  nand _50037_ (_17483_, _17482_, _17478_);
  nand _50038_ (_17484_, _17483_, _06751_);
  nand _50039_ (_17485_, _17484_, _17473_);
  nand _50040_ (_17486_, _17485_, _06761_);
  nor _50041_ (_17487_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  nor _50042_ (_17488_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  nor _50043_ (_17489_, _17488_, _17487_);
  nand _50044_ (_17490_, _17489_, _06717_);
  nor _50045_ (_17491_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  nor _50046_ (_17492_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  nor _50047_ (_17493_, _17492_, _17491_);
  nand _50048_ (_17494_, _17493_, _06716_);
  nand _50049_ (_17495_, _17494_, _17490_);
  nand _50050_ (_17496_, _17495_, _06748_);
  not _50051_ (_17497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  nand _50052_ (_17498_, _06774_, _17497_);
  nor _50053_ (_17499_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  nor _50054_ (_17500_, _17499_, _06716_);
  nand _50055_ (_17501_, _17500_, _17498_);
  nor _50056_ (_17502_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  nor _50057_ (_17503_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  nor _50058_ (_17504_, _17503_, _17502_);
  nand _50059_ (_17505_, _17504_, _06716_);
  nand _50060_ (_17506_, _17505_, _17501_);
  nand _50061_ (_17507_, _17506_, _06751_);
  nand _50062_ (_17508_, _17507_, _17496_);
  nand _50063_ (_17509_, _17508_, _06760_);
  nand _50064_ (_17510_, _17509_, _17486_);
  nand _50065_ (_17511_, _17510_, _06780_);
  nand _50066_ (_17512_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  nand _50067_ (_17513_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  nand _50068_ (_17514_, _17513_, _17512_);
  nand _50069_ (_17515_, _17514_, _06717_);
  nand _50070_ (_17516_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  nand _50071_ (_17517_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  nand _50072_ (_17518_, _17517_, _17516_);
  nand _50073_ (_17519_, _17518_, _06716_);
  nand _50074_ (_17520_, _17519_, _17515_);
  nand _50075_ (_17521_, _17520_, _06748_);
  nand _50076_ (_17522_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  nand _50077_ (_17523_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  nand _50078_ (_17524_, _17523_, _17522_);
  nand _50079_ (_17525_, _17524_, _06717_);
  nand _50080_ (_17526_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  nand _50081_ (_17527_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  nand _50082_ (_17528_, _17527_, _17526_);
  nand _50083_ (_17529_, _17528_, _06716_);
  nand _50084_ (_17530_, _17529_, _17525_);
  nand _50085_ (_17531_, _17530_, _06751_);
  nand _50086_ (_17532_, _17531_, _17521_);
  nand _50087_ (_17533_, _17532_, _06761_);
  not _50088_ (_17534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  nand _50089_ (_17535_, _06774_, _17534_);
  nor _50090_ (_17536_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nor _50091_ (_17537_, _17536_, _06716_);
  nand _50092_ (_17538_, _17537_, _17535_);
  nor _50093_ (_17539_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  nor _50094_ (_17540_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  nor _50095_ (_17541_, _17540_, _17539_);
  nand _50096_ (_17542_, _17541_, _06716_);
  nand _50097_ (_17543_, _17542_, _17538_);
  nand _50098_ (_17544_, _17543_, _06748_);
  nor _50099_ (_17545_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nor _50100_ (_17546_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  nor _50101_ (_17547_, _17546_, _17545_);
  nand _50102_ (_17548_, _17547_, _06717_);
  nor _50103_ (_17549_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  nor _50104_ (_17550_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  nor _50105_ (_17551_, _17550_, _17549_);
  nand _50106_ (_17552_, _17551_, _06716_);
  nand _50107_ (_17553_, _17552_, _17548_);
  nand _50108_ (_17554_, _17553_, _06751_);
  nand _50109_ (_17555_, _17554_, _17544_);
  nand _50110_ (_17556_, _17555_, _06760_);
  nand _50111_ (_17557_, _17556_, _17533_);
  nand _50112_ (_17558_, _17557_, _06731_);
  nand _50113_ (_17559_, _17558_, _17511_);
  nand _50114_ (_17560_, _17559_, _06733_);
  nand _50115_ (_17561_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  nand _50116_ (_17562_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nand _50117_ (_17563_, _17562_, _17561_);
  nand _50118_ (_17564_, _17563_, _06716_);
  nand _50119_ (_17565_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  nand _50120_ (_17566_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  nand _50121_ (_17567_, _17566_, _17565_);
  nand _50122_ (_17568_, _17567_, _06717_);
  nand _50123_ (_17569_, _17568_, _17564_);
  nand _50124_ (_17570_, _17569_, _06748_);
  nand _50125_ (_17571_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  nand _50126_ (_17572_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  nand _50127_ (_17573_, _17572_, _17571_);
  nand _50128_ (_17574_, _17573_, _06716_);
  nand _50129_ (_17575_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  nand _50130_ (_17576_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  nand _50131_ (_17577_, _17576_, _17575_);
  nand _50132_ (_17578_, _17577_, _06717_);
  nand _50133_ (_17579_, _17578_, _17574_);
  nand _50134_ (_17580_, _17579_, _06751_);
  nand _50135_ (_17581_, _17580_, _17570_);
  nand _50136_ (_17582_, _17581_, _06761_);
  nand _50137_ (_17583_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  nand _50138_ (_17584_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  nand _50139_ (_17585_, _17584_, _17583_);
  nand _50140_ (_17586_, _17585_, _06717_);
  nor _50141_ (_17587_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  nor _50142_ (_17588_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  nor _50143_ (_17589_, _17588_, _17587_);
  nand _50144_ (_17590_, _17589_, _06716_);
  nand _50145_ (_17591_, _17590_, _17586_);
  nand _50146_ (_17592_, _17591_, _06748_);
  nand _50147_ (_17593_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  nand _50148_ (_17594_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  nand _50149_ (_17595_, _17594_, _17593_);
  nand _50150_ (_17596_, _17595_, _06717_);
  nor _50151_ (_17597_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  nor _50152_ (_17598_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  nor _50153_ (_17599_, _17598_, _17597_);
  nand _50154_ (_17600_, _17599_, _06716_);
  nand _50155_ (_17601_, _17600_, _17596_);
  nand _50156_ (_17602_, _17601_, _06751_);
  nand _50157_ (_17603_, _17602_, _17592_);
  nand _50158_ (_17604_, _17603_, _06760_);
  nand _50159_ (_17605_, _17604_, _17582_);
  nand _50160_ (_17606_, _17605_, _06780_);
  nand _50161_ (_17607_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  nand _50162_ (_17608_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nand _50163_ (_17609_, _17608_, _17607_);
  nand _50164_ (_17610_, _17609_, _06717_);
  nand _50165_ (_17611_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  nand _50166_ (_17612_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  nand _50167_ (_17613_, _17612_, _17611_);
  nand _50168_ (_17614_, _17613_, _06716_);
  nand _50169_ (_17615_, _17614_, _17610_);
  nand _50170_ (_17616_, _17615_, _06748_);
  nand _50171_ (_17617_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  nand _50172_ (_17618_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  nand _50173_ (_17619_, _17618_, _17617_);
  nand _50174_ (_17620_, _17619_, _06717_);
  nand _50175_ (_17621_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  nand _50176_ (_17622_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  nand _50177_ (_17623_, _17622_, _17621_);
  nand _50178_ (_17624_, _17623_, _06716_);
  nand _50179_ (_17625_, _17624_, _17620_);
  nand _50180_ (_17626_, _17625_, _06751_);
  nand _50181_ (_17627_, _17626_, _17616_);
  nand _50182_ (_17628_, _17627_, _06761_);
  nor _50183_ (_17629_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  nor _50184_ (_17630_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  nor _50185_ (_17631_, _17630_, _17629_);
  nand _50186_ (_17632_, _17631_, _06717_);
  nor _50187_ (_17633_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  nor _50188_ (_17634_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  nor _50189_ (_17635_, _17634_, _17633_);
  nand _50190_ (_17636_, _17635_, _06716_);
  nand _50191_ (_17637_, _17636_, _17632_);
  nand _50192_ (_17638_, _17637_, _06748_);
  nor _50193_ (_17639_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  nor _50194_ (_17640_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  nor _50195_ (_17641_, _17640_, _17639_);
  nor _50196_ (_17642_, _17641_, _06716_);
  nor _50197_ (_17643_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  nor _50198_ (_17644_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  nor _50199_ (_17645_, _17644_, _17643_);
  nor _50200_ (_17646_, _17645_, _06717_);
  nor _50201_ (_17647_, _17646_, _17642_);
  nand _50202_ (_17648_, _17647_, _06751_);
  nand _50203_ (_17649_, _17648_, _17638_);
  nand _50204_ (_17650_, _17649_, _06760_);
  nand _50205_ (_17651_, _17650_, _17628_);
  nand _50206_ (_17652_, _17651_, _06731_);
  nand _50207_ (_17653_, _17652_, _17606_);
  nand _50208_ (_17654_, _17653_, _06734_);
  nand _50209_ (_17655_, _17654_, _17560_);
  nor _50210_ (_17656_, _17655_, _13106_);
  nor _50211_ (_17657_, _17656_, _17463_);
  nor _50212_ (_17658_, _17657_, _25929_);
  nand _50213_ (_17659_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  nand _50214_ (_17660_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  nand _50215_ (_17661_, _17660_, _17659_);
  nand _50216_ (_17662_, _17661_, _06717_);
  nand _50217_ (_17663_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  nand _50218_ (_17664_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  nand _50219_ (_17665_, _17664_, _17663_);
  nand _50220_ (_17666_, _17665_, _06716_);
  nand _50221_ (_17667_, _17666_, _17662_);
  nand _50222_ (_17668_, _17667_, _06748_);
  nand _50223_ (_17669_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  nand _50224_ (_17670_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  nand _50225_ (_17671_, _17670_, _17669_);
  nand _50226_ (_17672_, _17671_, _06717_);
  nand _50227_ (_17673_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  nand _50228_ (_17674_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  nand _50229_ (_17675_, _17674_, _17673_);
  nand _50230_ (_17676_, _17675_, _06716_);
  nand _50231_ (_17677_, _17676_, _17672_);
  nand _50232_ (_17678_, _17677_, _06751_);
  nand _50233_ (_17679_, _17678_, _17668_);
  nand _50234_ (_17680_, _17679_, _06761_);
  nor _50235_ (_17681_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  nor _50236_ (_17682_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  nor _50237_ (_17683_, _17682_, _17681_);
  nand _50238_ (_17684_, _17683_, _06717_);
  nor _50239_ (_17685_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  nor _50240_ (_17686_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  nor _50241_ (_17687_, _17686_, _17685_);
  nand _50242_ (_17688_, _17687_, _06716_);
  nand _50243_ (_17689_, _17688_, _17684_);
  nand _50244_ (_17690_, _17689_, _06748_);
  nor _50245_ (_17691_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  nor _50246_ (_17692_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  nor _50247_ (_17693_, _17692_, _17691_);
  nand _50248_ (_17694_, _17693_, _06717_);
  nor _50249_ (_17695_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  nor _50250_ (_17696_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  nor _50251_ (_17697_, _17696_, _17695_);
  nand _50252_ (_17698_, _17697_, _06716_);
  nand _50253_ (_17699_, _17698_, _17694_);
  nand _50254_ (_17700_, _17699_, _06751_);
  nand _50255_ (_17701_, _17700_, _17690_);
  nand _50256_ (_17702_, _17701_, _06760_);
  nand _50257_ (_17703_, _17702_, _17680_);
  nand _50258_ (_17704_, _17703_, _06731_);
  nand _50259_ (_17705_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  nand _50260_ (_17706_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  nand _50261_ (_17707_, _17706_, _17705_);
  nand _50262_ (_17708_, _17707_, _06717_);
  nand _50263_ (_17709_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  nand _50264_ (_17710_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  nand _50265_ (_17711_, _17710_, _17709_);
  nand _50266_ (_17712_, _17711_, _06716_);
  nand _50267_ (_17713_, _17712_, _17708_);
  nand _50268_ (_17714_, _17713_, _06748_);
  nand _50269_ (_17715_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  nand _50270_ (_17716_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  nand _50271_ (_17717_, _17716_, _17715_);
  nand _50272_ (_17718_, _17717_, _06717_);
  nand _50273_ (_17719_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  nand _50274_ (_17720_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  nand _50275_ (_17721_, _17720_, _17719_);
  nand _50276_ (_17722_, _17721_, _06716_);
  nand _50277_ (_17723_, _17722_, _17718_);
  nand _50278_ (_17724_, _17723_, _06751_);
  nand _50279_ (_17725_, _17724_, _17714_);
  nand _50280_ (_17726_, _17725_, _06761_);
  nor _50281_ (_17727_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  nor _50282_ (_17728_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  nor _50283_ (_17729_, _17728_, _17727_);
  nand _50284_ (_17730_, _17729_, _06716_);
  nand _50285_ (_17731_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  nand _50286_ (_17732_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  nand _50287_ (_17733_, _17732_, _17731_);
  nand _50288_ (_17734_, _17733_, _06717_);
  nand _50289_ (_17735_, _17734_, _17730_);
  nand _50290_ (_17736_, _17735_, _06748_);
  nor _50291_ (_17737_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  nor _50292_ (_17738_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  nor _50293_ (_17739_, _17738_, _17737_);
  nand _50294_ (_17740_, _17739_, _06716_);
  nand _50295_ (_17741_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  nand _50296_ (_17742_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  nand _50297_ (_17743_, _17742_, _17741_);
  nand _50298_ (_17744_, _17743_, _06717_);
  nand _50299_ (_17745_, _17744_, _17740_);
  nand _50300_ (_17746_, _17745_, _06751_);
  nand _50301_ (_17747_, _17746_, _17736_);
  nand _50302_ (_17748_, _17747_, _06760_);
  nand _50303_ (_17749_, _17748_, _17726_);
  nand _50304_ (_17750_, _17749_, _06780_);
  nand _50305_ (_17751_, _17750_, _17704_);
  nand _50306_ (_17752_, _17751_, _06734_);
  nand _50307_ (_17753_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  nand _50308_ (_17754_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  nand _50309_ (_17755_, _17754_, _17753_);
  nand _50310_ (_17756_, _17755_, _06717_);
  nand _50311_ (_17757_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  nand _50312_ (_17758_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  nand _50313_ (_17759_, _17758_, _17757_);
  nand _50314_ (_17760_, _17759_, _06716_);
  nand _50315_ (_17761_, _17760_, _17756_);
  nand _50316_ (_17762_, _17761_, _06748_);
  nand _50317_ (_17763_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  nand _50318_ (_17764_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nand _50319_ (_17765_, _17764_, _17763_);
  nand _50320_ (_17766_, _17765_, _06717_);
  nand _50321_ (_17767_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nand _50322_ (_17768_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  nand _50323_ (_17769_, _17768_, _17767_);
  nand _50324_ (_17770_, _17769_, _06716_);
  nand _50325_ (_17771_, _17770_, _17766_);
  nand _50326_ (_17772_, _17771_, _06751_);
  nand _50327_ (_17773_, _17772_, _17762_);
  nand _50328_ (_17774_, _17773_, _06761_);
  nor _50329_ (_17775_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  nor _50330_ (_17776_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  nor _50331_ (_17777_, _17776_, _17775_);
  nand _50332_ (_17778_, _17777_, _06716_);
  nand _50333_ (_17779_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  nand _50334_ (_17780_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  nand _50335_ (_17781_, _17780_, _17779_);
  nand _50336_ (_17782_, _17781_, _06717_);
  nand _50337_ (_17783_, _17782_, _17778_);
  nand _50338_ (_17784_, _17783_, _06748_);
  nor _50339_ (_17785_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  nor _50340_ (_17787_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  nor _50341_ (_17788_, _17787_, _17785_);
  nand _50342_ (_17789_, _17788_, _06716_);
  nand _50343_ (_17790_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nand _50344_ (_17791_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  nand _50345_ (_17792_, _17791_, _17790_);
  nand _50346_ (_17793_, _17792_, _06717_);
  nand _50347_ (_17794_, _17793_, _17789_);
  nand _50348_ (_17795_, _17794_, _06751_);
  nand _50349_ (_17796_, _17795_, _17784_);
  nand _50350_ (_17797_, _17796_, _06760_);
  nand _50351_ (_17798_, _17797_, _17774_);
  nand _50352_ (_17799_, _17798_, _06780_);
  nand _50353_ (_17800_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  nand _50354_ (_17801_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  nand _50355_ (_17802_, _17801_, _17800_);
  nand _50356_ (_17803_, _17802_, _06717_);
  nand _50357_ (_17804_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  nand _50358_ (_17805_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  nand _50359_ (_17806_, _17805_, _17804_);
  nand _50360_ (_17807_, _17806_, _06716_);
  nand _50361_ (_17808_, _17807_, _17803_);
  nand _50362_ (_17809_, _17808_, _06748_);
  nand _50363_ (_17810_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  nand _50364_ (_17811_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  nand _50365_ (_17812_, _17811_, _17810_);
  nand _50366_ (_17813_, _17812_, _06717_);
  nand _50367_ (_17814_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  nand _50368_ (_17815_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  nand _50369_ (_17816_, _17815_, _17814_);
  nand _50370_ (_17817_, _17816_, _06716_);
  nand _50371_ (_17818_, _17817_, _17813_);
  nand _50372_ (_17819_, _17818_, _06751_);
  nand _50373_ (_17820_, _17819_, _17809_);
  nand _50374_ (_17821_, _17820_, _06761_);
  nor _50375_ (_17822_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  nor _50376_ (_17823_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  nor _50377_ (_17824_, _17823_, _17822_);
  nand _50378_ (_17825_, _17824_, _06717_);
  nor _50379_ (_17826_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  nor _50380_ (_17827_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  nor _50381_ (_17828_, _17827_, _17826_);
  nand _50382_ (_17829_, _17828_, _06716_);
  nand _50383_ (_17830_, _17829_, _17825_);
  nand _50384_ (_17831_, _17830_, _06748_);
  nor _50385_ (_17832_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  nor _50386_ (_17833_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  nor _50387_ (_17834_, _17833_, _17832_);
  nand _50388_ (_17835_, _17834_, _06717_);
  nor _50389_ (_17836_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  nor _50390_ (_17837_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  nor _50391_ (_17838_, _17837_, _17836_);
  nand _50392_ (_17839_, _17838_, _06716_);
  nand _50393_ (_17840_, _17839_, _17835_);
  nand _50394_ (_17841_, _17840_, _06751_);
  nand _50395_ (_17842_, _17841_, _17831_);
  nand _50396_ (_17843_, _17842_, _06760_);
  nand _50397_ (_17844_, _17843_, _17821_);
  nand _50398_ (_17845_, _17844_, _06731_);
  nand _50399_ (_17846_, _17845_, _17799_);
  nand _50400_ (_17847_, _17846_, _06733_);
  nand _50401_ (_17848_, _17847_, _17752_);
  nor _50402_ (_17849_, _17848_, _06723_);
  nand _50403_ (_17850_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  nand _50404_ (_17851_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  nand _50405_ (_17852_, _17851_, _17850_);
  nand _50406_ (_17853_, _17852_, _06717_);
  nand _50407_ (_17854_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  nand _50408_ (_17855_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  nand _50409_ (_17856_, _17855_, _17854_);
  nand _50410_ (_17857_, _17856_, _06716_);
  nand _50411_ (_17858_, _17857_, _17853_);
  nand _50412_ (_17859_, _17858_, _06748_);
  nand _50413_ (_17860_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  nand _50414_ (_17861_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  nand _50415_ (_17862_, _17861_, _17860_);
  nand _50416_ (_17863_, _17862_, _06717_);
  nand _50417_ (_17864_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  nand _50418_ (_17865_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  nand _50419_ (_17866_, _17865_, _17864_);
  nand _50420_ (_17868_, _17866_, _06716_);
  nand _50421_ (_17869_, _17868_, _17863_);
  nand _50422_ (_17870_, _17869_, _06751_);
  nand _50423_ (_17871_, _17870_, _17859_);
  nand _50424_ (_17872_, _17871_, _06761_);
  nor _50425_ (_17873_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  nor _50426_ (_17874_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  nor _50427_ (_17875_, _17874_, _17873_);
  nand _50428_ (_17876_, _17875_, _06716_);
  nand _50429_ (_17877_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  nand _50430_ (_17878_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nand _50431_ (_17879_, _17878_, _17877_);
  nand _50432_ (_17880_, _17879_, _06717_);
  nand _50433_ (_17881_, _17880_, _17876_);
  nand _50434_ (_17882_, _17881_, _06748_);
  nor _50435_ (_17883_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  nor _50436_ (_17884_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  nor _50437_ (_17885_, _17884_, _17883_);
  nand _50438_ (_17886_, _17885_, _06716_);
  nand _50439_ (_17887_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  nand _50440_ (_17888_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  nand _50441_ (_17889_, _17888_, _17887_);
  nand _50442_ (_17890_, _17889_, _06717_);
  nand _50443_ (_17891_, _17890_, _17886_);
  nand _50444_ (_17892_, _17891_, _06751_);
  nand _50445_ (_17893_, _17892_, _17882_);
  nand _50446_ (_17894_, _17893_, _06760_);
  nand _50447_ (_17895_, _17894_, _17872_);
  nand _50448_ (_17896_, _17895_, _06780_);
  nand _50449_ (_17897_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  nand _50450_ (_17898_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  nand _50451_ (_17899_, _17898_, _17897_);
  nand _50452_ (_17900_, _17899_, _06717_);
  nand _50453_ (_17901_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  nand _50454_ (_17902_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  nand _50455_ (_17903_, _17902_, _17901_);
  nand _50456_ (_17904_, _17903_, _06716_);
  nand _50457_ (_17905_, _17904_, _17900_);
  nand _50458_ (_17906_, _17905_, _06748_);
  nand _50459_ (_17907_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  nand _50460_ (_17908_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  nand _50461_ (_17909_, _17908_, _17907_);
  nand _50462_ (_17910_, _17909_, _06717_);
  nand _50463_ (_17911_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  nand _50464_ (_17912_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  nand _50465_ (_17913_, _17912_, _17911_);
  nand _50466_ (_17914_, _17913_, _06716_);
  nand _50467_ (_17915_, _17914_, _17910_);
  nand _50468_ (_17916_, _17915_, _06751_);
  nand _50469_ (_17917_, _17916_, _17906_);
  nand _50470_ (_17918_, _17917_, _06761_);
  nor _50471_ (_17919_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  nor _50472_ (_17920_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  nor _50473_ (_17921_, _17920_, _17919_);
  nand _50474_ (_17922_, _17921_, _06717_);
  nor _50475_ (_17923_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  nor _50476_ (_17924_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  nor _50477_ (_17925_, _17924_, _17923_);
  nand _50478_ (_17926_, _17925_, _06716_);
  nand _50479_ (_17927_, _17926_, _17922_);
  nand _50480_ (_17929_, _17927_, _06748_);
  nor _50481_ (_17930_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  nor _50482_ (_17931_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  nor _50483_ (_17932_, _17931_, _17930_);
  nand _50484_ (_17933_, _17932_, _06717_);
  nor _50485_ (_17934_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  nor _50486_ (_17935_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  nor _50487_ (_17936_, _17935_, _17934_);
  nand _50488_ (_17937_, _17936_, _06716_);
  nand _50489_ (_17938_, _17937_, _17933_);
  nand _50490_ (_17939_, _17938_, _06751_);
  nand _50491_ (_17940_, _17939_, _17929_);
  nand _50492_ (_17941_, _17940_, _06760_);
  nand _50493_ (_17942_, _17941_, _17918_);
  nand _50494_ (_17943_, _17942_, _06731_);
  nand _50495_ (_17944_, _17943_, _17896_);
  nand _50496_ (_17945_, _17944_, _06734_);
  nor _50497_ (_17946_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  nor _50498_ (_17947_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  nor _50499_ (_17948_, _17947_, _17946_);
  nand _50500_ (_17949_, _17948_, _06717_);
  nor _50501_ (_17950_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  nor _50502_ (_17951_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nor _50503_ (_17952_, _17951_, _17950_);
  nand _50504_ (_17953_, _17952_, _06716_);
  nand _50505_ (_17954_, _17953_, _17949_);
  nand _50506_ (_17955_, _17954_, _06751_);
  nor _50507_ (_17956_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  nor _50508_ (_17957_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  nor _50509_ (_17958_, _17957_, _17956_);
  nand _50510_ (_17959_, _17958_, _06717_);
  nor _50511_ (_17960_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  nor _50512_ (_17961_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  nor _50513_ (_17962_, _17961_, _17960_);
  nand _50514_ (_17963_, _17962_, _06716_);
  nand _50515_ (_17964_, _17963_, _17959_);
  nand _50516_ (_17965_, _17964_, _06748_);
  nand _50517_ (_17966_, _17965_, _17955_);
  nand _50518_ (_17967_, _17966_, _06760_);
  nand _50519_ (_17968_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  nand _50520_ (_17969_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  nand _50521_ (_17970_, _17969_, _17968_);
  nand _50522_ (_17971_, _17970_, _06717_);
  nand _50523_ (_17972_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  nand _50524_ (_17973_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  nand _50525_ (_17974_, _17973_, _17972_);
  nand _50526_ (_17975_, _17974_, _06716_);
  nand _50527_ (_17976_, _17975_, _17971_);
  nand _50528_ (_17977_, _17976_, _06751_);
  nand _50529_ (_17978_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  nand _50530_ (_17979_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  nand _50531_ (_17980_, _17979_, _17978_);
  nand _50532_ (_17981_, _17980_, _06717_);
  nand _50533_ (_17982_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  nand _50534_ (_17983_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  nand _50535_ (_17984_, _17983_, _17982_);
  nand _50536_ (_17985_, _17984_, _06716_);
  nand _50537_ (_17986_, _17985_, _17981_);
  nand _50538_ (_17987_, _17986_, _06748_);
  nand _50539_ (_17988_, _17987_, _17977_);
  nand _50540_ (_17989_, _17988_, _06761_);
  nand _50541_ (_17990_, _17989_, _17967_);
  nand _50542_ (_17991_, _17990_, _06731_);
  nor _50543_ (_17992_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  nor _50544_ (_17993_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nor _50545_ (_17994_, _17993_, _17992_);
  nand _50546_ (_17995_, _17994_, _06716_);
  nand _50547_ (_17996_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  nand _50548_ (_17997_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nand _50549_ (_17998_, _17997_, _17996_);
  nand _50550_ (_17999_, _17998_, _06717_);
  nand _50551_ (_18000_, _17999_, _17995_);
  nand _50552_ (_18001_, _18000_, _06751_);
  nor _50553_ (_18002_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  nor _50554_ (_18003_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nor _50555_ (_18004_, _18003_, _18002_);
  nand _50556_ (_18005_, _18004_, _06716_);
  nand _50557_ (_18006_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  nand _50558_ (_18007_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  nand _50559_ (_18008_, _18007_, _18006_);
  nand _50560_ (_18009_, _18008_, _06717_);
  nand _50561_ (_18010_, _18009_, _18005_);
  nand _50562_ (_18011_, _18010_, _06748_);
  nand _50563_ (_18012_, _18011_, _18001_);
  nand _50564_ (_18013_, _18012_, _06760_);
  nand _50565_ (_18014_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  nand _50566_ (_18015_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  nand _50567_ (_18016_, _18015_, _18014_);
  nand _50568_ (_18017_, _18016_, _06717_);
  nand _50569_ (_18018_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  nand _50570_ (_18019_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  nand _50571_ (_18020_, _18019_, _18018_);
  nand _50572_ (_18021_, _18020_, _06716_);
  nand _50573_ (_18022_, _18021_, _18017_);
  nand _50574_ (_18023_, _18022_, _06751_);
  nand _50575_ (_18024_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  nand _50576_ (_18025_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  nand _50577_ (_18026_, _18025_, _18024_);
  nand _50578_ (_18027_, _18026_, _06717_);
  nand _50579_ (_18028_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  nand _50580_ (_18029_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  nand _50581_ (_18030_, _18029_, _18028_);
  nand _50582_ (_18031_, _18030_, _06716_);
  nand _50583_ (_18032_, _18031_, _18027_);
  nand _50584_ (_18033_, _18032_, _06748_);
  nand _50585_ (_18034_, _18033_, _18023_);
  nand _50586_ (_18035_, _18034_, _06761_);
  nand _50587_ (_18036_, _18035_, _18013_);
  nand _50588_ (_18037_, _18036_, _06780_);
  nand _50589_ (_18038_, _18037_, _17991_);
  nand _50590_ (_18039_, _18038_, _06733_);
  nand _50591_ (_18040_, _18039_, _17945_);
  nor _50592_ (_18041_, _18040_, _13106_);
  nor _50593_ (_18042_, _18041_, _17849_);
  nor _50594_ (_18043_, _18042_, _25843_);
  nor _50595_ (_18044_, _18043_, _17658_);
  nor _50596_ (_18045_, _18044_, _13105_);
  not _50597_ (_18046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nand _50598_ (_18047_, _13105_, _18046_);
  nand _50599_ (_18048_, _18047_, _26487_);
  nor _50600_ (_07173_, _18048_, _18045_);
  nand _50601_ (_18049_, _12567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nand _50602_ (_18050_, _12566_, _25203_);
  nand _50603_ (_07176_, _18050_, _18049_);
  nand _50604_ (_18051_, _09547_, _25099_);
  nand _50605_ (_18052_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nand _50606_ (_07180_, _18052_, _18051_);
  nand _50607_ (_18053_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  nand _50608_ (_18054_, _08230_, _24789_);
  nand _50609_ (_07187_, _18054_, _18053_);
  nand _50610_ (_18056_, _12465_, _24789_);
  nand _50611_ (_18057_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  nand _50612_ (_07195_, _18057_, _18056_);
  nor _50613_ (_18058_, _00631_, _24795_);
  nand _50614_ (_18059_, _18058_, _24789_);
  not _50615_ (_18060_, _18058_);
  nand _50616_ (_18061_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  nand _50617_ (_07199_, _18061_, _18059_);
  nand _50618_ (_18062_, _12465_, _25039_);
  nand _50619_ (_18063_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nand _50620_ (_28278_, _18063_, _18062_);
  nor _50621_ (_18064_, _07818_, _24882_);
  nand _50622_ (_18065_, _18064_, _25039_);
  not _50623_ (_18066_, _18064_);
  nand _50624_ (_18067_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nand _50625_ (_07203_, _18067_, _18065_);
  nand _50626_ (_18068_, _12699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nand _50627_ (_18069_, _12698_, _28096_);
  nand _50628_ (_07207_, _18069_, _18068_);
  nand _50629_ (_18070_, _12619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  nand _50630_ (_18071_, _12618_, _25039_);
  nand _50631_ (_07222_, _18071_, _18070_);
  nand _50632_ (_18072_, _12591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  nand _50633_ (_18073_, _12590_, _24927_);
  nand _50634_ (_07224_, _18073_, _18072_);
  nand _50635_ (_18074_, _18064_, _25203_);
  nand _50636_ (_18075_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  nand _50637_ (_07231_, _18075_, _18074_);
  nand _50638_ (_18076_, _18064_, _28096_);
  nand _50639_ (_18077_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nand _50640_ (_07233_, _18077_, _18076_);
  nand _50641_ (_18078_, _12465_, _24830_);
  nand _50642_ (_18079_, _12467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  nand _50643_ (_07253_, _18079_, _18078_);
  nand _50644_ (_18080_, _12522_, _25099_);
  nand _50645_ (_18081_, _12524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  nand _50646_ (_07256_, _18081_, _18080_);
  nand _50647_ (_18082_, _12498_, _28096_);
  nand _50648_ (_18083_, _12500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  nand _50649_ (_07261_, _18083_, _18082_);
  nand _50650_ (_18084_, _12483_, _25203_);
  nand _50651_ (_18085_, _12485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  nand _50652_ (_28277_, _18085_, _18084_);
  nand _50653_ (_18086_, _18058_, _25150_);
  nand _50654_ (_18087_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  nand _50655_ (_07267_, _18087_, _18086_);
  nand _50656_ (_18088_, _12672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  nand _50657_ (_18089_, _12671_, _25203_);
  nand _50658_ (_07270_, _18089_, _18088_);
  nand _50659_ (_18090_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nand _50660_ (_18091_, _08212_, _25099_);
  nand _50661_ (_07272_, _18091_, _18090_);
  nand _50662_ (_18092_, _12413_, _25099_);
  nand _50663_ (_18093_, _12415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nand _50664_ (_07276_, _18093_, _18092_);
  nand _50665_ (_18094_, _08213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  nand _50666_ (_18095_, _08212_, _28096_);
  nand _50667_ (_07278_, _18095_, _18094_);
  nand _50668_ (_18096_, _18064_, _24927_);
  nand _50669_ (_18097_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nand _50670_ (_07280_, _18097_, _18096_);
  nand _50671_ (_18098_, _18064_, _24789_);
  nand _50672_ (_18099_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  nand _50673_ (_07285_, _18099_, _18098_);
  nand _50674_ (_18100_, _18064_, _25150_);
  nand _50675_ (_18101_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  nand _50676_ (_07289_, _18101_, _18100_);
  nand _50677_ (_18102_, _12763_, _24927_);
  nand _50678_ (_18103_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  nand _50679_ (_07295_, _18103_, _18102_);
  nand _50680_ (_18104_, _12857_, _25099_);
  nand _50681_ (_18105_, _12859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  nand _50682_ (_07297_, _18105_, _18104_);
  nand _50683_ (_18106_, _12976_, _25203_);
  nand _50684_ (_18107_, _12978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nand _50685_ (_28276_, _18107_, _18106_);
  nand _50686_ (_18108_, _17220_, _25150_);
  nand _50687_ (_18109_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  nand _50688_ (_07300_, _18109_, _18108_);
  nand _50689_ (_18110_, _17220_, _24830_);
  nand _50690_ (_18112_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nand _50691_ (_28274_, _18112_, _18110_);
  nor _50692_ (_18113_, _07818_, _00114_);
  nand _50693_ (_18114_, _18113_, _25039_);
  not _50694_ (_18115_, _18113_);
  nand _50695_ (_18116_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nand _50696_ (_07307_, _18116_, _18114_);
  nor _50697_ (_18117_, _00926_, _24889_);
  nand _50698_ (_18118_, _18117_, _25099_);
  not _50699_ (_18119_, _18117_);
  nand _50700_ (_18120_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nand _50701_ (_07311_, _18120_, _18118_);
  nor _50702_ (_18121_, _24889_, _24795_);
  nand _50703_ (_18122_, _18121_, _25039_);
  not _50704_ (_18123_, _18121_);
  nand _50705_ (_18124_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  nand _50706_ (_07314_, _18124_, _18122_);
  nor _50707_ (_18125_, _24889_, _24059_);
  nand _50708_ (_18126_, _18125_, _25150_);
  not _50709_ (_18127_, _18125_);
  nand _50710_ (_18128_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nand _50711_ (_07317_, _18128_, _18126_);
  nand _50712_ (_18129_, _18125_, _25099_);
  nand _50713_ (_18130_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nand _50714_ (_07319_, _18130_, _18129_);
  nor _50715_ (_18131_, _24978_, _24889_);
  nand _50716_ (_18132_, _18131_, _25099_);
  not _50717_ (_18133_, _18131_);
  nand _50718_ (_18134_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nand _50719_ (_07322_, _18134_, _18132_);
  nor _50720_ (_18135_, _00122_, _24889_);
  nand _50721_ (_18136_, _18135_, _24830_);
  not _50722_ (_18137_, _18135_);
  nand _50723_ (_18138_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  nand _50724_ (_07329_, _18138_, _18136_);
  nand _50725_ (_18139_, _09547_, _24830_);
  nand _50726_ (_18140_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  nand _50727_ (_07333_, _18140_, _18139_);
  nand _50728_ (_18141_, _04006_, _24789_);
  nand _50729_ (_18142_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  nand _50730_ (_07335_, _18142_, _18141_);
  nor _50731_ (_18143_, _07818_, _00629_);
  nand _50732_ (_18144_, _18143_, _25203_);
  not _50733_ (_18145_, _18143_);
  nand _50734_ (_18146_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  nand _50735_ (_07338_, _18146_, _18144_);
  nand _50736_ (_18147_, _24890_, _24830_);
  nand _50737_ (_18148_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nand _50738_ (_07343_, _18148_, _18147_);
  nand _50739_ (_18149_, _05739_, _24789_);
  nand _50740_ (_18150_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  nand _50741_ (_28249_, _18150_, _18149_);
  nand _50742_ (_18151_, _18143_, _24927_);
  nand _50743_ (_18152_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  nand _50744_ (_07347_, _18152_, _18151_);
  nand _50745_ (_18153_, _09944_, _24927_);
  nand _50746_ (_18154_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  nand _50747_ (_07353_, _18154_, _18153_);
  nand _50748_ (_18155_, _18143_, _25039_);
  nand _50749_ (_18156_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  nand _50750_ (_07356_, _18156_, _18155_);
  nor _50751_ (_18157_, _28057_, _25057_);
  nand _50752_ (_18158_, _18157_, _25039_);
  not _50753_ (_18159_, _18157_);
  nand _50754_ (_18160_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  nand _50755_ (_07358_, _18160_, _18158_);
  nand _50756_ (_18161_, _18157_, _24830_);
  nand _50757_ (_18162_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  nand _50758_ (_07360_, _18162_, _18161_);
  nand _50759_ (_18163_, _12010_, _25039_);
  nand _50760_ (_18164_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nand _50761_ (_07380_, _18164_, _18163_);
  nand _50762_ (_18165_, _01371_, _25150_);
  nand _50763_ (_18166_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nand _50764_ (_07382_, _18166_, _18165_);
  nand _50765_ (_18167_, _01371_, _28096_);
  nand _50766_ (_18168_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  nand _50767_ (_07384_, _18168_, _18167_);
  nand _50768_ (_18169_, _08354_, _24927_);
  nand _50769_ (_18170_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  nand _50770_ (_28241_, _18170_, _18169_);
  nand _50771_ (_18171_, _12710_, _28096_);
  nand _50772_ (_18172_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  nand _50773_ (_07390_, _18172_, _18171_);
  nor _50774_ (_18173_, _00114_, _24889_);
  nand _50775_ (_18174_, _18173_, _24927_);
  not _50776_ (_18175_, _18173_);
  nand _50777_ (_18176_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  nand _50778_ (_28252_, _18176_, _18174_);
  nand _50779_ (_18177_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nand _50780_ (_18178_, _08230_, _25203_);
  nand _50781_ (_28310_, _18178_, _18177_);
  nand _50782_ (_18179_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  nand _50783_ (_18180_, _08230_, _28096_);
  nand _50784_ (_07397_, _18180_, _18179_);
  nand _50785_ (_18181_, _10222_, _24830_);
  nand _50786_ (_18182_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  nand _50787_ (_07401_, _18182_, _18181_);
  nor _50788_ (_18183_, _13042_, _02509_);
  nand _50789_ (_18184_, _13042_, _05277_);
  nand _50790_ (_18185_, _18184_, _25630_);
  nor _50791_ (_18186_, _18185_, _18183_);
  nand _50792_ (_18187_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _50793_ (_18188_, _13040_, _24842_);
  nand _50794_ (_18189_, _18188_, _24717_);
  nor _50795_ (_18190_, _18188_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _50796_ (_18191_, _18190_, _26245_);
  nand _50797_ (_18192_, _18191_, _18189_);
  nand _50798_ (_18193_, _18192_, _18187_);
  nor _50799_ (_18194_, _18193_, _18186_);
  nor _50800_ (_07403_, _18194_, rst);
  nor _50801_ (_18195_, _13042_, _01974_);
  nor _50802_ (_18196_, _13041_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _50803_ (_18197_, _18196_);
  nand _50804_ (_18198_, _18197_, _25630_);
  nor _50805_ (_18199_, _18198_, _18195_);
  nand _50806_ (_18200_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _50807_ (_18201_, _13041_, _24717_);
  nor _50808_ (_18202_, _18196_, _26245_);
  nand _50809_ (_18203_, _18202_, _18201_);
  nand _50810_ (_18204_, _18203_, _18200_);
  nor _50811_ (_18205_, _18204_, _18199_);
  nor _50812_ (_07405_, _18205_, rst);
  nand _50813_ (_18206_, _01402_, _28096_);
  nand _50814_ (_18207_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  nand _50815_ (_07407_, _18207_, _18206_);
  nor _50816_ (_18208_, _13042_, _02685_);
  nand _50817_ (_18209_, _13042_, _05290_);
  nand _50818_ (_18210_, _18209_, _25630_);
  nor _50819_ (_18211_, _18210_, _18208_);
  nand _50820_ (_18212_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _50821_ (_18213_, _13039_, _03583_);
  nand _50822_ (_18214_, _18213_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _50823_ (_18215_, _24051_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _50824_ (_18216_, _18215_, _00381_);
  nand _50825_ (_18217_, _18216_, _13039_);
  nand _50826_ (_18218_, _18217_, _18214_);
  nand _50827_ (_18219_, _18218_, _26244_);
  nand _50828_ (_18220_, _18219_, _18212_);
  nor _50829_ (_18221_, _18220_, _18211_);
  nor _50830_ (_07410_, _18221_, rst);
  nor _50831_ (_18223_, _13042_, _02620_);
  not _50832_ (_18224_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _50833_ (_18225_, _13042_, _18224_);
  nand _50834_ (_18226_, _18225_, _25630_);
  nor _50835_ (_18227_, _18226_, _18223_);
  nand _50836_ (_18228_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _50837_ (_18229_, _13040_, _00263_);
  nand _50838_ (_18230_, _18229_, _24717_);
  nor _50839_ (_18231_, _18229_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _50840_ (_18232_, _18231_, _26245_);
  nand _50841_ (_18233_, _18232_, _18230_);
  nand _50842_ (_18234_, _18233_, _18228_);
  nor _50843_ (_18235_, _18234_, _18227_);
  nor _50844_ (_07411_, _18235_, rst);
  nor _50845_ (_18236_, _13042_, _02096_);
  nand _50846_ (_18237_, _13042_, _05285_);
  nand _50847_ (_18238_, _18237_, _25630_);
  nor _50848_ (_18239_, _18238_, _18236_);
  nand _50849_ (_18240_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor _50850_ (_18242_, _13040_, _00276_);
  nand _50851_ (_18243_, _18242_, _24717_);
  nor _50852_ (_18244_, _18242_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor _50853_ (_18245_, _18244_, _26245_);
  nand _50854_ (_18246_, _18245_, _18243_);
  nand _50855_ (_18247_, _18246_, _18240_);
  nor _50856_ (_18248_, _18247_, _18239_);
  nor _50857_ (_07413_, _18248_, rst);
  nor _50858_ (_18249_, _13042_, _02761_);
  nand _50859_ (_18250_, _13042_, _05275_);
  nand _50860_ (_18251_, _18250_, _25630_);
  nor _50861_ (_18252_, _18251_, _18249_);
  nand _50862_ (_18253_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor _50863_ (_18254_, _13040_, _00135_);
  nand _50864_ (_18255_, _18254_, _24717_);
  nor _50865_ (_18256_, _18254_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor _50866_ (_18257_, _18256_, _26245_);
  nand _50867_ (_18258_, _18257_, _18255_);
  nand _50868_ (_18259_, _18258_, _18253_);
  nor _50869_ (_18260_, _18259_, _18252_);
  nor _50870_ (_07416_, _18260_, rst);
  nand _50871_ (_18262_, _13056_, _24927_);
  nand _50872_ (_18263_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  nand _50873_ (_28275_, _18263_, _18262_);
  nor _50874_ (_18264_, _13042_, _02373_);
  nand _50875_ (_18265_, _13042_, _05282_);
  nand _50876_ (_18266_, _18265_, _25630_);
  nor _50877_ (_18267_, _18266_, _18264_);
  nand _50878_ (_18268_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor _50879_ (_18269_, _13040_, _01666_);
  nand _50880_ (_18270_, _18269_, _24717_);
  nor _50881_ (_18271_, _18269_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor _50882_ (_18272_, _18271_, _26245_);
  nand _50883_ (_18273_, _18272_, _18270_);
  nand _50884_ (_18274_, _18273_, _18268_);
  nor _50885_ (_18275_, _18274_, _18267_);
  nor _50886_ (_07419_, _18275_, rst);
  nand _50887_ (_18276_, _18064_, _25099_);
  nand _50888_ (_18277_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  nand _50889_ (_28273_, _18277_, _18276_);
  nand _50890_ (_18278_, _03911_, _25150_);
  nand _50891_ (_18279_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nand _50892_ (_07425_, _18279_, _18278_);
  nand _50893_ (_18280_, _18143_, _24789_);
  nand _50894_ (_18281_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  nand _50895_ (_07427_, _18281_, _18280_);
  nand _50896_ (_18282_, _12710_, _25203_);
  nand _50897_ (_18283_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  nand _50898_ (_07429_, _18283_, _18282_);
  nand _50899_ (_18284_, _12010_, _25203_);
  nand _50900_ (_18285_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nand _50901_ (_07430_, _18285_, _18284_);
  nor _50902_ (_18286_, _25057_, _24889_);
  nand _50903_ (_18287_, _18286_, _25203_);
  not _50904_ (_18288_, _18286_);
  nand _50905_ (_18289_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nand _50906_ (_07436_, _18289_, _18287_);
  nand _50907_ (_18290_, _18143_, _25150_);
  nand _50908_ (_18291_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nand _50909_ (_07438_, _18291_, _18290_);
  nand _50910_ (_18292_, _11542_, _25039_);
  nand _50911_ (_18293_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nand _50912_ (_07442_, _18293_, _18292_);
  nand _50913_ (_18294_, _04006_, _25099_);
  nand _50914_ (_18295_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nand _50915_ (_07446_, _18295_, _18294_);
  nand _50916_ (_18296_, _24890_, _24789_);
  nand _50917_ (_18297_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  nand _50918_ (_28253_, _18297_, _18296_);
  nand _50919_ (_18298_, _13080_, _25039_);
  nand _50920_ (_18299_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  nand _50921_ (_07455_, _18299_, _18298_);
  nand _50922_ (_18300_, _01182_, _24830_);
  nand _50923_ (_18301_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  nand _50924_ (_07458_, _18301_, _18300_);
  nand _50925_ (_18302_, _12710_, _25150_);
  nand _50926_ (_18303_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nand _50927_ (_28240_, _18303_, _18302_);
  nand _50928_ (_18304_, _08231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  nand _50929_ (_18305_, _08230_, _24927_);
  nand _50930_ (_07479_, _18305_, _18304_);
  nand _50931_ (_18306_, _00296_, _25628_);
  nor _50932_ (_18307_, _18306_, rst);
  nand _50933_ (_18308_, _18307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _50934_ (_18309_, _07948_, _25088_);
  not _50935_ (_18310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _50936_ (_18311_, _07960_, _18310_);
  not _50937_ (_18312_, _18311_);
  nor _50938_ (_18313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _50939_ (_18314_, _18313_);
  nor _50940_ (_18315_, _18314_, _07967_);
  not _50941_ (_18316_, _07946_);
  nor _50942_ (_18317_, _07979_, _07967_);
  not _50943_ (_18318_, _18317_);
  nor _50944_ (_18319_, _18318_, _18316_);
  nor _50945_ (_18320_, _18319_, _18315_);
  nor _50946_ (_18321_, _18320_, _18312_);
  not _50947_ (_18322_, _18321_);
  nand _50948_ (_18323_, _18322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not _50949_ (_18324_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _50950_ (_18325_, _18321_, _18324_);
  nand _50951_ (_18326_, _18325_, _18323_);
  nor _50952_ (_18327_, _18326_, _07948_);
  nor _50953_ (_18328_, _07941_, rst);
  not _50954_ (_18329_, _18328_);
  nor _50955_ (_18330_, _18329_, _18327_);
  nand _50956_ (_18331_, _18330_, _18309_);
  nand _50957_ (_07482_, _18331_, _18308_);
  nand _50958_ (_18332_, _18113_, _24789_);
  nand _50959_ (_18333_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  nand _50960_ (_07484_, _18333_, _18332_);
  nor _50961_ (_18334_, _00926_, _28057_);
  nand _50962_ (_18335_, _18334_, _24789_);
  not _50963_ (_18336_, _18334_);
  nand _50964_ (_18337_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  nand _50965_ (_07489_, _18337_, _18335_);
  nand _50966_ (_18338_, _18113_, _25150_);
  nand _50967_ (_18339_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  nand _50968_ (_07492_, _18339_, _18338_);
  nand _50969_ (_18340_, _17220_, _24789_);
  nand _50970_ (_18341_, _17222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  nand _50971_ (_07495_, _18341_, _18340_);
  nand _50972_ (_18342_, _18113_, _24927_);
  nand _50973_ (_18343_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  nand _50974_ (_07497_, _18343_, _18342_);
  nand _50975_ (_18344_, _18125_, _24789_);
  nand _50976_ (_18345_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  nand _50977_ (_28270_, _18345_, _18344_);
  nand _50978_ (_18346_, _09944_, _25099_);
  nand _50979_ (_18347_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nand _50980_ (_28243_, _18347_, _18346_);
  nand _50981_ (_18348_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nand _50982_ (_18349_, _08343_, _25099_);
  nand _50983_ (_07516_, _18349_, _18348_);
  nand _50984_ (_18350_, _18058_, _24927_);
  nand _50985_ (_18351_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  nand _50986_ (_07520_, _18351_, _18350_);
  nand _50987_ (_18352_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  nand _50988_ (_18353_, _08264_, _25150_);
  nand _50989_ (_07523_, _18353_, _18352_);
  nand _50990_ (_18354_, _18143_, _25099_);
  nand _50991_ (_18355_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nand _50992_ (_07524_, _18355_, _18354_);
  nand _50993_ (_18356_, _18143_, _24830_);
  nand _50994_ (_18357_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  nand _50995_ (_07527_, _18357_, _18356_);
  nand _50996_ (_18358_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nand _50997_ (_18359_, _08264_, _24927_);
  nand _50998_ (_07532_, _18359_, _18358_);
  nand _50999_ (_18360_, _18334_, _25203_);
  nand _51000_ (_18362_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nand _51001_ (_07543_, _18362_, _18360_);
  nand _51002_ (_18363_, _18334_, _25099_);
  nand _51003_ (_18364_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nand _51004_ (_07545_, _18364_, _18363_);
  nand _51005_ (_18365_, _18334_, _25150_);
  nand _51006_ (_18366_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nand _51007_ (_28250_, _18366_, _18365_);
  nand _51008_ (_18367_, _18173_, _25099_);
  nand _51009_ (_18368_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  nand _51010_ (_07569_, _18368_, _18367_);
  nand _51011_ (_18369_, _18173_, _28096_);
  nand _51012_ (_18370_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  nand _51013_ (_28251_, _18370_, _18369_);
  nand _51014_ (_18371_, _12710_, _25099_);
  nand _51015_ (_18372_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  nand _51016_ (_07579_, _18372_, _18371_);
  nor _51017_ (_07583_, _25886_, rst);
  nand _51018_ (_18373_, _12710_, _24927_);
  nand _51019_ (_18374_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  nand _51020_ (_07586_, _18374_, _18373_);
  nand _51021_ (_18375_, _12710_, _25039_);
  nand _51022_ (_18376_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nand _51023_ (_07588_, _18376_, _18375_);
  nor _51024_ (_07590_, _25717_, rst);
  nand _51025_ (_18377_, _08354_, _25099_);
  nand _51026_ (_18378_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  nand _51027_ (_07592_, _18378_, _18377_);
  nand _51028_ (_18379_, _08354_, _25203_);
  nand _51029_ (_18380_, _08356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nand _51030_ (_07594_, _18380_, _18379_);
  nor _51031_ (_18381_, _04950_, _25593_);
  nand _51032_ (_18382_, _18381_, _06599_);
  nand _51033_ (_18383_, _25802_, _25402_);
  nand _51034_ (_18384_, _18383_, _06559_);
  nand _51035_ (_18385_, _01048_, _25402_);
  nand _51036_ (_18386_, _18385_, _11889_);
  nor _51037_ (_18387_, _18386_, _18384_);
  nand _51038_ (_18388_, _18387_, _25409_);
  nor _51039_ (_18389_, _18388_, _18382_);
  not _51040_ (_18390_, _04042_);
  nor _51041_ (_18391_, _06494_, _04954_);
  not _51042_ (_18392_, _06678_);
  nor _51043_ (_18393_, _18392_, _25329_);
  nor _51044_ (_18394_, _18393_, _11896_);
  nand _51045_ (_18395_, _18394_, _18391_);
  nor _51046_ (_18396_, _18395_, _18390_);
  nand _51047_ (_18397_, _18396_, _18389_);
  not _51048_ (_18398_, _04276_);
  nand _51049_ (_18399_, _26201_, _25561_);
  nand _51050_ (_18401_, _18399_, _18398_);
  nand _51051_ (_18402_, _06630_, _04967_);
  nor _51052_ (_18403_, _18402_, _18401_);
  nand _51053_ (_18404_, _18403_, _06492_);
  nor _51054_ (_18405_, _18404_, _18397_);
  nor _51055_ (_18406_, _18405_, _24864_);
  nand _51056_ (_18407_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _51057_ (_18408_, _18407_, _11749_);
  nor _51058_ (_18409_, _18408_, _18406_);
  nor _51059_ (_28188_[0], _18409_, rst);
  nand _51060_ (_18410_, _18113_, _24830_);
  nand _51061_ (_18411_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nand _51062_ (_07599_, _18411_, _18410_);
  nand _51063_ (_18412_, _12010_, _25099_);
  nand _51064_ (_18413_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  nand _51065_ (_07604_, _18413_, _18412_);
  nor _51066_ (_18414_, _25627_, _25629_);
  nand _51067_ (_18415_, _18414_, _24717_);
  nor _51068_ (_18416_, _18414_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor _51069_ (_18417_, _18416_, _26245_);
  nand _51070_ (_18418_, _18417_, _18415_);
  nand _51071_ (_18419_, _03094_, _25088_);
  nor _51072_ (_18420_, _03094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor _51073_ (_18421_, _18420_, _25631_);
  nand _51074_ (_18422_, _18421_, _18419_);
  nand _51075_ (_18423_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nand _51076_ (_18424_, _18423_, _18422_);
  nor _51077_ (_18425_, _18424_, rst);
  nand _51078_ (_07608_, _18425_, _18418_);
  nand _51079_ (_18426_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  nand _51080_ (_18427_, _08264_, _24789_);
  nand _51081_ (_07611_, _18427_, _18426_);
  nand _51082_ (_18428_, _03894_, _24789_);
  nand _51083_ (_18429_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  nand _51084_ (_28371_, _18429_, _18428_);
  nand _51085_ (_18430_, _18157_, _25150_);
  nand _51086_ (_18431_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nand _51087_ (_07613_, _18431_, _18430_);
  nand _51088_ (_18432_, _01182_, _25039_);
  nand _51089_ (_18433_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  nand _51090_ (_07615_, _18433_, _18432_);
  nand _51091_ (_18434_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  nand _51092_ (_18435_, _03867_, _25039_);
  nand _51093_ (_07617_, _18435_, _18434_);
  nor _51094_ (_18436_, _01913_, _00276_);
  nand _51095_ (_18437_, _18436_, _24717_);
  nor _51096_ (_18438_, _18436_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor _51097_ (_18439_, _18438_, _26245_);
  nand _51098_ (_18440_, _18439_, _18437_);
  nand _51099_ (_18441_, _01919_, _25703_);
  nor _51100_ (_18442_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor _51101_ (_18443_, _18442_, _25631_);
  nand _51102_ (_18444_, _18443_, _18441_);
  nand _51103_ (_18445_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nand _51104_ (_18446_, _18445_, _18444_);
  nor _51105_ (_18447_, _18446_, rst);
  nand _51106_ (_07621_, _18447_, _18440_);
  nand _51107_ (_18448_, _09944_, _24830_);
  nand _51108_ (_18449_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  nand _51109_ (_07623_, _18449_, _18448_);
  nand _51110_ (_18450_, _18113_, _25203_);
  nand _51111_ (_18451_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nand _51112_ (_07628_, _18451_, _18450_);
  nor _51113_ (_18452_, _01714_, _00147_);
  nand _51114_ (_18453_, _18452_, _24717_);
  nor _51115_ (_18454_, _18452_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _51116_ (_18455_, _18454_, _26245_);
  nand _51117_ (_18456_, _18455_, _18453_);
  nand _51118_ (_18457_, _01720_, _25029_);
  nor _51119_ (_18458_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _51120_ (_18459_, _18458_, _25631_);
  nand _51121_ (_18460_, _18459_, _18457_);
  nand _51122_ (_18461_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand _51123_ (_18462_, _18461_, _18460_);
  nor _51124_ (_18463_, _18462_, rst);
  nand _51125_ (_07631_, _18463_, _18456_);
  nand _51126_ (_18464_, _09944_, _25203_);
  nand _51127_ (_18465_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  nand _51128_ (_07640_, _18465_, _18464_);
  nand _51129_ (_18466_, _13080_, _25203_);
  nand _51130_ (_18467_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nand _51131_ (_07642_, _18467_, _18466_);
  nand _51132_ (_18468_, _13080_, _24830_);
  nand _51133_ (_18469_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  nand _51134_ (_28244_, _18469_, _18468_);
  nand _51135_ (_18470_, _18113_, _28096_);
  nand _51136_ (_18471_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nand _51137_ (_07647_, _18471_, _18470_);
  nand _51138_ (_18472_, _05739_, _25099_);
  nand _51139_ (_18473_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  nand _51140_ (_28247_, _18473_, _18472_);
  nand _51141_ (_18474_, _13080_, _24789_);
  nand _51142_ (_18475_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  nand _51143_ (_28245_, _18475_, _18474_);
  nand _51144_ (_18476_, _05739_, _25039_);
  nand _51145_ (_18477_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nand _51146_ (_07667_, _18477_, _18476_);
  nand _51147_ (_18478_, _00276_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nand _51148_ (_18479_, _18478_, _03603_);
  nand _51149_ (_18480_, _18479_, _01541_);
  nand _51150_ (_18481_, _01542_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nand _51151_ (_18482_, _18481_, _18480_);
  nand _51152_ (_18483_, _18482_, _26244_);
  nand _51153_ (_18484_, _01551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nand _51154_ (_18485_, _01552_, _25680_);
  nand _51155_ (_18486_, _18485_, _18484_);
  nand _51156_ (_18487_, _18486_, _25630_);
  nand _51157_ (_18488_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nand _51158_ (_18489_, _18488_, _18487_);
  nor _51159_ (_18490_, _18489_, rst);
  nand _51160_ (_07671_, _18490_, _18483_);
  nand _51161_ (_18491_, _01402_, _24927_);
  nand _51162_ (_18492_, _01404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  nand _51163_ (_07673_, _18492_, _18491_);
  nand _51164_ (_18493_, _25203_, _24890_);
  nand _51165_ (_18494_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  nand _51166_ (_07676_, _18494_, _18493_);
  nand _51167_ (_18495_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  nand _51168_ (_18496_, _08501_, _24789_);
  nand _51169_ (_07678_, _18496_, _18495_);
  nand _51170_ (_18497_, _03442_, _25203_);
  nand _51171_ (_18498_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  nand _51172_ (_07680_, _18498_, _18497_);
  nand _51173_ (_18499_, _03442_, _25099_);
  nand _51174_ (_18500_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  nand _51175_ (_07681_, _18500_, _18499_);
  nand _51176_ (_18501_, _18117_, _25039_);
  nand _51177_ (_18502_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  nand _51178_ (_07684_, _18502_, _18501_);
  nand _51179_ (_18503_, _04006_, _24830_);
  nand _51180_ (_18504_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nand _51181_ (_28254_, _18504_, _18503_);
  nand _51182_ (_18505_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  nand _51183_ (_18506_, _08501_, _25150_);
  nand _51184_ (_28309_, _18506_, _18505_);
  nand _51185_ (_18507_, _18117_, _25203_);
  nand _51186_ (_18508_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  nand _51187_ (_07687_, _18508_, _18507_);
  nand _51188_ (_18509_, _03442_, _25150_);
  nand _51189_ (_18510_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  nand _51190_ (_07688_, _18510_, _18509_);
  nand _51191_ (_18511_, _07882_, _24830_);
  nand _51192_ (_18512_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  nand _51193_ (_07690_, _18512_, _18511_);
  nand _51194_ (_18513_, _11542_, _25203_);
  nand _51195_ (_18514_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  nand _51196_ (_07694_, _18514_, _18513_);
  nand _51197_ (_18515_, _11542_, _25099_);
  nand _51198_ (_18516_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nand _51199_ (_07695_, _18516_, _18515_);
  nand _51200_ (_18517_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  nand _51201_ (_18518_, _08501_, _24927_);
  nand _51202_ (_07697_, _18518_, _18517_);
  nor _51203_ (_18519_, _00393_, _25059_);
  nand _51204_ (_18520_, _18519_, _24830_);
  not _51205_ (_18521_, _18519_);
  nand _51206_ (_18522_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nand _51207_ (_07701_, _18522_, _18520_);
  nor _51208_ (_18523_, _25047_, _24889_);
  nand _51209_ (_18524_, _18523_, _24927_);
  not _51210_ (_18525_, _18523_);
  nand _51211_ (_18526_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  nand _51212_ (_07703_, _18526_, _18524_);
  nand _51213_ (_18527_, _18135_, _25150_);
  nand _51214_ (_18528_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  nand _51215_ (_28260_, _18528_, _18527_);
  nand _51216_ (_18529_, _18117_, _28096_);
  nand _51217_ (_18530_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  nand _51218_ (_07705_, _18530_, _18529_);
  nand _51219_ (_18531_, _18135_, _25039_);
  nand _51220_ (_18532_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  nand _51221_ (_07707_, _18532_, _18531_);
  nor _51222_ (_18533_, _28073_, _24889_);
  nand _51223_ (_18534_, _18533_, _25039_);
  not _51224_ (_18535_, _18533_);
  nand _51225_ (_18536_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nand _51226_ (_28262_, _18536_, _18534_);
  nor _51227_ (_18537_, _24889_, _28080_);
  nand _51228_ (_18538_, _18537_, _25039_);
  not _51229_ (_18539_, _18537_);
  nand _51230_ (_18540_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nand _51231_ (_07715_, _18540_, _18538_);
  nand _51232_ (_18541_, _18537_, _24830_);
  nand _51233_ (_18542_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  nand _51234_ (_07720_, _18542_, _18541_);
  nand _51235_ (_18543_, _18286_, _28096_);
  nand _51236_ (_18544_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  nand _51237_ (_07723_, _18544_, _18543_);
  nor _51238_ (_18545_, _24999_, _24889_);
  nand _51239_ (_18546_, _18545_, _28096_);
  not _51240_ (_18547_, _18545_);
  nand _51241_ (_18548_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nand _51242_ (_07729_, _18548_, _18546_);
  nand _51243_ (_18549_, _18286_, _24789_);
  nand _51244_ (_18550_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  nand _51245_ (_07731_, _18550_, _18549_);
  nand _51246_ (_18551_, _18307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  not _51247_ (_18552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _51248_ (_18553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not _51249_ (_18554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _51250_ (_18555_, _18554_, _18553_);
  not _51251_ (_18556_, _18555_);
  nor _51252_ (_18557_, _18556_, _18552_);
  not _51253_ (_18558_, _18557_);
  nor _51254_ (_18559_, _18324_, _18310_);
  not _51255_ (_18560_, _18559_);
  nor _51256_ (_18561_, _18560_, _07967_);
  nor _51257_ (_18562_, _07960_, _17063_);
  nand _51258_ (_18563_, _18562_, _18561_);
  nor _51259_ (_18564_, _18563_, _18558_);
  nor _51260_ (_18565_, _18564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _51261_ (_18566_, _18564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _51262_ (_18567_, _18566_, _18313_);
  not _51263_ (_18568_, _18567_);
  not _51264_ (_18569_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _51265_ (_18570_, _07967_, _07952_);
  nand _51266_ (_18571_, _18570_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _51267_ (_18572_, _18571_, _07944_);
  nand _51268_ (_18573_, _18572_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _51269_ (_18574_, _18573_, _18324_);
  nand _51270_ (_18575_, _18574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _51271_ (_18576_, _18575_, _07960_);
  nand _51272_ (_18577_, _18576_, _18557_);
  nor _51273_ (_18578_, _18577_, _18569_);
  nor _51274_ (_18579_, _18578_, _18316_);
  nor _51275_ (_18580_, _18579_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _51276_ (_18581_, _07979_, _18316_);
  nor _51277_ (_18582_, _18581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _51278_ (_18583_, _18582_, _18580_);
  nor _51279_ (_18584_, _18583_, _18568_);
  nor _51280_ (_18586_, _18584_, _18565_);
  nand _51281_ (_18587_, _18586_, _07983_);
  nand _51282_ (_18588_, _07948_, _25139_);
  nand _51283_ (_18589_, _18588_, _18587_);
  nand _51284_ (_18590_, _18589_, _18328_);
  nand _51285_ (_07735_, _18590_, _18551_);
  nand _51286_ (_18591_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  nand _51287_ (_18592_, _08264_, _25099_);
  nand _51288_ (_07737_, _18592_, _18591_);
  nand _51289_ (_18593_, _18545_, _25150_);
  nand _51290_ (_18594_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nand _51291_ (_07745_, _18594_, _18593_);
  nand _51292_ (_18595_, _09547_, _25039_);
  nand _51293_ (_18596_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  nand _51294_ (_28294_, _18596_, _18595_);
  nand _51295_ (_18597_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nand _51296_ (_18598_, _08264_, _25203_);
  nand _51297_ (_07759_, _18598_, _18597_);
  nand _51298_ (_18599_, _18117_, _24789_);
  nand _51299_ (_18600_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  nand _51300_ (_07770_, _18600_, _18599_);
  nand _51301_ (_18601_, _18121_, _28096_);
  nand _51302_ (_18602_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  nand _51303_ (_07772_, _18602_, _18601_);
  nand _51304_ (_18603_, _18117_, _25150_);
  nand _51305_ (_18604_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nand _51306_ (_07784_, _18604_, _18603_);
  nand _51307_ (_18605_, _08265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nand _51308_ (_18606_, _08264_, _28096_);
  nand _51309_ (_07786_, _18606_, _18605_);
  nand _51310_ (_18607_, _00991_, _24789_);
  nand _51311_ (_18608_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  nand _51312_ (_07788_, _18608_, _18607_);
  nand _51313_ (_18609_, _18121_, _24789_);
  nand _51314_ (_18610_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  nand _51315_ (_07792_, _18610_, _18609_);
  nand _51316_ (_18611_, _04006_, _25203_);
  nand _51317_ (_18612_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nand _51318_ (_28255_, _18612_, _18611_);
  nand _51319_ (_18613_, _18117_, _24927_);
  nand _51320_ (_18614_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  nand _51321_ (_28272_, _18614_, _18613_);
  nand _51322_ (_18615_, _18121_, _25150_);
  nand _51323_ (_18616_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  nand _51324_ (_07815_, _18616_, _18615_);
  nand _51325_ (_18617_, _18113_, _25099_);
  nand _51326_ (_18618_, _18115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  nand _51327_ (_07817_, _18618_, _18617_);
  nand _51328_ (_18619_, _18121_, _24927_);
  nand _51329_ (_18620_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nand _51330_ (_07820_, _18620_, _18619_);
  nand _51331_ (_18621_, _18143_, _28096_);
  nand _51332_ (_18622_, _18145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  nand _51333_ (_07822_, _18622_, _18621_);
  nand _51334_ (_18623_, _18064_, _24830_);
  nand _51335_ (_18624_, _18066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  nand _51336_ (_07837_, _18624_, _18623_);
  nand _51337_ (_18625_, _09547_, _25203_);
  nand _51338_ (_18626_, _09549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nand _51339_ (_07842_, _18626_, _18625_);
  nand _51340_ (_18627_, _01371_, _24789_);
  nand _51341_ (_18628_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  nand _51342_ (_07845_, _18628_, _18627_);
  nand _51343_ (_18629_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  nand _51344_ (_18630_, _08319_, _24789_);
  nand _51345_ (_07847_, _18630_, _18629_);
  nor _51346_ (_18631_, _18563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _51347_ (_18632_, _18631_);
  nor _51348_ (_18633_, _18632_, _07979_);
  nor _51349_ (_18634_, _18633_, _18313_);
  nand _51350_ (_18636_, _18563_, _18313_);
  nand _51351_ (_18637_, _18636_, _18555_);
  nor _51352_ (_18638_, _18637_, _18634_);
  nand _51353_ (_18639_, _18638_, _18552_);
  not _51354_ (_18640_, _18638_);
  nand _51355_ (_18641_, _18640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand _51356_ (_18642_, _18641_, _18639_);
  nand _51357_ (_18643_, _18642_, _07983_);
  nand _51358_ (_18644_, _07948_, _24920_);
  nand _51359_ (_18645_, _18644_, _18643_);
  nand _51360_ (_18646_, _18645_, _18328_);
  nand _51361_ (_18647_, _18307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand _51362_ (_08057_, _18647_, _18646_);
  nand _51363_ (_18648_, _17136_, _24927_);
  nand _51364_ (_18649_, _17138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  nand _51365_ (_08060_, _18649_, _18648_);
  nand _51366_ (_18650_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nand _51367_ (_18651_, _08319_, _25150_);
  nand _51368_ (_28308_, _18651_, _18650_);
  nand _51369_ (_18652_, _13056_, _25039_);
  nand _51370_ (_18654_, _13058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nand _51371_ (_08074_, _18654_, _18652_);
  nand _51372_ (_18655_, _18117_, _24830_);
  nand _51373_ (_18656_, _18119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  nand _51374_ (_28271_, _18656_, _18655_);
  nand _51375_ (_18657_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  nand _51376_ (_18658_, _08501_, _28096_);
  nand _51377_ (_08093_, _18658_, _18657_);
  nand _51378_ (_18659_, _08502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nand _51379_ (_18660_, _08501_, _25099_);
  nand _51380_ (_08098_, _18660_, _18659_);
  nand _51381_ (_18661_, _07979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand _51382_ (_18662_, _18661_, _05826_);
  not _51383_ (_18663_, _18662_);
  nand _51384_ (_18664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _51385_ (_18665_, _18664_, _18558_);
  nand _51386_ (_18666_, _18665_, _18663_);
  nor _51387_ (_18667_, _18666_, _18563_);
  not _51388_ (_18668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _51389_ (_18669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _18668_);
  nand _51390_ (_18670_, _18669_, _07960_);
  not _51391_ (_18671_, _07960_);
  nand _51392_ (_18672_, _18671_, _07664_);
  nor _51393_ (_18673_, _05826_, _18668_);
  nand _51394_ (_18674_, _18673_, _18672_);
  nand _51395_ (_18675_, _18674_, _18670_);
  nor _51396_ (_18676_, _18675_, _18667_);
  nand _51397_ (_18677_, _18676_, _17064_);
  nand _51398_ (_18678_, _18677_, _07983_);
  nor _51399_ (_08140_, _18678_, _18329_);
  nand _51400_ (_18679_, _12763_, _28096_);
  nand _51401_ (_18680_, _12765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  nand _51402_ (_08143_, _18680_, _18679_);
  nand _51403_ (_18681_, _12401_, _28096_);
  nand _51404_ (_18682_, _12403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nand _51405_ (_08145_, _18682_, _18681_);
  nand _51406_ (_18683_, _11919_, _25150_);
  nand _51407_ (_18684_, _11921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nand _51408_ (_08155_, _18684_, _18683_);
  nand _51409_ (_18685_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nand _51410_ (_18686_, _08343_, _24830_);
  nand _51411_ (_08162_, _18686_, _18685_);
  nand _51412_ (_18687_, _18307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _51413_ (_18688_, _07948_, _25029_);
  nand _51414_ (_18689_, _18661_, _18631_);
  nor _51415_ (_18690_, _18689_, _18553_);
  not _51416_ (_18691_, _18690_);
  nand _51417_ (_18692_, _18691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _51418_ (_18693_, _18690_, _18554_);
  nand _51419_ (_18694_, _18693_, _18692_);
  nor _51420_ (_18695_, _18694_, _07948_);
  nor _51421_ (_18696_, _18695_, _18329_);
  nand _51422_ (_18697_, _18696_, _18688_);
  nand _51423_ (_08169_, _18697_, _18687_);
  nand _51424_ (_18698_, _05739_, _25203_);
  nand _51425_ (_18699_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  nand _51426_ (_28248_, _18699_, _18698_);
  nand _51427_ (_18700_, _07908_, _25099_);
  nand _51428_ (_18701_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  nand _51429_ (_08268_, _18701_, _18700_);
  nand _51430_ (_18702_, _06826_, _28096_);
  nand _51431_ (_18703_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  nand _51432_ (_08288_, _18703_, _18702_);
  nand _51433_ (_18704_, _06826_, _25203_);
  nand _51434_ (_18705_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  nand _51435_ (_08292_, _18705_, _18704_);
  nand _51436_ (_18706_, _01066_, _01056_);
  nor _51437_ (_18707_, _18706_, _01041_);
  nor _51438_ (_18708_, _18707_, _24864_);
  nand _51439_ (_18709_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _51440_ (_18711_, _18709_, _01078_);
  nor _51441_ (_18712_, _18711_, _18708_);
  nor _51442_ (_28190_[0], _18712_, rst);
  nor _51443_ (_18713_, _00631_, _00393_);
  nand _51444_ (_18714_, _18713_, _25099_);
  not _51445_ (_18715_, _18713_);
  nand _51446_ (_18716_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nand _51447_ (_08303_, _18716_, _18714_);
  nand _51448_ (_18717_, _12910_, _28096_);
  nand _51449_ (_18718_, _12912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nand _51450_ (_08316_, _18718_, _18717_);
  nand _51451_ (_18719_, _11533_, _25203_);
  nand _51452_ (_18720_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nand _51453_ (_08318_, _18720_, _18719_);
  nand _51454_ (_18721_, _18713_, _28096_);
  nand _51455_ (_18722_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nand _51456_ (_08322_, _18722_, _18721_);
  nor _51457_ (_18723_, _05824_, _24782_);
  not _51458_ (_18724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nand _51459_ (_18725_, _05824_, _18724_);
  nand _51460_ (_18726_, _18725_, _26487_);
  nor _51461_ (_08328_, _18726_, _18723_);
  nand _51462_ (_18727_, _03911_, _24927_);
  nand _51463_ (_18728_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  nand _51464_ (_08330_, _18728_, _18727_);
  nand _51465_ (_18729_, _07882_, _28096_);
  nand _51466_ (_18730_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nand _51467_ (_08335_, _18730_, _18729_);
  nand _51468_ (_18731_, _18713_, _25203_);
  nand _51469_ (_18732_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  nand _51470_ (_08350_, _18732_, _18731_);
  nand _51471_ (_18733_, _06437_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor _51472_ (_18734_, _25469_, _25596_);
  nor _51473_ (_18735_, _26490_, _25802_);
  nor _51474_ (_18736_, _18735_, _18734_);
  not _51475_ (_18737_, _25585_);
  nor _51476_ (_18738_, _18737_, _25427_);
  nand _51477_ (_18739_, _18738_, _11902_);
  nor _51478_ (_18740_, _18739_, _18736_);
  nand _51479_ (_18741_, _25403_, _04949_);
  nor _51480_ (_18743_, _25510_, _25489_);
  nand _51481_ (_18744_, _18743_, _25514_);
  nor _51482_ (_18745_, _18744_, _18741_);
  nor _51483_ (_18746_, _18745_, _25803_);
  nor _51484_ (_18747_, _11892_, _11745_);
  nor _51485_ (_18748_, _06642_, _25509_);
  nor _51486_ (_18749_, _18748_, _18401_);
  nand _51487_ (_18750_, _18749_, _18747_);
  nor _51488_ (_18751_, _18750_, _18746_);
  nand _51489_ (_18752_, _18751_, _18740_);
  nand _51490_ (_18753_, _18752_, _00883_);
  nand _51491_ (_28189_[0], _18753_, _18733_);
  nand _51492_ (_18754_, _03876_, _25150_);
  nand _51493_ (_18755_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  nand _51494_ (_08364_, _18755_, _18754_);
  nand _51495_ (_18756_, _11533_, _24830_);
  nand _51496_ (_18757_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nand _51497_ (_08372_, _18757_, _18756_);
  nand _51498_ (_18758_, _12010_, _24789_);
  nand _51499_ (_18759_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  nand _51500_ (_08377_, _18759_, _18758_);
  nand _51501_ (_18760_, _11533_, _25150_);
  nand _51502_ (_18761_, _11535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nand _51503_ (_08388_, _18761_, _18760_);
  nand _51504_ (_18762_, _10222_, _25150_);
  nand _51505_ (_18763_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nand _51506_ (_08392_, _18763_, _18762_);
  nand _51507_ (_18764_, _03876_, _24789_);
  nand _51508_ (_18765_, _03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  nand _51509_ (_28280_, _18765_, _18764_);
  nand _51510_ (_18766_, _03139_, _24830_);
  nand _51511_ (_18767_, _03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nand _51512_ (_28246_, _18767_, _18766_);
  nand _51513_ (_18768_, _04111_, _25150_);
  nand _51514_ (_18769_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nand _51515_ (_08430_, _18769_, _18768_);
  nand _51516_ (_18770_, _08806_, _25203_);
  nand _51517_ (_18771_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  nand _51518_ (_08432_, _18771_, _18770_);
  nand _51519_ (_18772_, _18713_, _24830_);
  nand _51520_ (_18773_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nand _51521_ (_08446_, _18773_, _18772_);
  nand _51522_ (_18774_, _18713_, _24789_);
  nand _51523_ (_18775_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  nand _51524_ (_08484_, _18775_, _18774_);
  nand _51525_ (_18776_, _12104_, _24830_);
  nand _51526_ (_18777_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  nand _51527_ (_08488_, _18777_, _18776_);
  nand _51528_ (_18778_, _12104_, _25099_);
  nand _51529_ (_18779_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nand _51530_ (_08493_, _18779_, _18778_);
  nand _51531_ (_18780_, _12104_, _28096_);
  nand _51532_ (_18781_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  nand _51533_ (_08495_, _18781_, _18780_);
  nand _51534_ (_18782_, _12010_, _24927_);
  nand _51535_ (_18783_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  nand _51536_ (_08497_, _18783_, _18782_);
  nand _51537_ (_18784_, _12010_, _25150_);
  nand _51538_ (_18785_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  nand _51539_ (_08507_, _18785_, _18784_);
  nand _51540_ (_18786_, _18713_, _24927_);
  nand _51541_ (_18787_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  nand _51542_ (_08514_, _18787_, _18786_);
  nand _51543_ (_18788_, _11659_, _25099_);
  nand _51544_ (_18789_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  nand _51545_ (_08523_, _18789_, _18788_);
  nand _51546_ (_18790_, _07882_, _25203_);
  nand _51547_ (_18791_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nand _51548_ (_08530_, _18791_, _18790_);
  nand _51549_ (_18792_, _18713_, _25150_);
  nand _51550_ (_18793_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nand _51551_ (_08535_, _18793_, _18792_);
  nand _51552_ (_18794_, _06826_, _25150_);
  nand _51553_ (_18795_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nand _51554_ (_08539_, _18795_, _18794_);
  nor _51555_ (_18796_, _07637_, _04214_);
  nand _51556_ (_18797_, _07633_, _04215_);
  not _51557_ (_18798_, _07633_);
  nand _51558_ (_18799_, _18798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _51559_ (_18800_, _18799_, _18797_);
  nor _51560_ (_18801_, _18800_, _18796_);
  nor _51561_ (_18802_, _18801_, _01644_);
  nor _51562_ (_18803_, _01642_, _04215_);
  nor _51563_ (_18804_, _18803_, _18802_);
  nor _51564_ (_18805_, _18804_, _01573_);
  nor _51565_ (_18806_, _04175_, _25140_);
  nor _51566_ (_18807_, _18806_, _18805_);
  nor _51567_ (_08542_, _18807_, rst);
  nand _51568_ (_18808_, _04308_, _25150_);
  nand _51569_ (_18809_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  nand _51570_ (_08550_, _18809_, _18808_);
  nand _51571_ (_18810_, _06826_, _24789_);
  nand _51572_ (_18811_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  nand _51573_ (_08553_, _18811_, _18810_);
  nand _51574_ (_18812_, _06826_, _24927_);
  nand _51575_ (_18813_, _06828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  nand _51576_ (_08555_, _18813_, _18812_);
  nand _51577_ (_18814_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  nand _51578_ (_18815_, _28074_, _24927_);
  nand _51579_ (_08559_, _18815_, _18814_);
  nor _51580_ (_18816_, _00954_, _00631_);
  nand _51581_ (_18817_, _18816_, _24927_);
  not _51582_ (_18818_, _18816_);
  nand _51583_ (_18819_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  nand _51584_ (_28317_, _18819_, _18817_);
  nand _51585_ (_18820_, _00979_, _25150_);
  nand _51586_ (_18821_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  nand _51587_ (_28279_, _18821_, _18820_);
  nand _51588_ (_18822_, _18816_, _25150_);
  nand _51589_ (_18823_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  nand _51590_ (_08578_, _18823_, _18822_);
  nand _51591_ (_18824_, _08806_, _28096_);
  nand _51592_ (_18825_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nand _51593_ (_08582_, _18825_, _18824_);
  nand _51594_ (_18826_, _12100_, _24830_);
  nand _51595_ (_18827_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nand _51596_ (_08586_, _18827_, _18826_);
  nand _51597_ (_18828_, _18816_, _25099_);
  nand _51598_ (_18829_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  nand _51599_ (_08589_, _18829_, _18828_);
  nand _51600_ (_18830_, _18816_, _28096_);
  nand _51601_ (_18831_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  nand _51602_ (_08591_, _18831_, _18830_);
  nand _51603_ (_18832_, _12100_, _25099_);
  nand _51604_ (_18833_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  nand _51605_ (_08598_, _18833_, _18832_);
  nand _51606_ (_18834_, _04312_, _25150_);
  nand _51607_ (_18835_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  nand _51608_ (_08600_, _18835_, _18834_);
  nand _51609_ (_18836_, _18816_, _25203_);
  nand _51610_ (_18837_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nand _51611_ (_08601_, _18837_, _18836_);
  nand _51612_ (_18838_, _08806_, _25099_);
  nand _51613_ (_18839_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  nand _51614_ (_28295_, _18839_, _18838_);
  nor _51615_ (_18840_, _00631_, _00415_);
  nand _51616_ (_18841_, _18840_, _28096_);
  not _51617_ (_18842_, _18840_);
  nand _51618_ (_18843_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  nand _51619_ (_28320_, _18843_, _18841_);
  nand _51620_ (_18844_, _18840_, _25203_);
  nand _51621_ (_18845_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nand _51622_ (_08621_, _18845_, _18844_);
  nand _51623_ (_18846_, _18157_, _25203_);
  nand _51624_ (_18847_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  nand _51625_ (_08626_, _18847_, _18846_);
  nand _51626_ (_18848_, _18840_, _25039_);
  nand _51627_ (_18849_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  nand _51628_ (_08628_, _18849_, _18848_);
  nand _51629_ (_18850_, _12104_, _25150_);
  nand _51630_ (_18852_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nand _51631_ (_08632_, _18852_, _18850_);
  nand _51632_ (_18853_, _12104_, _24927_);
  nand _51633_ (_18854_, _12107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  nand _51634_ (_08634_, _18854_, _18853_);
  nand _51635_ (_18855_, _18816_, _24789_);
  nand _51636_ (_18856_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  nand _51637_ (_08646_, _18856_, _18855_);
  nand _51638_ (_18857_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  nand _51639_ (_18858_, _01388_, _28096_);
  nand _51640_ (_08648_, _18858_, _18857_);
  nand _51641_ (_18859_, _18840_, _24830_);
  nand _51642_ (_18860_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  nand _51643_ (_28318_, _18860_, _18859_);
  nand _51644_ (_18861_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nand _51645_ (_18862_, _04021_, _25203_);
  nand _51646_ (_08657_, _18862_, _18861_);
  nand _51647_ (_18863_, _18840_, _25099_);
  nand _51648_ (_18864_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nand _51649_ (_28319_, _18864_, _18863_);
  nand _51650_ (_18865_, _12100_, _25150_);
  nand _51651_ (_18866_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  nand _51652_ (_28283_, _18866_, _18865_);
  nand _51653_ (_18867_, _12100_, _24789_);
  nand _51654_ (_18868_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  nand _51655_ (_08662_, _18868_, _18867_);
  nand _51656_ (_18869_, _01389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nand _51657_ (_18870_, _01388_, _25203_);
  nand _51658_ (_08664_, _18870_, _18869_);
  nor _51659_ (_18871_, _00631_, _25047_);
  nand _51660_ (_18872_, _18871_, _25099_);
  not _51661_ (_18873_, _18871_);
  nand _51662_ (_18874_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  nand _51663_ (_08675_, _18874_, _18872_);
  nand _51664_ (_18875_, _12100_, _25039_);
  nand _51665_ (_18876_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  nand _51666_ (_08689_, _18876_, _18875_);
  nand _51667_ (_18877_, _18840_, _24927_);
  nand _51668_ (_18878_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  nand _51669_ (_08701_, _18878_, _18877_);
  nand _51670_ (_18880_, _18840_, _25150_);
  nand _51671_ (_18881_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  nand _51672_ (_08703_, _18881_, _18880_);
  nand _51673_ (_18882_, _12100_, _24927_);
  nand _51674_ (_18883_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  nand _51675_ (_08704_, _18883_, _18882_);
  nand _51676_ (_18884_, _18840_, _24789_);
  nand _51677_ (_18885_, _18842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  nand _51678_ (_08706_, _18885_, _18884_);
  nand _51679_ (_18886_, _12100_, _25203_);
  nand _51680_ (_18887_, _12102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nand _51681_ (_28282_, _18887_, _18886_);
  nand _51682_ (_18888_, _11659_, _25203_);
  nand _51683_ (_18889_, _11661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  nand _51684_ (_08718_, _18889_, _18888_);
  nand _51685_ (_18890_, _11827_, _25099_);
  nand _51686_ (_18891_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nand _51687_ (_28330_, _18891_, _18890_);
  nand _51688_ (_18892_, _11720_, _25203_);
  nand _51689_ (_18893_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  nand _51690_ (_08722_, _18893_, _18892_);
  nand _51691_ (_18894_, _11720_, _24927_);
  nand _51692_ (_18895_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nand _51693_ (_08724_, _18895_, _18894_);
  nand _51694_ (_18896_, _11827_, _24830_);
  nand _51695_ (_18897_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  nand _51696_ (_08726_, _18897_, _18896_);
  nand _51697_ (_18898_, _05739_, _28096_);
  nand _51698_ (_18899_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nand _51699_ (_08734_, _18899_, _18898_);
  nand _51700_ (_18900_, _07908_, _24830_);
  nand _51701_ (_18901_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  nand _51702_ (_08743_, _18901_, _18900_);
  nand _51703_ (_18902_, _18121_, _25099_);
  nand _51704_ (_18903_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  nand _51705_ (_08748_, _18903_, _18902_);
  nand _51706_ (_18904_, _18121_, _24830_);
  nand _51707_ (_18905_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  nand _51708_ (_08752_, _18905_, _18904_);
  nand _51709_ (_18906_, _11720_, _24789_);
  nand _51710_ (_18907_, _11724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  nand _51711_ (_08755_, _18907_, _18906_);
  nand _51712_ (_18908_, _11907_, _24830_);
  nand _51713_ (_18909_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  nand _51714_ (_28286_, _18909_, _18908_);
  nand _51715_ (_18910_, _12663_, _28096_);
  nand _51716_ (_18911_, _12665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand _51717_ (_08798_, _18911_, _18910_);
  nand _51718_ (_18912_, _18871_, _24927_);
  nand _51719_ (_18913_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  nand _51720_ (_28322_, _18913_, _18912_);
  nand _51721_ (_18914_, _10226_, _24927_);
  nand _51722_ (_18915_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand _51723_ (_08810_, _18915_, _18914_);
  nand _51724_ (_18916_, _18871_, _25150_);
  nand _51725_ (_18917_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nand _51726_ (_28323_, _18917_, _18916_);
  nand _51727_ (_18918_, _10226_, _25203_);
  nand _51728_ (_18919_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nand _51729_ (_08823_, _18919_, _18918_);
  nand _51730_ (_18920_, _18871_, _24789_);
  nand _51731_ (_18921_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  nand _51732_ (_08826_, _18921_, _18920_);
  nand _51733_ (_18922_, _04006_, _25039_);
  nand _51734_ (_18923_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  nand _51735_ (_08830_, _18923_, _18922_);
  nand _51736_ (_18924_, _12096_, _28096_);
  nand _51737_ (_18925_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nand _51738_ (_08832_, _18925_, _18924_);
  nand _51739_ (_18926_, _12096_, _25203_);
  nand _51740_ (_18927_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  nand _51741_ (_08846_, _18927_, _18926_);
  nand _51742_ (_18928_, _08806_, _24789_);
  nand _51743_ (_18929_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  nand _51744_ (_08850_, _18929_, _18928_);
  nand _51745_ (_18930_, _12096_, _25039_);
  nand _51746_ (_18931_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  nand _51747_ (_08855_, _18931_, _18930_);
  nand _51748_ (_18932_, _11907_, _28096_);
  nand _51749_ (_18933_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  nand _51750_ (_28287_, _18933_, _18932_);
  nand _51751_ (_18934_, _11907_, _25039_);
  nand _51752_ (_18935_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  nand _51753_ (_08867_, _18935_, _18934_);
  nand _51754_ (_18936_, _18058_, _24830_);
  nand _51755_ (_18937_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nand _51756_ (_08869_, _18937_, _18936_);
  nand _51757_ (_18938_, _11907_, _25150_);
  nand _51758_ (_18939_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nand _51759_ (_08871_, _18939_, _18938_);
  nand _51760_ (_18940_, _07819_, _25039_);
  nand _51761_ (_18941_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nand _51762_ (_08886_, _18941_, _18940_);
  nand _51763_ (_18942_, _07819_, _28096_);
  nand _51764_ (_18943_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  nand _51765_ (_08888_, _18943_, _18942_);
  nand _51766_ (_18944_, _07819_, _25099_);
  nand _51767_ (_18945_, _07823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  nand _51768_ (_08890_, _18945_, _18944_);
  nor _51769_ (_18946_, _00631_, _24059_);
  nand _51770_ (_18947_, _18946_, _24789_);
  not _51771_ (_18948_, _18946_);
  nand _51772_ (_18949_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  nand _51773_ (_08893_, _18949_, _18947_);
  nand _51774_ (_18950_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  nand _51775_ (_18951_, _08324_, _24789_);
  nand _51776_ (_08895_, _18951_, _18950_);
  nand _51777_ (_18952_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  nand _51778_ (_18953_, _08319_, _24830_);
  nand _51779_ (_08897_, _18953_, _18952_);
  nand _51780_ (_18954_, _18121_, _25203_);
  nand _51781_ (_18955_, _18123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  nand _51782_ (_08899_, _18955_, _18954_);
  nand _51783_ (_18956_, _18307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not _51784_ (_18957_, _18689_);
  nor _51785_ (_18958_, _18957_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _51786_ (_18959_, _18958_, _18690_);
  nand _51787_ (_18960_, _18959_, _07983_);
  nand _51788_ (_18961_, _07948_, _25194_);
  nand _51789_ (_18962_, _18961_, _18960_);
  nand _51790_ (_18963_, _18962_, _18328_);
  nand _51791_ (_08904_, _18963_, _18956_);
  nand _51792_ (_18964_, _03958_, _25039_);
  nand _51793_ (_18965_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  nand _51794_ (_28238_, _18965_, _18964_);
  nand _51795_ (_18966_, _03958_, _28096_);
  nand _51796_ (_18967_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nand _51797_ (_28237_, _18967_, _18966_);
  nand _51798_ (_18968_, _11907_, _24789_);
  nand _51799_ (_18969_, _11909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  nand _51800_ (_08923_, _18969_, _18968_);
  nand _51801_ (_18970_, _11874_, _28096_);
  nand _51802_ (_18971_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nand _51803_ (_08926_, _18971_, _18970_);
  nand _51804_ (_18972_, _04022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  nand _51805_ (_18973_, _04021_, _24830_);
  nand _51806_ (_08928_, _18973_, _18972_);
  nand _51807_ (_18974_, _09944_, _28096_);
  nand _51808_ (_18975_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nand _51809_ (_08930_, _18975_, _18974_);
  nand _51810_ (_18976_, _11874_, _25203_);
  nand _51811_ (_18977_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nand _51812_ (_08932_, _18977_, _18976_);
  nand _51813_ (_18978_, _11874_, _24927_);
  nand _51814_ (_18979_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  nand _51815_ (_08939_, _18979_, _18978_);
  nand _51816_ (_18980_, _00955_, _25203_);
  nand _51817_ (_18981_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nand _51818_ (_08941_, _18981_, _18980_);
  nand _51819_ (_18982_, _11874_, _24789_);
  nand _51820_ (_18984_, _11876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  nand _51821_ (_08944_, _18984_, _18982_);
  nand _51822_ (_18985_, _00394_, _24789_);
  nand _51823_ (_18986_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nand _51824_ (_08948_, _18986_, _18985_);
  nand _51825_ (_18987_, _18307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _51826_ (_18988_, _07948_, _25703_);
  nand _51827_ (_18989_, _18689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _51828_ (_18990_, _18561_, _18313_);
  nand _51829_ (_18991_, _18559_, _18319_);
  nand _51830_ (_18992_, _18991_, _18990_);
  nor _51831_ (_18993_, _07960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _51832_ (_18994_, _18993_, _18992_);
  nand _51833_ (_18995_, _18994_, _18989_);
  nor _51834_ (_18996_, _18995_, _07948_);
  nor _51835_ (_18997_, _18996_, _18329_);
  nand _51836_ (_18998_, _18997_, _18988_);
  nand _51837_ (_08950_, _18998_, _18987_);
  nand _51838_ (_18999_, _00394_, _28096_);
  nand _51839_ (_19000_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nand _51840_ (_08952_, _19000_, _18999_);
  nand _51841_ (_19001_, _28059_, _24789_);
  nand _51842_ (_19002_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  nand _51843_ (_28375_, _19002_, _19001_);
  nand _51844_ (_19003_, _28096_, _28059_);
  nand _51845_ (_19004_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  nand _51846_ (_08957_, _19004_, _19003_);
  nand _51847_ (_19005_, _01153_, _25203_);
  nand _51848_ (_19006_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  nand _51849_ (_08962_, _19006_, _19005_);
  nand _51850_ (_19007_, _01153_, _25099_);
  nand _51851_ (_19008_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nand _51852_ (_08963_, _19008_, _19007_);
  nand _51853_ (_19009_, _11633_, _24789_);
  nand _51854_ (_19010_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  nand _51855_ (_08965_, _19010_, _19009_);
  nand _51856_ (_19011_, _11633_, _25203_);
  nand _51857_ (_19012_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  nand _51858_ (_08969_, _19012_, _19011_);
  nand _51859_ (_19013_, _04251_, _24789_);
  nand _51860_ (_19014_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  nand _51861_ (_08971_, _19014_, _19013_);
  nand _51862_ (_19015_, _03894_, _25039_);
  nand _51863_ (_19016_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nand _51864_ (_08976_, _19016_, _19015_);
  nand _51865_ (_19017_, _03894_, _28096_);
  nand _51866_ (_19018_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  nand _51867_ (_08978_, _19018_, _19017_);
  nand _51868_ (_19019_, _18058_, _25203_);
  nand _51869_ (_19020_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nand _51870_ (_08980_, _19020_, _19019_);
  nand _51871_ (_19022_, _04006_, _24927_);
  nand _51872_ (_19023_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  nand _51873_ (_28256_, _19023_, _19022_);
  nor _51874_ (_19024_, _00631_, _00122_);
  nand _51875_ (_19025_, _19024_, _24927_);
  not _51876_ (_19026_, _19024_);
  nand _51877_ (_19027_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  nand _51878_ (_09009_, _19027_, _19025_);
  nand _51879_ (_19028_, _19024_, _24789_);
  nand _51880_ (_19029_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  nand _51881_ (_09011_, _19029_, _19028_);
  nand _51882_ (_19030_, _19024_, _25150_);
  nand _51883_ (_19031_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nand _51884_ (_09014_, _19031_, _19030_);
  nand _51885_ (_19032_, _12807_, _25150_);
  nand _51886_ (_19033_, _12809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nand _51887_ (_09016_, _19033_, _19032_);
  nand _51888_ (_19034_, _12096_, _25099_);
  nand _51889_ (_19035_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nand _51890_ (_09020_, _19035_, _19034_);
  nand _51891_ (_19036_, _18157_, _28096_);
  nand _51892_ (_19037_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  nand _51893_ (_09024_, _19037_, _19036_);
  nand _51894_ (_19038_, _28059_, _25203_);
  nand _51895_ (_19039_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nand _51896_ (_09026_, _19039_, _19038_);
  nand _51897_ (_19040_, _12096_, _24830_);
  nand _51898_ (_19041_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  nand _51899_ (_09039_, _19041_, _19040_);
  nand _51900_ (_19042_, _18157_, _25099_);
  nand _51901_ (_19043_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nand _51902_ (_28242_, _19043_, _19042_);
  nand _51903_ (_19044_, _18871_, _25039_);
  nand _51904_ (_19045_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  nand _51905_ (_09050_, _19045_, _19044_);
  nand _51906_ (_19046_, _18871_, _25203_);
  nand _51907_ (_19047_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  nand _51908_ (_28321_, _19047_, _19046_);
  nand _51909_ (_19048_, _03858_, _24927_);
  nand _51910_ (_19049_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  nand _51911_ (_09060_, _19049_, _19048_);
  nand _51912_ (_19050_, _03958_, _25150_);
  nand _51913_ (_19051_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  nand _51914_ (_09062_, _19051_, _19050_);
  nand _51915_ (_19052_, _03911_, _28096_);
  nand _51916_ (_19053_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  nand _51917_ (_09066_, _19053_, _19052_);
  nand _51918_ (_19054_, _11867_, _25099_);
  nand _51919_ (_19055_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nand _51920_ (_09068_, _19055_, _19054_);
  nand _51921_ (_19056_, _25039_, _24985_);
  nand _51922_ (_19057_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  nand _51923_ (_09072_, _19057_, _19056_);
  nand _51924_ (_19058_, _18125_, _25203_);
  nand _51925_ (_19059_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nand _51926_ (_09077_, _19059_, _19058_);
  nand _51927_ (_19060_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  nand _51928_ (_19061_, _08319_, _28096_);
  nand _51929_ (_09081_, _19061_, _19060_);
  nand _51930_ (_19062_, _18125_, _28096_);
  nand _51931_ (_19063_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nand _51932_ (_28269_, _19063_, _19062_);
  nand _51933_ (_19064_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  nand _51934_ (_19065_, _08319_, _25039_);
  nand _51935_ (_09089_, _19065_, _19064_);
  nand _51936_ (_19066_, _08320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nand _51937_ (_19067_, _08319_, _25203_);
  nand _51938_ (_28307_, _19067_, _19066_);
  nor _51939_ (_19068_, _24999_, _24984_);
  nand _51940_ (_19069_, _19068_, _25039_);
  not _51941_ (_19070_, _19068_);
  nand _51942_ (_19071_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nand _51943_ (_09095_, _19071_, _19069_);
  nand _51944_ (_19072_, _18058_, _28096_);
  nand _51945_ (_19073_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  nand _51946_ (_28329_, _19073_, _19072_);
  nand _51947_ (_19074_, _18125_, _24927_);
  nand _51948_ (_19075_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  nand _51949_ (_09106_, _19075_, _19074_);
  nand _51950_ (_19076_, _04251_, _25039_);
  nand _51951_ (_19077_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nand _51952_ (_09108_, _19077_, _19076_);
  nand _51953_ (_19078_, _18125_, _25039_);
  nand _51954_ (_19079_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nand _51955_ (_09110_, _19079_, _19078_);
  nand _51956_ (_19080_, _00979_, _28096_);
  nand _51957_ (_19081_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  nand _51958_ (_09112_, _19081_, _19080_);
  nand _51959_ (_19082_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  nand _51960_ (_19083_, _08324_, _24830_);
  nand _51961_ (_09114_, _19083_, _19082_);
  nand _51962_ (_19084_, _11867_, _28096_);
  nand _51963_ (_19085_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  nand _51964_ (_09141_, _19085_, _19084_);
  nand _51965_ (_19086_, _11867_, _25039_);
  nand _51966_ (_19087_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  nand _51967_ (_09155_, _19087_, _19086_);
  nand _51968_ (_19088_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  nand _51969_ (_19089_, _03867_, _24789_);
  nand _51970_ (_09159_, _19089_, _19088_);
  nand _51971_ (_19090_, _11867_, _25150_);
  nand _51972_ (_19091_, _11870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nand _51973_ (_28288_, _19091_, _19090_);
  nand _51974_ (_19092_, _11855_, _25099_);
  nand _51975_ (_19093_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nand _51976_ (_09183_, _19093_, _19092_);
  nor _51977_ (_19094_, _00415_, _25059_);
  nand _51978_ (_19095_, _19094_, _25203_);
  not _51979_ (_19096_, _19094_);
  nand _51980_ (_19098_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  nand _51981_ (_09239_, _19098_, _19095_);
  nand _51982_ (_19099_, _01153_, _25039_);
  nand _51983_ (_19100_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  nand _51984_ (_09252_, _19100_, _19099_);
  nand _51985_ (_19101_, _19094_, _28096_);
  nand _51986_ (_19102_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  nand _51987_ (_09261_, _19102_, _19101_);
  nand _51988_ (_19103_, _19094_, _25099_);
  nand _51989_ (_19104_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  nand _51990_ (_09263_, _19104_, _19103_);
  nand _51991_ (_19105_, _18946_, _25099_);
  nand _51992_ (_19106_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nand _51993_ (_09266_, _19106_, _19105_);
  nand _51994_ (_19107_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  nand _51995_ (_19108_, _08343_, _28096_);
  nand _51996_ (_09277_, _19108_, _19107_);
  nand _51997_ (_19109_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  nand _51998_ (_19110_, _08343_, _25039_);
  nand _51999_ (_09305_, _19110_, _19109_);
  nand _52000_ (_19111_, _05739_, _25150_);
  nand _52001_ (_19112_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  nand _52002_ (_09346_, _19112_, _19111_);
  nand _52003_ (_19113_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  nand _52004_ (_19114_, _08343_, _25203_);
  nand _52005_ (_28297_, _19114_, _19113_);
  nand _52006_ (_19115_, _19094_, _24927_);
  nand _52007_ (_19116_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  nand _52008_ (_09350_, _19116_, _19115_);
  nand _52009_ (_19117_, _19094_, _25150_);
  nand _52010_ (_19118_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nand _52011_ (_09360_, _19118_, _19117_);
  nor _52012_ (_19119_, _00954_, _25059_);
  nand _52013_ (_19120_, _19119_, _24927_);
  not _52014_ (_19121_, _19119_);
  nand _52015_ (_19122_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  nand _52016_ (_09413_, _19122_, _19120_);
  nand _52017_ (_19123_, _19119_, _25039_);
  nand _52018_ (_19124_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  nand _52019_ (_09419_, _19124_, _19123_);
  nand _52020_ (_19125_, _19119_, _25203_);
  nand _52021_ (_19126_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nand _52022_ (_09428_, _19126_, _19125_);
  nand _52023_ (_19127_, _18946_, _24830_);
  nand _52024_ (_19128_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  nand _52025_ (_09457_, _19128_, _19127_);
  nand _52026_ (_19129_, _11855_, _28096_);
  nand _52027_ (_19130_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nand _52028_ (_09471_, _19130_, _19129_);
  nand _52029_ (_19131_, _12688_, _24830_);
  nand _52030_ (_19132_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand _52031_ (_09474_, _19132_, _19131_);
  nand _52032_ (_19133_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nand _52033_ (_19134_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  nand _52034_ (_19135_, _19134_, _19133_);
  nand _52035_ (_19136_, _19135_, _06716_);
  nand _52036_ (_19137_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  nand _52037_ (_19138_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  nand _52038_ (_19139_, _19138_, _19137_);
  nand _52039_ (_19140_, _19139_, _06717_);
  nand _52040_ (_19141_, _19140_, _19136_);
  nand _52041_ (_19142_, _19141_, _06748_);
  nand _52042_ (_19143_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  nand _52043_ (_19144_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  nand _52044_ (_19145_, _19144_, _19143_);
  nand _52045_ (_19146_, _19145_, _06716_);
  nand _52046_ (_19147_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  nand _52047_ (_19148_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nand _52048_ (_19149_, _19148_, _19147_);
  nand _52049_ (_19150_, _19149_, _06717_);
  nand _52050_ (_19151_, _19150_, _19146_);
  nand _52051_ (_19152_, _19151_, _06751_);
  nand _52052_ (_19153_, _19152_, _19142_);
  nand _52053_ (_19154_, _19153_, _06761_);
  nand _52054_ (_19155_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nand _52055_ (_19156_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nand _52056_ (_19157_, _19156_, _19155_);
  nand _52057_ (_19158_, _19157_, _06717_);
  nor _52058_ (_19159_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  nor _52059_ (_19160_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  nor _52060_ (_19161_, _19160_, _19159_);
  nand _52061_ (_19162_, _19161_, _06716_);
  nand _52062_ (_19163_, _19162_, _19158_);
  nand _52063_ (_19164_, _19163_, _06748_);
  nand _52064_ (_19165_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nand _52065_ (_19166_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  nand _52066_ (_19167_, _19166_, _19165_);
  nand _52067_ (_19168_, _19167_, _06717_);
  nor _52068_ (_19169_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nor _52069_ (_19170_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nor _52070_ (_19171_, _19170_, _19169_);
  nand _52071_ (_19172_, _19171_, _06716_);
  nand _52072_ (_19173_, _19172_, _19168_);
  nand _52073_ (_19174_, _19173_, _06751_);
  nand _52074_ (_19175_, _19174_, _19164_);
  nand _52075_ (_19176_, _19175_, _06760_);
  nand _52076_ (_19177_, _19176_, _19154_);
  nand _52077_ (_19178_, _19177_, _06780_);
  nand _52078_ (_19179_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  nand _52079_ (_19180_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nand _52080_ (_19181_, _19180_, _19179_);
  nand _52081_ (_19182_, _19181_, _06717_);
  nand _52082_ (_19183_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nand _52083_ (_19184_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  nand _52084_ (_19185_, _19184_, _19183_);
  nand _52085_ (_19186_, _19185_, _06716_);
  nand _52086_ (_19187_, _19186_, _19182_);
  nand _52087_ (_19188_, _19187_, _06748_);
  nand _52088_ (_19189_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  nand _52089_ (_19190_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  nand _52090_ (_19191_, _19190_, _19189_);
  nand _52091_ (_19192_, _19191_, _06717_);
  nand _52092_ (_19193_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  nand _52093_ (_19194_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nand _52094_ (_19195_, _19194_, _19193_);
  nand _52095_ (_19196_, _19195_, _06716_);
  nand _52096_ (_19197_, _19196_, _19192_);
  nand _52097_ (_19198_, _19197_, _06751_);
  nand _52098_ (_19199_, _19198_, _19188_);
  nand _52099_ (_19200_, _19199_, _06761_);
  nor _52100_ (_19201_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  nor _52101_ (_19202_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  nor _52102_ (_19203_, _19202_, _19201_);
  nand _52103_ (_19204_, _19203_, _06717_);
  nor _52104_ (_19205_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  nor _52105_ (_19206_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nor _52106_ (_19207_, _19206_, _19205_);
  nand _52107_ (_19208_, _19207_, _06716_);
  nand _52108_ (_19209_, _19208_, _19204_);
  nand _52109_ (_19210_, _19209_, _06748_);
  nor _52110_ (_19211_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nor _52111_ (_19212_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  nor _52112_ (_19213_, _19212_, _19211_);
  nor _52113_ (_19214_, _19213_, _06716_);
  nor _52114_ (_19215_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  nor _52115_ (_19216_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  nor _52116_ (_19217_, _19216_, _19215_);
  nor _52117_ (_19218_, _19217_, _06717_);
  nor _52118_ (_19219_, _19218_, _19214_);
  nand _52119_ (_19220_, _19219_, _06751_);
  nand _52120_ (_19221_, _19220_, _19210_);
  nand _52121_ (_19222_, _19221_, _06760_);
  nand _52122_ (_19223_, _19222_, _19200_);
  nand _52123_ (_19224_, _19223_, _06731_);
  nand _52124_ (_19225_, _19224_, _19178_);
  nand _52125_ (_19226_, _19225_, _06734_);
  nand _52126_ (_19227_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand _52127_ (_19228_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nand _52128_ (_19229_, _19228_, _19227_);
  nand _52129_ (_19230_, _19229_, _06717_);
  nand _52130_ (_19231_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand _52131_ (_19232_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nand _52132_ (_19233_, _19232_, _19231_);
  nand _52133_ (_19234_, _19233_, _06716_);
  nand _52134_ (_19235_, _19234_, _19230_);
  nand _52135_ (_19236_, _19235_, _06748_);
  nand _52136_ (_19237_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand _52137_ (_19238_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nand _52138_ (_19239_, _19238_, _19237_);
  nand _52139_ (_19240_, _19239_, _06717_);
  nand _52140_ (_19241_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand _52141_ (_19242_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nand _52142_ (_19243_, _19242_, _19241_);
  nand _52143_ (_19244_, _19243_, _06716_);
  nand _52144_ (_19245_, _19244_, _19240_);
  nand _52145_ (_19246_, _19245_, _06751_);
  nand _52146_ (_19247_, _19246_, _19236_);
  nand _52147_ (_19248_, _19247_, _06761_);
  nor _52148_ (_19249_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _52149_ (_19250_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _52150_ (_19251_, _19250_, _19249_);
  nand _52151_ (_19252_, _19251_, _06717_);
  nor _52152_ (_19253_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _52153_ (_19254_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _52154_ (_19255_, _19254_, _19253_);
  nand _52155_ (_19256_, _19255_, _06716_);
  nand _52156_ (_19257_, _19256_, _19252_);
  nand _52157_ (_19258_, _19257_, _06748_);
  nor _52158_ (_19259_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _52159_ (_19260_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _52160_ (_19261_, _19260_, _19259_);
  nand _52161_ (_19262_, _19261_, _06717_);
  nor _52162_ (_19263_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor _52163_ (_19264_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _52164_ (_19265_, _19264_, _19263_);
  nand _52165_ (_19266_, _19265_, _06716_);
  nand _52166_ (_19267_, _19266_, _19262_);
  nand _52167_ (_19268_, _19267_, _06751_);
  nand _52168_ (_19269_, _19268_, _19258_);
  nand _52169_ (_19270_, _19269_, _06760_);
  nand _52170_ (_19271_, _19270_, _19248_);
  nand _52171_ (_19272_, _19271_, _06780_);
  nand _52172_ (_19273_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  nand _52173_ (_19274_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  nand _52174_ (_19275_, _19274_, _19273_);
  nand _52175_ (_19276_, _19275_, _06717_);
  nand _52176_ (_19277_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nand _52177_ (_19278_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nand _52178_ (_19279_, _19278_, _19277_);
  nand _52179_ (_19280_, _19279_, _06716_);
  nand _52180_ (_19281_, _19280_, _19276_);
  nand _52181_ (_19282_, _19281_, _06748_);
  nand _52182_ (_19283_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  nand _52183_ (_19284_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  nand _52184_ (_19285_, _19284_, _19283_);
  nand _52185_ (_19286_, _19285_, _06717_);
  nand _52186_ (_19287_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nand _52187_ (_19288_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nand _52188_ (_19289_, _19288_, _19287_);
  nand _52189_ (_19290_, _19289_, _06716_);
  nand _52190_ (_19291_, _19290_, _19286_);
  nand _52191_ (_19292_, _19291_, _06751_);
  nand _52192_ (_19293_, _19292_, _19282_);
  nand _52193_ (_19294_, _19293_, _06761_);
  nor _52194_ (_19295_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  nor _52195_ (_19296_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nor _52196_ (_19297_, _19296_, _19295_);
  nand _52197_ (_19298_, _19297_, _06717_);
  nor _52198_ (_19299_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nor _52199_ (_19300_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  nor _52200_ (_19301_, _19300_, _19299_);
  nand _52201_ (_19302_, _19301_, _06716_);
  nand _52202_ (_19303_, _19302_, _19298_);
  nand _52203_ (_19304_, _19303_, _06748_);
  nor _52204_ (_19305_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  nor _52205_ (_19306_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  nor _52206_ (_19307_, _19306_, _19305_);
  nand _52207_ (_19308_, _19307_, _06717_);
  nor _52208_ (_19309_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nor _52209_ (_19310_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nor _52210_ (_19312_, _19310_, _19309_);
  nand _52211_ (_19313_, _19312_, _06716_);
  nand _52212_ (_19314_, _19313_, _19308_);
  nand _52213_ (_19315_, _19314_, _06751_);
  nand _52214_ (_19316_, _19315_, _19304_);
  nand _52215_ (_19317_, _19316_, _06760_);
  nand _52216_ (_19318_, _19317_, _19294_);
  nand _52217_ (_19319_, _19318_, _06731_);
  nand _52218_ (_19320_, _19319_, _19272_);
  nand _52219_ (_19321_, _19320_, _06733_);
  nand _52220_ (_19322_, _19321_, _19226_);
  nor _52221_ (_19323_, _19322_, _06723_);
  nand _52222_ (_19324_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  nand _52223_ (_19325_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  nand _52224_ (_19326_, _19325_, _19324_);
  nand _52225_ (_19327_, _19326_, _06717_);
  nand _52226_ (_19328_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  nand _52227_ (_19329_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  nand _52228_ (_19330_, _19329_, _19328_);
  nand _52229_ (_19331_, _19330_, _06716_);
  nand _52230_ (_19332_, _19331_, _19327_);
  nand _52231_ (_19333_, _19332_, _06748_);
  nand _52232_ (_19334_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  nand _52233_ (_19335_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nand _52234_ (_19336_, _19335_, _19334_);
  nand _52235_ (_19337_, _19336_, _06717_);
  nand _52236_ (_19338_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nand _52237_ (_19339_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nand _52238_ (_19340_, _19339_, _19338_);
  nand _52239_ (_19341_, _19340_, _06716_);
  nand _52240_ (_19342_, _19341_, _19337_);
  nand _52241_ (_19343_, _19342_, _06751_);
  nand _52242_ (_19344_, _19343_, _19333_);
  nand _52243_ (_19345_, _19344_, _06761_);
  nor _52244_ (_19346_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  nor _52245_ (_19347_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  nor _52246_ (_19348_, _19347_, _19346_);
  nand _52247_ (_19349_, _19348_, _06716_);
  nand _52248_ (_19350_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  nand _52249_ (_19351_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nand _52250_ (_19352_, _19351_, _19350_);
  nand _52251_ (_19353_, _19352_, _06717_);
  nand _52252_ (_19354_, _19353_, _19349_);
  nand _52253_ (_19355_, _19354_, _06748_);
  nor _52254_ (_19356_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nor _52255_ (_19357_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  nor _52256_ (_19358_, _19357_, _19356_);
  nand _52257_ (_19359_, _19358_, _06716_);
  nand _52258_ (_19360_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nand _52259_ (_19361_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  nand _52260_ (_19362_, _19361_, _19360_);
  nand _52261_ (_19363_, _19362_, _06717_);
  nand _52262_ (_19364_, _19363_, _19359_);
  nand _52263_ (_19365_, _19364_, _06751_);
  nand _52264_ (_19366_, _19365_, _19355_);
  nand _52265_ (_19367_, _19366_, _06760_);
  nand _52266_ (_19368_, _19367_, _19345_);
  nand _52267_ (_19369_, _19368_, _06780_);
  nand _52268_ (_19370_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nand _52269_ (_19371_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  nand _52270_ (_19372_, _19371_, _19370_);
  nand _52271_ (_19373_, _19372_, _06717_);
  nand _52272_ (_19374_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nand _52273_ (_19375_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nand _52274_ (_19376_, _19375_, _19374_);
  nand _52275_ (_19377_, _19376_, _06716_);
  nand _52276_ (_19378_, _19377_, _19373_);
  nand _52277_ (_19379_, _19378_, _06748_);
  nand _52278_ (_19380_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  nand _52279_ (_19381_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nand _52280_ (_19382_, _19381_, _19380_);
  nand _52281_ (_19383_, _19382_, _06717_);
  nand _52282_ (_19384_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  nand _52283_ (_19385_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  nand _52284_ (_19386_, _19385_, _19384_);
  nand _52285_ (_19387_, _19386_, _06716_);
  nand _52286_ (_19388_, _19387_, _19383_);
  nand _52287_ (_19389_, _19388_, _06751_);
  nand _52288_ (_19390_, _19389_, _19379_);
  nand _52289_ (_19391_, _19390_, _06761_);
  nor _52290_ (_19392_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nor _52291_ (_19393_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nor _52292_ (_19394_, _19393_, _19392_);
  nand _52293_ (_19395_, _19394_, _06717_);
  nor _52294_ (_19396_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nor _52295_ (_19397_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  nor _52296_ (_19398_, _19397_, _19396_);
  nand _52297_ (_19399_, _19398_, _06716_);
  nand _52298_ (_19400_, _19399_, _19395_);
  nand _52299_ (_19401_, _19400_, _06748_);
  nor _52300_ (_19402_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  nor _52301_ (_19403_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nor _52302_ (_19404_, _19403_, _19402_);
  nand _52303_ (_19405_, _19404_, _06717_);
  nor _52304_ (_19406_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  nor _52305_ (_19407_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  nor _52306_ (_19408_, _19407_, _19406_);
  nand _52307_ (_19409_, _19408_, _06716_);
  nand _52308_ (_19410_, _19409_, _19405_);
  nand _52309_ (_19411_, _19410_, _06751_);
  nand _52310_ (_19412_, _19411_, _19401_);
  nand _52311_ (_19413_, _19412_, _06760_);
  nand _52312_ (_19414_, _19413_, _19391_);
  nand _52313_ (_19415_, _19414_, _06731_);
  nand _52314_ (_19416_, _19415_, _19369_);
  nand _52315_ (_19417_, _19416_, _06734_);
  nor _52316_ (_19418_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  nor _52317_ (_19419_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nor _52318_ (_19420_, _19419_, _19418_);
  nand _52319_ (_19421_, _19420_, _06717_);
  nor _52320_ (_19423_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nor _52321_ (_19424_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  nor _52322_ (_19425_, _19424_, _19423_);
  nand _52323_ (_19426_, _19425_, _06716_);
  nand _52324_ (_19427_, _19426_, _19421_);
  nand _52325_ (_19428_, _19427_, _06751_);
  nor _52326_ (_19429_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nor _52327_ (_19430_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  nor _52328_ (_19431_, _19430_, _19429_);
  nand _52329_ (_19432_, _19431_, _06717_);
  nor _52330_ (_19433_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nor _52331_ (_19434_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nor _52332_ (_19435_, _19434_, _19433_);
  nand _52333_ (_19436_, _19435_, _06716_);
  nand _52334_ (_19437_, _19436_, _19432_);
  nand _52335_ (_19438_, _19437_, _06748_);
  nand _52336_ (_19439_, _19438_, _19428_);
  nand _52337_ (_19440_, _19439_, _06760_);
  nand _52338_ (_19441_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  nand _52339_ (_19442_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  nand _52340_ (_19443_, _19442_, _19441_);
  nand _52341_ (_19444_, _19443_, _06717_);
  nand _52342_ (_19445_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  nand _52343_ (_19446_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nand _52344_ (_19447_, _19446_, _19445_);
  nand _52345_ (_19448_, _19447_, _06716_);
  nand _52346_ (_19449_, _19448_, _19444_);
  nand _52347_ (_19450_, _19449_, _06751_);
  nand _52348_ (_19451_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nand _52349_ (_19452_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  nand _52350_ (_19453_, _19452_, _19451_);
  nand _52351_ (_19454_, _19453_, _06717_);
  nand _52352_ (_19455_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nand _52353_ (_19456_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nand _52354_ (_19457_, _19456_, _19455_);
  nand _52355_ (_19458_, _19457_, _06716_);
  nand _52356_ (_19459_, _19458_, _19454_);
  nand _52357_ (_19460_, _19459_, _06748_);
  nand _52358_ (_19461_, _19460_, _19450_);
  nand _52359_ (_19462_, _19461_, _06761_);
  nand _52360_ (_19463_, _19462_, _19440_);
  nand _52361_ (_19464_, _19463_, _06731_);
  nor _52362_ (_19465_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nor _52363_ (_19466_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  nor _52364_ (_19467_, _19466_, _19465_);
  nand _52365_ (_19468_, _19467_, _06716_);
  nand _52366_ (_19469_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nand _52367_ (_19470_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  nand _52368_ (_19471_, _19470_, _19469_);
  nand _52369_ (_19472_, _19471_, _06717_);
  nand _52370_ (_19473_, _19472_, _19468_);
  nand _52371_ (_19474_, _19473_, _06751_);
  nor _52372_ (_19475_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  nor _52373_ (_19476_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  nor _52374_ (_19477_, _19476_, _19475_);
  nand _52375_ (_19478_, _19477_, _06716_);
  nand _52376_ (_19479_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  nand _52377_ (_19480_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  nand _52378_ (_19481_, _19480_, _19479_);
  nand _52379_ (_19482_, _19481_, _06717_);
  nand _52380_ (_19483_, _19482_, _19478_);
  nand _52381_ (_19484_, _19483_, _06748_);
  nand _52382_ (_19485_, _19484_, _19474_);
  nand _52383_ (_19486_, _19485_, _06760_);
  nand _52384_ (_19487_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  nand _52385_ (_19488_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  nand _52386_ (_19489_, _19488_, _19487_);
  nand _52387_ (_19490_, _19489_, _06717_);
  nand _52388_ (_19491_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  nand _52389_ (_19492_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  nand _52390_ (_19493_, _19492_, _19491_);
  nand _52391_ (_19494_, _19493_, _06716_);
  nand _52392_ (_19495_, _19494_, _19490_);
  nand _52393_ (_19496_, _19495_, _06751_);
  nand _52394_ (_19497_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  nand _52395_ (_19498_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nand _52396_ (_19499_, _19498_, _19497_);
  nand _52397_ (_19500_, _19499_, _06717_);
  nand _52398_ (_19501_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nand _52399_ (_19502_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  nand _52400_ (_19504_, _19502_, _19501_);
  nand _52401_ (_19505_, _19504_, _06716_);
  nand _52402_ (_19506_, _19505_, _19500_);
  nand _52403_ (_19507_, _19506_, _06748_);
  nand _52404_ (_19508_, _19507_, _19496_);
  nand _52405_ (_19509_, _19508_, _06761_);
  nand _52406_ (_19510_, _19509_, _19486_);
  nand _52407_ (_19511_, _19510_, _06780_);
  nand _52408_ (_19512_, _19511_, _19464_);
  nand _52409_ (_19513_, _19512_, _06733_);
  nand _52410_ (_19514_, _19513_, _19417_);
  nor _52411_ (_19515_, _19514_, _13106_);
  nor _52412_ (_19516_, _19515_, _19323_);
  nor _52413_ (_19517_, _19516_, _25929_);
  nand _52414_ (_19518_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  nand _52415_ (_19519_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nand _52416_ (_19520_, _19519_, _19518_);
  nand _52417_ (_19521_, _19520_, _06717_);
  nand _52418_ (_19522_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nand _52419_ (_19523_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  nand _52420_ (_19524_, _19523_, _19522_);
  nand _52421_ (_19525_, _19524_, _06716_);
  nand _52422_ (_19526_, _19525_, _19521_);
  nand _52423_ (_19527_, _19526_, _06748_);
  nand _52424_ (_19528_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nand _52425_ (_19529_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nand _52426_ (_19530_, _19529_, _19528_);
  nand _52427_ (_19531_, _19530_, _06717_);
  nand _52428_ (_19532_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  nand _52429_ (_19533_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  nand _52430_ (_19534_, _19533_, _19532_);
  nand _52431_ (_19535_, _19534_, _06716_);
  nand _52432_ (_19536_, _19535_, _19531_);
  nand _52433_ (_19537_, _19536_, _06751_);
  nand _52434_ (_19538_, _19537_, _19527_);
  nand _52435_ (_19539_, _19538_, _06761_);
  nor _52436_ (_19540_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nor _52437_ (_19541_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  nor _52438_ (_19542_, _19541_, _19540_);
  nand _52439_ (_19543_, _19542_, _06716_);
  nand _52440_ (_19544_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nand _52441_ (_19545_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  nand _52442_ (_19546_, _19545_, _19544_);
  nand _52443_ (_19547_, _19546_, _06717_);
  nand _52444_ (_19548_, _19547_, _19543_);
  nand _52445_ (_19549_, _19548_, _06748_);
  nor _52446_ (_19550_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nor _52447_ (_19551_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  nor _52448_ (_19552_, _19551_, _19550_);
  nand _52449_ (_19553_, _19552_, _06716_);
  nand _52450_ (_19555_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  nand _52451_ (_19556_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  nand _52452_ (_19557_, _19556_, _19555_);
  nand _52453_ (_19558_, _19557_, _06717_);
  nand _52454_ (_19559_, _19558_, _19553_);
  nand _52455_ (_19560_, _19559_, _06751_);
  nand _52456_ (_19561_, _19560_, _19549_);
  nand _52457_ (_19562_, _19561_, _06760_);
  nand _52458_ (_19563_, _19562_, _19539_);
  nand _52459_ (_19564_, _19563_, _06780_);
  nand _52460_ (_19565_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  nand _52461_ (_19566_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nand _52462_ (_19567_, _19566_, _19565_);
  nand _52463_ (_19568_, _19567_, _06717_);
  nand _52464_ (_19569_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nand _52465_ (_19570_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  nand _52466_ (_19571_, _19570_, _19569_);
  nand _52467_ (_19572_, _19571_, _06716_);
  nand _52468_ (_19573_, _19572_, _19568_);
  nand _52469_ (_19574_, _19573_, _06748_);
  nand _52470_ (_19575_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  nand _52471_ (_19576_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  nand _52472_ (_19577_, _19576_, _19575_);
  nand _52473_ (_19578_, _19577_, _06717_);
  nand _52474_ (_19579_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nand _52475_ (_19580_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nand _52476_ (_19581_, _19580_, _19579_);
  nand _52477_ (_19582_, _19581_, _06716_);
  nand _52478_ (_19583_, _19582_, _19578_);
  nand _52479_ (_19584_, _19583_, _06751_);
  nand _52480_ (_19585_, _19584_, _19574_);
  nand _52481_ (_19586_, _19585_, _06761_);
  nor _52482_ (_19587_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  nor _52483_ (_19588_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nor _52484_ (_19589_, _19588_, _19587_);
  nand _52485_ (_19590_, _19589_, _06717_);
  nor _52486_ (_19591_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nor _52487_ (_19592_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  nor _52488_ (_19593_, _19592_, _19591_);
  nand _52489_ (_19594_, _19593_, _06716_);
  nand _52490_ (_19595_, _19594_, _19590_);
  nand _52491_ (_19596_, _19595_, _06748_);
  nor _52492_ (_19597_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  nor _52493_ (_19598_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nor _52494_ (_19599_, _19598_, _19597_);
  nand _52495_ (_19600_, _19599_, _06717_);
  nor _52496_ (_19601_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nor _52497_ (_19602_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  nor _52498_ (_19603_, _19602_, _19601_);
  nand _52499_ (_19604_, _19603_, _06716_);
  nand _52500_ (_19606_, _19604_, _19600_);
  nand _52501_ (_19607_, _19606_, _06751_);
  nand _52502_ (_19608_, _19607_, _19596_);
  nand _52503_ (_19609_, _19608_, _06760_);
  nand _52504_ (_19610_, _19609_, _19586_);
  nand _52505_ (_19611_, _19610_, _06731_);
  nand _52506_ (_19612_, _19611_, _19564_);
  nand _52507_ (_19613_, _19612_, _06733_);
  nand _52508_ (_19614_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  nand _52509_ (_19615_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nand _52510_ (_19616_, _19615_, _19614_);
  nand _52511_ (_19617_, _19616_, _06717_);
  nand _52512_ (_19618_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nand _52513_ (_19619_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  nand _52514_ (_19620_, _19619_, _19618_);
  nand _52515_ (_19621_, _19620_, _06716_);
  nand _52516_ (_19622_, _19621_, _19617_);
  nand _52517_ (_19623_, _19622_, _06748_);
  nand _52518_ (_19624_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  nand _52519_ (_19625_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  nand _52520_ (_19626_, _19625_, _19624_);
  nand _52521_ (_19627_, _19626_, _06717_);
  nand _52522_ (_19628_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  nand _52523_ (_19629_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  nand _52524_ (_19630_, _19629_, _19628_);
  nand _52525_ (_19631_, _19630_, _06716_);
  nand _52526_ (_19632_, _19631_, _19627_);
  nand _52527_ (_19633_, _19632_, _06751_);
  nand _52528_ (_19634_, _19633_, _19623_);
  nand _52529_ (_19635_, _19634_, _06761_);
  nor _52530_ (_19636_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  nor _52531_ (_19637_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  nor _52532_ (_19638_, _19637_, _19636_);
  nand _52533_ (_19639_, _19638_, _06717_);
  nor _52534_ (_19640_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  nor _52535_ (_19641_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nor _52536_ (_19642_, _19641_, _19640_);
  nand _52537_ (_19643_, _19642_, _06716_);
  nand _52538_ (_19644_, _19643_, _19639_);
  nand _52539_ (_19645_, _19644_, _06748_);
  nor _52540_ (_19646_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nor _52541_ (_19647_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nor _52542_ (_19648_, _19647_, _19646_);
  nand _52543_ (_19649_, _19648_, _06717_);
  nor _52544_ (_19650_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nor _52545_ (_19651_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  nor _52546_ (_19652_, _19651_, _19650_);
  nand _52547_ (_19653_, _19652_, _06716_);
  nand _52548_ (_19654_, _19653_, _19649_);
  nand _52549_ (_19655_, _19654_, _06751_);
  nand _52550_ (_19657_, _19655_, _19645_);
  nand _52551_ (_19658_, _19657_, _06760_);
  nand _52552_ (_19659_, _19658_, _19635_);
  nand _52553_ (_19660_, _19659_, _06731_);
  nand _52554_ (_19661_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nand _52555_ (_19662_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  nand _52556_ (_19663_, _19662_, _19661_);
  nand _52557_ (_19664_, _19663_, _06717_);
  nand _52558_ (_19665_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  nand _52559_ (_19666_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nand _52560_ (_19667_, _19666_, _19665_);
  nand _52561_ (_19668_, _19667_, _06716_);
  nand _52562_ (_19669_, _19668_, _19664_);
  nand _52563_ (_19670_, _19669_, _06748_);
  nand _52564_ (_19671_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  nand _52565_ (_19672_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  nand _52566_ (_19673_, _19672_, _19671_);
  nand _52567_ (_19674_, _19673_, _06717_);
  nand _52568_ (_19675_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nand _52569_ (_19676_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  nand _52570_ (_19677_, _19676_, _19675_);
  nand _52571_ (_19678_, _19677_, _06716_);
  nand _52572_ (_19679_, _19678_, _19674_);
  nand _52573_ (_19680_, _19679_, _06751_);
  nand _52574_ (_19681_, _19680_, _19670_);
  nand _52575_ (_19682_, _19681_, _06761_);
  nor _52576_ (_19683_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  nor _52577_ (_19684_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nor _52578_ (_19685_, _19684_, _19683_);
  nand _52579_ (_19686_, _19685_, _06716_);
  nand _52580_ (_19687_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nand _52581_ (_19688_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nand _52582_ (_19689_, _19688_, _19687_);
  nand _52583_ (_19690_, _19689_, _06717_);
  nand _52584_ (_19691_, _19690_, _19686_);
  nand _52585_ (_19692_, _19691_, _06748_);
  nor _52586_ (_19693_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nor _52587_ (_19694_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nor _52588_ (_19695_, _19694_, _19693_);
  nand _52589_ (_19696_, _19695_, _06716_);
  nand _52590_ (_19697_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  nand _52591_ (_19698_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  nand _52592_ (_19699_, _19698_, _19697_);
  nand _52593_ (_19700_, _19699_, _06717_);
  nand _52594_ (_19701_, _19700_, _19696_);
  nand _52595_ (_19702_, _19701_, _06751_);
  nand _52596_ (_19703_, _19702_, _19692_);
  nand _52597_ (_19704_, _19703_, _06760_);
  nand _52598_ (_19705_, _19704_, _19682_);
  nand _52599_ (_19706_, _19705_, _06780_);
  nand _52600_ (_19707_, _19706_, _19660_);
  nand _52601_ (_19708_, _19707_, _06734_);
  nand _52602_ (_19709_, _19708_, _19613_);
  nor _52603_ (_19710_, _19709_, _06723_);
  nand _52604_ (_19711_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nand _52605_ (_19712_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  nand _52606_ (_19713_, _19712_, _19711_);
  nand _52607_ (_19714_, _19713_, _06716_);
  nand _52608_ (_19715_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  nand _52609_ (_19716_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nand _52610_ (_19718_, _19716_, _19715_);
  nand _52611_ (_19719_, _19718_, _06717_);
  nand _52612_ (_19720_, _19719_, _19714_);
  nand _52613_ (_19721_, _19720_, _06748_);
  nand _52614_ (_19722_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nand _52615_ (_19723_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  nand _52616_ (_19724_, _19723_, _19722_);
  nand _52617_ (_19725_, _19724_, _06716_);
  nand _52618_ (_19726_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  nand _52619_ (_19727_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nand _52620_ (_19728_, _19727_, _19726_);
  nand _52621_ (_19729_, _19728_, _06717_);
  nand _52622_ (_19730_, _19729_, _19725_);
  nand _52623_ (_19731_, _19730_, _06751_);
  nand _52624_ (_19732_, _19731_, _19721_);
  nand _52625_ (_19733_, _19732_, _06761_);
  nand _52626_ (_19734_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nand _52627_ (_19735_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  nand _52628_ (_19736_, _19735_, _19734_);
  nand _52629_ (_19737_, _19736_, _06717_);
  nor _52630_ (_19738_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  nor _52631_ (_19739_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  nor _52632_ (_19740_, _19739_, _19738_);
  nand _52633_ (_19741_, _19740_, _06716_);
  nand _52634_ (_19742_, _19741_, _19737_);
  nand _52635_ (_19743_, _19742_, _06748_);
  nand _52636_ (_19744_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  nand _52637_ (_19745_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nand _52638_ (_19746_, _19745_, _19744_);
  nand _52639_ (_19747_, _19746_, _06717_);
  nor _52640_ (_19748_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  nor _52641_ (_19749_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nor _52642_ (_19750_, _19749_, _19748_);
  nand _52643_ (_19751_, _19750_, _06716_);
  nand _52644_ (_19752_, _19751_, _19747_);
  nand _52645_ (_19753_, _19752_, _06751_);
  nand _52646_ (_19754_, _19753_, _19743_);
  nand _52647_ (_19755_, _19754_, _06760_);
  nand _52648_ (_19756_, _19755_, _19733_);
  nand _52649_ (_19757_, _19756_, _06780_);
  nand _52650_ (_19758_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  nand _52651_ (_19759_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nand _52652_ (_19760_, _19759_, _19758_);
  nand _52653_ (_19761_, _19760_, _06717_);
  nand _52654_ (_19762_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nand _52655_ (_19763_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  nand _52656_ (_19764_, _19763_, _19762_);
  nand _52657_ (_19765_, _19764_, _06716_);
  nand _52658_ (_19766_, _19765_, _19761_);
  nand _52659_ (_19767_, _19766_, _06748_);
  nand _52660_ (_19768_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  nand _52661_ (_19769_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  nand _52662_ (_19770_, _19769_, _19768_);
  nand _52663_ (_19771_, _19770_, _06717_);
  nand _52664_ (_19772_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  nand _52665_ (_19773_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nand _52666_ (_19774_, _19773_, _19772_);
  nand _52667_ (_19775_, _19774_, _06716_);
  nand _52668_ (_19776_, _19775_, _19771_);
  nand _52669_ (_19777_, _19776_, _06751_);
  nand _52670_ (_19778_, _19777_, _19767_);
  nand _52671_ (_19779_, _19778_, _06761_);
  nor _52672_ (_19780_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nor _52673_ (_19781_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  nor _52674_ (_19782_, _19781_, _19780_);
  nand _52675_ (_19783_, _19782_, _06717_);
  nor _52676_ (_19784_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  nor _52677_ (_19785_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nor _52678_ (_19786_, _19785_, _19784_);
  nand _52679_ (_19787_, _19786_, _06716_);
  nand _52680_ (_19788_, _19787_, _19783_);
  nand _52681_ (_19789_, _19788_, _06748_);
  nor _52682_ (_19790_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nor _52683_ (_19791_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  nor _52684_ (_19792_, _19791_, _19790_);
  nor _52685_ (_19793_, _19792_, _06716_);
  nor _52686_ (_19794_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  nor _52687_ (_19795_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  nor _52688_ (_19796_, _19795_, _19794_);
  nor _52689_ (_19797_, _19796_, _06717_);
  nor _52690_ (_19798_, _19797_, _19793_);
  nand _52691_ (_19799_, _19798_, _06751_);
  nand _52692_ (_19800_, _19799_, _19789_);
  nand _52693_ (_19801_, _19800_, _06760_);
  nand _52694_ (_19802_, _19801_, _19779_);
  nand _52695_ (_19803_, _19802_, _06731_);
  nand _52696_ (_19804_, _19803_, _19757_);
  nand _52697_ (_19805_, _19804_, _06734_);
  nand _52698_ (_19806_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  nand _52699_ (_19807_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  nand _52700_ (_19808_, _19807_, _19806_);
  nand _52701_ (_19809_, _19808_, _06717_);
  nand _52702_ (_19810_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nand _52703_ (_19811_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nand _52704_ (_19812_, _19811_, _19810_);
  nand _52705_ (_19813_, _19812_, _06716_);
  nand _52706_ (_19814_, _19813_, _19809_);
  nand _52707_ (_19815_, _19814_, _06748_);
  nand _52708_ (_19816_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  nand _52709_ (_19817_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nand _52710_ (_19818_, _19817_, _19816_);
  nand _52711_ (_19819_, _19818_, _06717_);
  nand _52712_ (_19820_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  nand _52713_ (_19821_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  nand _52714_ (_19822_, _19821_, _19820_);
  nand _52715_ (_19823_, _19822_, _06716_);
  nand _52716_ (_19824_, _19823_, _19819_);
  nand _52717_ (_19825_, _19824_, _06751_);
  nand _52718_ (_19826_, _19825_, _19815_);
  nand _52719_ (_19827_, _19826_, _06761_);
  nor _52720_ (_19828_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  nor _52721_ (_19829_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nor _52722_ (_19830_, _19829_, _19828_);
  nand _52723_ (_19831_, _19830_, _06717_);
  nor _52724_ (_19832_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nor _52725_ (_19833_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  nor _52726_ (_19834_, _19833_, _19832_);
  nand _52727_ (_19835_, _19834_, _06716_);
  nand _52728_ (_19836_, _19835_, _19831_);
  nand _52729_ (_19837_, _19836_, _06748_);
  nor _52730_ (_19838_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  nor _52731_ (_19839_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  nor _52732_ (_19840_, _19839_, _19838_);
  nand _52733_ (_19841_, _19840_, _06717_);
  nor _52734_ (_19842_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  nor _52735_ (_19843_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nor _52736_ (_19844_, _19843_, _19842_);
  nand _52737_ (_19845_, _19844_, _06716_);
  nand _52738_ (_19846_, _19845_, _19841_);
  nand _52739_ (_19847_, _19846_, _06751_);
  nand _52740_ (_19848_, _19847_, _19837_);
  nand _52741_ (_19849_, _19848_, _06760_);
  nand _52742_ (_19850_, _19849_, _19827_);
  nand _52743_ (_19851_, _19850_, _06731_);
  nand _52744_ (_19852_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  nand _52745_ (_19853_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  nand _52746_ (_19854_, _19853_, _19852_);
  nand _52747_ (_19855_, _19854_, _06717_);
  nand _52748_ (_19856_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  nand _52749_ (_19857_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nand _52750_ (_19858_, _19857_, _19856_);
  nand _52751_ (_19859_, _19858_, _06716_);
  nand _52752_ (_19860_, _19859_, _19855_);
  nand _52753_ (_19861_, _19860_, _06748_);
  nand _52754_ (_19862_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nand _52755_ (_19863_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  nand _52756_ (_19864_, _19863_, _19862_);
  nand _52757_ (_19865_, _19864_, _06717_);
  nand _52758_ (_19866_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  nand _52759_ (_19867_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nand _52760_ (_19868_, _19867_, _19866_);
  nand _52761_ (_19869_, _19868_, _06716_);
  nand _52762_ (_19870_, _19869_, _19865_);
  nand _52763_ (_19871_, _19870_, _06751_);
  nand _52764_ (_19872_, _19871_, _19861_);
  nand _52765_ (_19873_, _19872_, _06761_);
  nor _52766_ (_19874_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nor _52767_ (_19875_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  nor _52768_ (_19876_, _19875_, _19874_);
  nand _52769_ (_19877_, _19876_, _06717_);
  nor _52770_ (_19878_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  nor _52771_ (_19879_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  nor _52772_ (_19880_, _19879_, _19878_);
  nand _52773_ (_19881_, _19880_, _06716_);
  nand _52774_ (_19882_, _19881_, _19877_);
  nand _52775_ (_19883_, _19882_, _06748_);
  nor _52776_ (_19884_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nor _52777_ (_19885_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  nor _52778_ (_19886_, _19885_, _19884_);
  nand _52779_ (_19887_, _19886_, _06717_);
  nor _52780_ (_19888_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nor _52781_ (_19889_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  nor _52782_ (_19890_, _19889_, _19888_);
  nand _52783_ (_19891_, _19890_, _06716_);
  nand _52784_ (_19892_, _19891_, _19887_);
  nand _52785_ (_19893_, _19892_, _06751_);
  nand _52786_ (_19894_, _19893_, _19883_);
  nand _52787_ (_19895_, _19894_, _06760_);
  nand _52788_ (_19896_, _19895_, _19873_);
  nand _52789_ (_19897_, _19896_, _06780_);
  nand _52790_ (_19898_, _19897_, _19851_);
  nand _52791_ (_19899_, _19898_, _06733_);
  nand _52792_ (_19900_, _19899_, _19805_);
  nor _52793_ (_19901_, _19900_, _13106_);
  nor _52794_ (_19902_, _19901_, _19710_);
  nor _52795_ (_19903_, _19902_, _25843_);
  nor _52796_ (_19904_, _19903_, _19517_);
  nor _52797_ (_19905_, _19904_, _13105_);
  nand _52798_ (_19906_, _13105_, _24225_);
  nand _52799_ (_19907_, _19906_, _26487_);
  nor _52800_ (_09502_, _19907_, _19905_);
  nand _52801_ (_19908_, _05739_, _24927_);
  nand _52802_ (_19909_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  nand _52803_ (_09529_, _19909_, _19908_);
  nand _52804_ (_19910_, _12688_, _24927_);
  nand _52805_ (_19911_, _12690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nand _52806_ (_09546_, _19911_, _19910_);
  nand _52807_ (_19912_, _11855_, _25039_);
  nand _52808_ (_19913_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  nand _52809_ (_28289_, _19913_, _19912_);
  nand _52810_ (_19914_, _19119_, _24789_);
  nand _52811_ (_19915_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  nand _52812_ (_09578_, _19915_, _19914_);
  nand _52813_ (_19916_, _11855_, _25150_);
  nand _52814_ (_19917_, _11857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nand _52815_ (_28290_, _19917_, _19916_);
  nand _52816_ (_19918_, _11848_, _24830_);
  nand _52817_ (_19919_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  nand _52818_ (_28291_, _19919_, _19918_);
  nand _52819_ (_19920_, _09944_, _25039_);
  nand _52820_ (_19922_, _09946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nand _52821_ (_09621_, _19922_, _19920_);
  nand _52822_ (_19923_, _18946_, _28096_);
  nand _52823_ (_19924_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nand _52824_ (_09636_, _19924_, _19923_);
  nand _52825_ (_19925_, _11848_, _25099_);
  nand _52826_ (_19926_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  nand _52827_ (_09638_, _19926_, _19925_);
  nor _52828_ (_19927_, _00219_, _26260_);
  nand _52829_ (_19928_, _19927_, _23940_);
  nor _52830_ (_19929_, _19928_, _25723_);
  not _52831_ (_19930_, _19929_);
  nor _52832_ (_19931_, _19930_, _24716_);
  nor _52833_ (_19932_, _19929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor _52834_ (_19933_, _19932_, _19931_);
  nor _52835_ (_19934_, _19933_, _00374_);
  nand _52836_ (_19935_, _00374_, _24820_);
  nand _52837_ (_19936_, _19935_, _26487_);
  nor _52838_ (_09641_, _19936_, _19934_);
  nor _52839_ (_19937_, _19928_, _00263_);
  not _52840_ (_19938_, _19937_);
  nor _52841_ (_19939_, _19938_, _24716_);
  nor _52842_ (_19940_, _19937_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _52843_ (_19941_, _19940_, _19939_);
  nor _52844_ (_19942_, _19941_, _00374_);
  nand _52845_ (_19943_, _00236_, _25195_);
  nand _52846_ (_19944_, _19943_, _26487_);
  nor _52847_ (_09643_, _19944_, _19942_);
  nor _52848_ (_19945_, _19928_, _00276_);
  not _52849_ (_19946_, _19945_);
  nor _52850_ (_19947_, _19946_, _24716_);
  nor _52851_ (_19948_, _19945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  nor _52852_ (_19949_, _19948_, _19947_);
  nor _52853_ (_19950_, _19949_, _00374_);
  nand _52854_ (_19951_, _00236_, _25703_);
  nand _52855_ (_19952_, _19951_, _26487_);
  nor _52856_ (_09646_, _19952_, _19950_);
  not _52857_ (_19953_, _00153_);
  nand _52858_ (_19954_, _19953_, _00216_);
  nand _52859_ (_19955_, _19954_, _05060_);
  nor _52860_ (_19956_, _19955_, _00223_);
  nand _52861_ (_19957_, _01666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _52862_ (_19958_, _19957_, _00223_);
  nor _52863_ (_19959_, _19958_, _07866_);
  nor _52864_ (_19960_, _19959_, _19956_);
  nor _52865_ (_19961_, _19960_, _00236_);
  nand _52866_ (_19962_, _00236_, _25140_);
  nand _52867_ (_19963_, _19962_, _26487_);
  nor _52868_ (_09648_, _19963_, _19961_);
  nand _52869_ (_19964_, _00223_, _03356_);
  nand _52870_ (_19965_, _19964_, _05076_);
  nand _52871_ (_19966_, _19965_, _00375_);
  nor _52872_ (_19967_, _19964_, _24716_);
  nor _52873_ (_19968_, _19967_, _19966_);
  nor _52874_ (_19969_, _00375_, _26096_);
  nor _52875_ (_19970_, _19969_, _19968_);
  nor _52876_ (_09651_, _19970_, rst);
  nand _52877_ (_19971_, _10226_, _25039_);
  nand _52878_ (_19972_, _10230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand _52879_ (_09667_, _19972_, _19971_);
  nand _52880_ (_19974_, _18946_, _25203_);
  nand _52881_ (_19975_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  nand _52882_ (_28326_, _19975_, _19974_);
  nand _52883_ (_19976_, _12096_, _24789_);
  nand _52884_ (_19977_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  nand _52885_ (_09683_, _19977_, _19976_);
  nand _52886_ (_19978_, _19119_, _25150_);
  nand _52887_ (_19979_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nand _52888_ (_09691_, _19979_, _19978_);
  nand _52889_ (_19980_, _11848_, _25203_);
  nand _52890_ (_19981_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nand _52891_ (_09693_, _19981_, _19980_);
  nand _52892_ (_19982_, _11848_, _24927_);
  nand _52893_ (_19983_, _11850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  nand _52894_ (_09695_, _19983_, _19982_);
  nand _52895_ (_09702_, _26396_, _26487_);
  nand _52896_ (_19984_, _04251_, _25099_);
  nand _52897_ (_19985_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  nand _52898_ (_09707_, _19985_, _19984_);
  nor _52899_ (_19986_, _18662_, _07977_);
  not _52900_ (_19988_, _19986_);
  nor _52901_ (_19989_, _19988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _52902_ (_19990_, _19986_, _18310_);
  nor _52903_ (_19991_, _19990_, _19989_);
  nor _52904_ (_19992_, _19991_, _07948_);
  nand _52905_ (_19993_, _07948_, _24821_);
  nand _52906_ (_19994_, _19993_, _18306_);
  nor _52907_ (_19995_, _19994_, _19992_);
  nand _52908_ (_19996_, _07941_, _18310_);
  nand _52909_ (_19997_, _19996_, _26487_);
  nor _52910_ (_09714_, _19997_, _19995_);
  nand _52911_ (_19998_, _10222_, _25203_);
  nand _52912_ (_19999_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nand _52913_ (_09725_, _19999_, _19998_);
  nand _52914_ (_20000_, _12710_, _24830_);
  nand _52915_ (_20001_, _12712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  nand _52916_ (_09728_, _20001_, _20000_);
  nor _52917_ (_09732_, _26070_, rst);
  nand _52918_ (_20002_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  nand _52919_ (_20003_, _08324_, _25099_);
  nand _52920_ (_09742_, _20003_, _20002_);
  nand _52921_ (_20004_, _00955_, _24927_);
  nand _52922_ (_20005_, _00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  nand _52923_ (_09759_, _20005_, _20004_);
  nor _52924_ (_20006_, _05481_, _04760_);
  not _52925_ (_20007_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor _52926_ (_20008_, _25726_, _25627_);
  nand _52927_ (_20009_, _20008_, _00444_);
  nand _52928_ (_20010_, _20009_, _20007_);
  nand _52929_ (_20011_, _20010_, _05481_);
  nor _52930_ (_20012_, _20009_, _02415_);
  nor _52931_ (_20013_, _20012_, _20011_);
  nor _52932_ (_20014_, _20013_, _20006_);
  nor _52933_ (_09770_, _20014_, rst);
  nand _52934_ (_09774_, _26440_, _26487_);
  nand _52935_ (_09777_, _26277_, _26487_);
  nand _52936_ (_20015_, _00394_, _25039_);
  nand _52937_ (_20016_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  nand _52938_ (_09781_, _20016_, _20015_);
  nand _52939_ (_20017_, _18131_, _24927_);
  nand _52940_ (_20018_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  nand _52941_ (_09791_, _20018_, _20017_);
  nand _52942_ (_20019_, _28059_, _25039_);
  nand _52943_ (_20020_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  nand _52944_ (_09801_, _20020_, _20019_);
  nand _52945_ (_20021_, _28059_, _24830_);
  nand _52946_ (_20022_, _28061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nand _52947_ (_09805_, _20022_, _20021_);
  nand _52948_ (_20023_, _01153_, _24927_);
  nand _52949_ (_20024_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  nand _52950_ (_09806_, _20024_, _20023_);
  nand _52951_ (_20025_, _11839_, _25099_);
  nand _52952_ (_20026_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  nand _52953_ (_09809_, _20026_, _20025_);
  not _52954_ (_20027_, _20008_);
  nor _52955_ (_20028_, _20027_, _00276_);
  nor _52956_ (_20029_, _20028_, _05469_);
  nor _52957_ (_20030_, _20029_, _02415_);
  not _52958_ (_20031_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand _52959_ (_20032_, _20029_, _20031_);
  nand _52960_ (_20033_, _20032_, _26487_);
  nor _52961_ (_09814_, _20033_, _20030_);
  nand _52962_ (_20034_, _11633_, _24830_);
  nand _52963_ (_20035_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  nand _52964_ (_28374_, _20035_, _20034_);
  nand _52965_ (_20036_, _10222_, _25099_);
  nand _52966_ (_20037_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nand _52967_ (_09817_, _20037_, _20036_);
  nand _52968_ (_20038_, _03894_, _25150_);
  nand _52969_ (_20039_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  nand _52970_ (_09820_, _20039_, _20038_);
  nand _52971_ (_20040_, _25099_, _24985_);
  nand _52972_ (_20041_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nand _52973_ (_09829_, _20041_, _20040_);
  nand _52974_ (_20042_, _19068_, _25150_);
  nand _52975_ (_20043_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  nand _52976_ (_09831_, _20043_, _20042_);
  nand _52977_ (_20044_, _18131_, _25039_);
  nand _52978_ (_20045_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  nand _52979_ (_09838_, _20045_, _20044_);
  nand _52980_ (_20046_, _10222_, _24927_);
  nand _52981_ (_20047_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  nand _52982_ (_09849_, _20047_, _20046_);
  nand _52983_ (_20048_, _11839_, _25203_);
  nand _52984_ (_20049_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nand _52985_ (_09855_, _20049_, _20048_);
  nor _52986_ (_09861_, _25938_, rst);
  nand _52987_ (_20050_, _18131_, _25203_);
  nand _52988_ (_20051_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nand _52989_ (_09864_, _20051_, _20050_);
  nand _52990_ (_20052_, _19024_, _25099_);
  nand _52991_ (_20053_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nand _52992_ (_28324_, _20053_, _20052_);
  nor _52993_ (_09876_, _26052_, rst);
  nand _52994_ (_20054_, _18131_, _28096_);
  nand _52995_ (_20055_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  nand _52996_ (_28266_, _20055_, _20054_);
  nand _52997_ (_20056_, _18157_, _24927_);
  nand _52998_ (_20057_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  nand _52999_ (_09887_, _20057_, _20056_);
  nor _53000_ (_09889_, _25892_, rst);
  nand _53001_ (_20058_, _07908_, _25203_);
  nand _53002_ (_20059_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  nand _53003_ (_09898_, _20059_, _20058_);
  nand _53004_ (_20060_, _07908_, _24927_);
  nand _53005_ (_20061_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  nand _53006_ (_09900_, _20061_, _20060_);
  nand _53007_ (_20062_, _11633_, _25039_);
  nand _53008_ (_20063_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  nand _53009_ (_09902_, _20063_, _20062_);
  nor _53010_ (_20064_, _05481_, _02802_);
  not _53011_ (_20065_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand _53012_ (_20066_, _20009_, _20065_);
  nand _53013_ (_20067_, _20066_, _05481_);
  nor _53014_ (_20068_, _20009_, _02761_);
  nor _53015_ (_20069_, _20068_, _20067_);
  nor _53016_ (_20070_, _20069_, _20064_);
  nor _53017_ (_09911_, _20070_, rst);
  nand _53018_ (_20071_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nand _53019_ (_20072_, _04601_, _25203_);
  nand _53020_ (_09913_, _20072_, _20071_);
  nand _53021_ (_20073_, _24985_, _24927_);
  nand _53022_ (_20074_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  nand _53023_ (_28370_, _20074_, _20073_);
  nand _53024_ (_20075_, _11633_, _25099_);
  nand _53025_ (_20076_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  nand _53026_ (_09926_, _20076_, _20075_);
  nand _53027_ (_20077_, _04251_, _24927_);
  nand _53028_ (_20078_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  nand _53029_ (_28373_, _20078_, _20077_);
  nand _53030_ (_20079_, _10222_, _24789_);
  nand _53031_ (_20080_, _10224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  nand _53032_ (_28372_, _20080_, _20079_);
  nor _53033_ (_20081_, _20029_, _01974_);
  not _53034_ (_20082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _53035_ (_20083_, _20029_, _20082_);
  nand _53036_ (_20084_, _20083_, _26487_);
  nor _53037_ (_09935_, _20084_, _20081_);
  nand _53038_ (_20085_, _00394_, _24830_);
  nand _53039_ (_20086_, _00396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nand _53040_ (_09948_, _20086_, _20085_);
  nor _53041_ (_20087_, _05481_, _02478_);
  nand _53042_ (_20088_, _20009_, _05931_);
  nand _53043_ (_20089_, _20088_, _05481_);
  nor _53044_ (_20090_, _20009_, _01974_);
  nor _53045_ (_20091_, _20090_, _20089_);
  nor _53046_ (_20092_, _20091_, _20087_);
  nor _53047_ (_09965_, _20092_, rst);
  nor _53048_ (_20093_, _20029_, _02620_);
  not _53049_ (_20094_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand _53050_ (_20095_, _20029_, _20094_);
  nand _53051_ (_20096_, _20095_, _26487_);
  nor _53052_ (_09967_, _20096_, _20093_);
  nand _53053_ (_20097_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  nand _53054_ (_20098_, _04601_, _24789_);
  nand _53055_ (_09972_, _20098_, _20097_);
  nand _53056_ (_20099_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nand _53057_ (_20100_, _08324_, _28096_);
  nand _53058_ (_09980_, _20100_, _20099_);
  nand _53059_ (_20101_, _11839_, _25039_);
  nand _53060_ (_20102_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nand _53061_ (_28292_, _20102_, _20101_);
  nand _53062_ (_20103_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  nand _53063_ (_20104_, _08324_, _24927_);
  nand _53064_ (_28306_, _20104_, _20103_);
  nand _53065_ (_20105_, _28081_, _24927_);
  nand _53066_ (_20106_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  nand _53067_ (_09992_, _20106_, _20105_);
  nand _53068_ (_20107_, _01398_, _24789_);
  nand _53069_ (_20108_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  nand _53070_ (_09995_, _20108_, _20107_);
  nand _53071_ (_20110_, _01398_, _25099_);
  nand _53072_ (_20111_, _01400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  nand _53073_ (_09997_, _20111_, _20110_);
  nand _53074_ (_20112_, _07423_, _25203_);
  nand _53075_ (_20113_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nand _53076_ (_09999_, _20113_, _20112_);
  nor _53077_ (_20114_, _26135_, _24490_);
  nor _53078_ (_20115_, _20114_, _00226_);
  nor _53079_ (_20116_, _20115_, _26262_);
  not _53080_ (_20117_, _25729_);
  nand _53081_ (_20118_, _26253_, _24717_);
  nor _53082_ (_20119_, _26253_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _53083_ (_20120_, _20119_, _26261_);
  nand _53084_ (_20121_, _20120_, _20118_);
  nand _53085_ (_20122_, _20121_, _20117_);
  nor _53086_ (_20123_, _20122_, _20116_);
  nand _53087_ (_20124_, _25729_, _25625_);
  nand _53088_ (_20125_, _20124_, _26487_);
  nor _53089_ (_10002_, _20125_, _20123_);
  nand _53090_ (_20126_, _11839_, _24789_);
  nand _53091_ (_20127_, _11841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  nand _53092_ (_10005_, _20127_, _20126_);
  nor _53093_ (_20128_, _20029_, _02373_);
  not _53094_ (_20129_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand _53095_ (_20130_, _20029_, _20129_);
  nand _53096_ (_20131_, _20130_, _26487_);
  nor _53097_ (_10007_, _20131_, _20128_);
  nor _53098_ (_20132_, _20029_, _02096_);
  not _53099_ (_20133_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand _53100_ (_20134_, _20029_, _20133_);
  nand _53101_ (_20135_, _20134_, _26487_);
  nor _53102_ (_10010_, _20135_, _20132_);
  nand _53103_ (_20136_, _19094_, _24789_);
  nand _53104_ (_20137_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  nand _53105_ (_28332_, _20137_, _20136_);
  nand _53106_ (_20138_, _03958_, _24789_);
  nand _53107_ (_20139_, _03960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  nand _53108_ (_28239_, _20139_, _20138_);
  nand _53109_ (_20140_, _19119_, _25099_);
  nand _53110_ (_20141_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  nand _53111_ (_28331_, _20141_, _20140_);
  nand _53112_ (_20142_, _18519_, _28096_);
  nand _53113_ (_20143_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  nand _53114_ (_10018_, _20143_, _20142_);
  nand _53115_ (_20144_, _00991_, _25203_);
  nand _53116_ (_20145_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  nand _53117_ (_10020_, _20145_, _20144_);
  nand _53118_ (_20146_, _18307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _53119_ (_20147_, _07948_, _25625_);
  nand _53120_ (_20148_, _18580_, _18567_);
  nand _53121_ (_20149_, _20148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _53122_ (_20150_, _18578_, _07946_);
  nor _53123_ (_20151_, _20150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _53124_ (_20152_, _18313_, _07984_);
  nor _53125_ (_20153_, _20152_, _18566_);
  nor _53126_ (_20154_, _20153_, _20151_);
  nand _53127_ (_20155_, _20154_, _20149_);
  nor _53128_ (_20156_, _20155_, _07948_);
  nor _53129_ (_20157_, _20156_, _18329_);
  nand _53130_ (_20158_, _20157_, _20147_);
  nand _53131_ (_10027_, _20158_, _20146_);
  nand _53132_ (_20159_, _11827_, _28096_);
  nand _53133_ (_20160_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  nand _53134_ (_10039_, _20160_, _20159_);
  nor _53135_ (_20161_, _05481_, _02726_);
  not _53136_ (_20162_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand _53137_ (_20163_, _20009_, _20162_);
  nand _53138_ (_20164_, _20163_, _05481_);
  nor _53139_ (_20165_, _20009_, _02685_);
  nor _53140_ (_20166_, _20165_, _20164_);
  nor _53141_ (_20167_, _20166_, _20161_);
  nor _53142_ (_10048_, _20167_, rst);
  nand _53143_ (_20168_, _18946_, _25039_);
  nand _53144_ (_20169_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  nand _53145_ (_10052_, _20169_, _20168_);
  nor _53146_ (_20170_, _00631_, _24978_);
  nand _53147_ (_20171_, _20170_, _24789_);
  not _53148_ (_20172_, _20170_);
  nand _53149_ (_20173_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  nand _53150_ (_10056_, _20173_, _20171_);
  nand _53151_ (_20175_, _03822_, _24927_);
  nand _53152_ (_20176_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  nand _53153_ (_10061_, _20176_, _20175_);
  nand _53154_ (_20177_, _07908_, _25150_);
  nand _53155_ (_20178_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nand _53156_ (_10065_, _20178_, _20177_);
  nor _53157_ (_20179_, _05481_, _02652_);
  not _53158_ (_20180_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nand _53159_ (_20181_, _20009_, _20180_);
  nand _53160_ (_20182_, _20181_, _05481_);
  nor _53161_ (_20183_, _20009_, _02620_);
  nor _53162_ (_20184_, _20183_, _20182_);
  nor _53163_ (_20185_, _20184_, _20179_);
  nor _53164_ (_10072_, _20185_, rst);
  nand _53165_ (_20186_, _18125_, _24830_);
  nand _53166_ (_20187_, _18127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nand _53167_ (_28268_, _20187_, _20186_);
  nand _53168_ (_20188_, _03858_, _24830_);
  nand _53169_ (_20189_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  nand _53170_ (_10079_, _20189_, _20188_);
  nand _53171_ (_20190_, _19024_, _24830_);
  nand _53172_ (_20191_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nand _53173_ (_10080_, _20191_, _20190_);
  nand _53174_ (_20192_, _18713_, _25039_);
  nand _53175_ (_20193_, _18715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  nand _53176_ (_10083_, _20193_, _20192_);
  nand _53177_ (_20194_, _03840_, _25099_);
  nand _53178_ (_20195_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nand _53179_ (_10086_, _20195_, _20194_);
  nand _53180_ (_20196_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nand _53181_ (_20197_, _08324_, _25039_);
  nand _53182_ (_10088_, _20197_, _20196_);
  nand _53183_ (_20198_, _04312_, _24789_);
  nand _53184_ (_20199_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  nand _53185_ (_10094_, _20199_, _20198_);
  nor _53186_ (_20200_, _20029_, _02509_);
  not _53187_ (_20201_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand _53188_ (_20202_, _20029_, _20201_);
  nand _53189_ (_20203_, _20202_, _26487_);
  nor _53190_ (_10099_, _20203_, _20200_);
  nor _53191_ (_20204_, _20029_, _02761_);
  not _53192_ (_20205_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand _53193_ (_20206_, _20029_, _20205_);
  nand _53194_ (_20207_, _20206_, _26487_);
  nor _53195_ (_10101_, _20207_, _20204_);
  nor _53196_ (_20208_, _20029_, _02685_);
  not _53197_ (_20209_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand _53198_ (_20210_, _20029_, _20209_);
  nand _53199_ (_20211_, _20210_, _26487_);
  nor _53200_ (_10103_, _20211_, _20208_);
  nor _53201_ (_20212_, _05481_, _02598_);
  not _53202_ (_20213_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand _53203_ (_20214_, _20009_, _20213_);
  nand _53204_ (_20215_, _20214_, _05481_);
  nor _53205_ (_20216_, _20009_, _02096_);
  nor _53206_ (_20217_, _20216_, _20215_);
  nor _53207_ (_20218_, _20217_, _20212_);
  nor _53208_ (_10106_, _20218_, rst);
  nor _53209_ (_20219_, _05481_, _02540_);
  not _53210_ (_20220_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand _53211_ (_20221_, _20009_, _20220_);
  nand _53212_ (_20222_, _20221_, _05481_);
  nor _53213_ (_20223_, _20009_, _02509_);
  nor _53214_ (_20224_, _20223_, _20222_);
  nor _53215_ (_20225_, _20224_, _20219_);
  nor _53216_ (_10109_, _20225_, rst);
  nand _53217_ (_20226_, _11633_, _25150_);
  nand _53218_ (_20227_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nand _53219_ (_10112_, _20227_, _20226_);
  nand _53220_ (_20228_, _18131_, _24789_);
  nand _53221_ (_20229_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  nand _53222_ (_28267_, _20229_, _20228_);
  nand _53223_ (_20230_, _18131_, _25150_);
  nand _53224_ (_20231_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  nand _53225_ (_10116_, _20231_, _20230_);
  nand _53226_ (_20232_, _25099_, _24852_);
  nand _53227_ (_20233_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nand _53228_ (_10118_, _20233_, _20232_);
  nand _53229_ (_20234_, _20170_, _25039_);
  nand _53230_ (_20235_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nand _53231_ (_10128_, _20235_, _20234_);
  nand _53232_ (_20236_, _00150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _53233_ (_20237_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  not _53234_ (_20238_, _00200_);
  nand _53235_ (_20239_, _20238_, _00242_);
  nand _53236_ (_20240_, _20239_, _00201_);
  nand _53237_ (_20241_, _20240_, _00158_);
  not _53238_ (_20242_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand _53239_ (_20243_, _00245_, _00205_);
  nor _53240_ (_20244_, _20243_, _20242_);
  nor _53241_ (_20245_, _20244_, _20241_);
  nor _53242_ (_20246_, _20245_, _20237_);
  nand _53243_ (_20247_, _20246_, _00240_);
  nand _53244_ (_20248_, _20247_, _20236_);
  nor _53245_ (_20249_, _00141_, _25140_);
  nor _53246_ (_20250_, _20249_, _20248_);
  nor _53247_ (_10130_, _20250_, rst);
  nor _53248_ (_20251_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand _53249_ (_20252_, _00199_, _00161_);
  nand _53250_ (_20253_, _20252_, _20238_);
  nand _53251_ (_20254_, _20253_, _00158_);
  not _53252_ (_20255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor _53253_ (_20256_, _20243_, _20255_);
  nor _53254_ (_20257_, _20256_, _20254_);
  nor _53255_ (_20258_, _20257_, _20251_);
  nand _53256_ (_20259_, _20258_, _00240_);
  nand _53257_ (_20260_, _00150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand _53258_ (_20261_, _20260_, _20259_);
  nor _53259_ (_20262_, _00141_, _26096_);
  nor _53260_ (_20264_, _20262_, _20261_);
  nor _53261_ (_10132_, _20264_, rst);
  nand _53262_ (_20265_, _00150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _53263_ (_20266_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand _53264_ (_20267_, _00197_, _00162_);
  nand _53265_ (_20268_, _20267_, _00199_);
  nand _53266_ (_20269_, _20268_, _00158_);
  not _53267_ (_20270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _53268_ (_20271_, _20243_, _20270_);
  nor _53269_ (_20272_, _20271_, _20269_);
  nor _53270_ (_20273_, _20272_, _20266_);
  nand _53271_ (_20274_, _20273_, _00240_);
  nand _53272_ (_20275_, _20274_, _20265_);
  nor _53273_ (_20276_, _00141_, _25029_);
  nor _53274_ (_20277_, _20276_, _20275_);
  nor _53275_ (_10134_, _20277_, rst);
  nand _53276_ (_20278_, _00356_, _25039_);
  nand _53277_ (_20279_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nand _53278_ (_10136_, _20279_, _20278_);
  nand _53279_ (_20280_, _00416_, _24789_);
  nand _53280_ (_20281_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  nand _53281_ (_10139_, _20281_, _20280_);
  nand _53282_ (_20282_, _07670_, _24830_);
  nand _53283_ (_20283_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  nand _53284_ (_10141_, _20283_, _20282_);
  nand _53285_ (_20284_, _20170_, _25203_);
  nand _53286_ (_20285_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nand _53287_ (_10143_, _20285_, _20284_);
  nand _53288_ (_20286_, _01587_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nand _53289_ (_20287_, _20286_, _08000_);
  not _53290_ (_20288_, _20286_);
  nor _53291_ (_20289_, _20288_, _01631_);
  nor _53292_ (_20290_, _20289_, _04226_);
  nand _53293_ (_20291_, _20290_, _20287_);
  nor _53294_ (_20292_, _20288_, _12077_);
  nor _53295_ (_20293_, _20292_, _04208_);
  nor _53296_ (_20294_, _20289_, _01609_);
  nor _53297_ (_20295_, _20294_, _20293_);
  nand _53298_ (_20296_, _20295_, _20291_);
  nor _53299_ (_20297_, _04172_, rst);
  nand _53300_ (_20298_, _20297_, _20296_);
  nor _53301_ (_10145_, _20298_, _01573_);
  not _53302_ (_20299_, _02861_);
  nor _53303_ (_20300_, _05481_, _20299_);
  not _53304_ (_20301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand _53305_ (_20302_, _20009_, _20301_);
  nand _53306_ (_20303_, _20302_, _05481_);
  nor _53307_ (_20304_, _20009_, _02373_);
  nor _53308_ (_20305_, _20304_, _20303_);
  nor _53309_ (_20306_, _20305_, _20300_);
  nor _53310_ (_10146_, _20306_, rst);
  nand _53311_ (_20307_, _08325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  nand _53312_ (_20308_, _08324_, _25203_);
  nand _53313_ (_10151_, _20308_, _20307_);
  nand _53314_ (_20309_, _00632_, _24830_);
  nand _53315_ (_20310_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  nand _53316_ (_10153_, _20310_, _20309_);
  nand _53317_ (_20311_, _00735_, _25150_);
  nand _53318_ (_20312_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  nand _53319_ (_10155_, _20312_, _20311_);
  nand _53320_ (_20313_, _00927_, _25203_);
  nand _53321_ (_20314_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  nand _53322_ (_10159_, _20314_, _20313_);
  nand _53323_ (_20315_, _00927_, _24830_);
  nand _53324_ (_20316_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nand _53325_ (_10164_, _20316_, _20315_);
  nand _53326_ (_20317_, _25203_, _25061_);
  nand _53327_ (_20318_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  nand _53328_ (_28333_, _20318_, _20317_);
  nand _53329_ (_20319_, _00150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor _53330_ (_20320_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _53331_ (_20321_, _00196_, _00193_);
  not _53332_ (_20322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nand _53333_ (_20323_, _00257_, _00205_);
  nor _53334_ (_20324_, _20323_, _20322_);
  nor _53335_ (_20325_, _20324_, _20321_);
  nor _53336_ (_20326_, _20325_, _00170_);
  nand _53337_ (_20327_, _00197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _53338_ (_20328_, _20327_, _00158_);
  nor _53339_ (_20329_, _20328_, _20326_);
  nor _53340_ (_20331_, _20329_, _20320_);
  nand _53341_ (_20332_, _20331_, _00240_);
  nand _53342_ (_20333_, _20332_, _20319_);
  nor _53343_ (_20334_, _00141_, _25195_);
  nor _53344_ (_20335_, _20334_, _20333_);
  nor _53345_ (_10172_, _20335_, rst);
  nand _53346_ (_20336_, _18545_, _25203_);
  nand _53347_ (_20337_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  nand _53348_ (_28265_, _20337_, _20336_);
  nand _53349_ (_20338_, _04624_, _25150_);
  nand _53350_ (_20339_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nand _53351_ (_10194_, _20339_, _20338_);
  nand _53352_ (_20340_, _20170_, _28096_);
  nand _53353_ (_20341_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  nand _53354_ (_10199_, _20341_, _20340_);
  nand _53355_ (_20342_, _04006_, _28096_);
  nand _53356_ (_20343_, _04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nand _53357_ (_10203_, _20343_, _20342_);
  nand _53358_ (_20344_, _04308_, _24927_);
  nand _53359_ (_20345_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  nand _53360_ (_10208_, _20345_, _20344_);
  nand _53361_ (_20346_, _03858_, _24789_);
  nand _53362_ (_20347_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  nand _53363_ (_10210_, _20347_, _20346_);
  nand _53364_ (_20348_, _18545_, _24927_);
  nand _53365_ (_20349_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  nand _53366_ (_10219_, _20349_, _20348_);
  nand _53367_ (_20350_, _03840_, _24789_);
  nand _53368_ (_20351_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  nand _53369_ (_10221_, _20351_, _20350_);
  nand _53370_ (_20352_, _28063_, _25099_);
  nand _53371_ (_20353_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  nand _53372_ (_28314_, _20353_, _20352_);
  nand _53373_ (_20354_, _25150_, _25000_);
  nand _53374_ (_20355_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  nand _53375_ (_28313_, _20355_, _20354_);
  nand _53376_ (_20356_, _04312_, _25203_);
  nand _53377_ (_20357_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  nand _53378_ (_10227_, _20357_, _20356_);
  nand _53379_ (_20358_, _28099_, _28096_);
  nand _53380_ (_20359_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nand _53381_ (_10229_, _20359_, _20358_);
  nand _53382_ (_20360_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _53383_ (_20361_, _20360_);
  nor _53384_ (_20362_, _20361_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _53385_ (_20363_, _24639_, _24591_);
  nand _53386_ (_20364_, _02203_, _24088_);
  nor _53387_ (_20365_, _27447_, _02078_);
  nor _53388_ (_20366_, _20365_, _20360_);
  nand _53389_ (_20367_, _20366_, _20364_);
  nor _53390_ (_20368_, _20367_, _20363_);
  nor _53391_ (_20369_, _20368_, _20362_);
  nor _53392_ (_20370_, _20369_, _26261_);
  nand _53393_ (_20371_, _01666_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _53394_ (_20372_, _20371_, _26261_);
  nor _53395_ (_20373_, _20372_, _07866_);
  nor _53396_ (_20374_, _20373_, _20370_);
  nor _53397_ (_20375_, _20374_, _25729_);
  nand _53398_ (_20376_, _25729_, _25140_);
  nand _53399_ (_20377_, _20376_, _26487_);
  nor _53400_ (_10231_, _20377_, _20375_);
  nor _53401_ (_10236_, _04762_, rst);
  nand _53402_ (_20378_, _00123_, _24830_);
  nand _53403_ (_20379_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nand _53404_ (_10239_, _20379_, _20378_);
  nand _53405_ (_20380_, _00632_, _25039_);
  nand _53406_ (_20381_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  nand _53407_ (_10261_, _20381_, _20380_);
  nand _53408_ (_20382_, _19119_, _28096_);
  nand _53409_ (_20383_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nand _53410_ (_10269_, _20383_, _20382_);
  nand _53411_ (_20384_, _18946_, _24927_);
  nand _53412_ (_20385_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  nand _53413_ (_28327_, _20385_, _20384_);
  nor _53414_ (_20386_, _04175_, _24782_);
  nor _53415_ (_20387_, _07637_, _07998_);
  nor _53416_ (_20388_, _18798_, _04215_);
  nand _53417_ (_20389_, _20388_, _01618_);
  not _53418_ (_20390_, _20388_);
  nand _53419_ (_20391_, _20390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand _53420_ (_20392_, _20391_, _20389_);
  nor _53421_ (_20393_, _20392_, _20387_);
  nor _53422_ (_20394_, _20393_, _01644_);
  nor _53423_ (_20395_, _01642_, _01618_);
  nor _53424_ (_20396_, _20395_, _20394_);
  nand _53425_ (_20397_, _20396_, _04175_);
  nand _53426_ (_20398_, _20397_, _26487_);
  nor _53427_ (_10279_, _20398_, _20386_);
  not _53428_ (_20399_, _25741_);
  nand _53429_ (_20400_, _26261_, _00444_);
  nor _53430_ (_20401_, _20400_, _24716_);
  nand _53431_ (_20402_, _20400_, _25738_);
  nand _53432_ (_20403_, _20402_, _20117_);
  nor _53433_ (_20404_, _20403_, _20401_);
  nor _53434_ (_20405_, _20404_, _20399_);
  nor _53435_ (_10295_, _20405_, rst);
  not _53436_ (_20406_, _04585_);
  nand _53437_ (_20407_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  nand _53438_ (_10301_, _20407_, _20406_);
  nor _53439_ (_20408_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor _53440_ (_20410_, _24647_, _24645_);
  not _53441_ (_20411_, _24592_);
  nand _53442_ (_20412_, _24645_, _20411_);
  nand _53443_ (_20413_, _20412_, _24590_);
  nor _53444_ (_20414_, _20413_, _20410_);
  nand _53445_ (_20415_, _24574_, _24761_);
  nor _53446_ (_20416_, _24574_, _24577_);
  nor _53447_ (_20417_, _20416_, _24089_);
  nand _53448_ (_20418_, _20417_, _20415_);
  nor _53449_ (_20419_, _24353_, _24296_);
  nor _53450_ (_20420_, _24508_, _24439_);
  nand _53451_ (_20421_, _20420_, _20419_);
  nand _53452_ (_20422_, _27533_, _26911_);
  nor _53453_ (_20423_, _20422_, _20421_);
  nand _53454_ (_20424_, _20423_, _24767_);
  nand _53455_ (_20425_, _20424_, _20418_);
  nor _53456_ (_20426_, _20425_, _20414_);
  nand _53457_ (_20427_, _02338_, _27396_);
  not _53458_ (_20428_, _02200_);
  nor _53459_ (_20429_, _02000_, _01952_);
  nand _53460_ (_20430_, _20429_, _02067_);
  nor _53461_ (_20431_, _20430_, _02132_);
  nand _53462_ (_20432_, _20431_, _20428_);
  nor _53463_ (_20433_, _20432_, _02269_);
  nand _53464_ (_20434_, _20433_, _20427_);
  nand _53465_ (_20435_, _20434_, _24770_);
  nand _53466_ (_20436_, _20435_, _20426_);
  nand _53467_ (_20437_, _27417_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor _53468_ (_20438_, _20437_, _20436_);
  nor _53469_ (_20439_, _20438_, _20408_);
  nor _53470_ (_20440_, _20439_, _26261_);
  nand _53471_ (_20441_, _00276_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand _53472_ (_20442_, _20441_, _03603_);
  nor _53473_ (_20443_, _20442_, _26262_);
  nor _53474_ (_20444_, _20443_, _20440_);
  nor _53475_ (_20445_, _20444_, _25729_);
  nand _53476_ (_20446_, _25729_, _25703_);
  nand _53477_ (_20447_, _20446_, _26487_);
  nor _53478_ (_10304_, _20447_, _20445_);
  not _53479_ (_20448_, _25732_);
  nor _53480_ (_20449_, _26262_, _00147_);
  not _53481_ (_20450_, _20449_);
  nor _53482_ (_20451_, _20450_, _24716_);
  nand _53483_ (_20452_, _20450_, _25720_);
  nand _53484_ (_20453_, _20452_, _20117_);
  nor _53485_ (_20454_, _20453_, _20451_);
  nor _53486_ (_20455_, _20454_, _20448_);
  nor _53487_ (_10307_, _20455_, rst);
  nand _53488_ (_20456_, _18545_, _25039_);
  nand _53489_ (_20457_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nand _53490_ (_10310_, _20457_, _20456_);
  nand _53491_ (_20459_, _26261_, _24840_);
  nor _53492_ (_20460_, _20459_, _24716_);
  nand _53493_ (_20461_, _20459_, _04901_);
  nand _53494_ (_20462_, _20461_, _20117_);
  nor _53495_ (_20463_, _20462_, _20460_);
  nor _53496_ (_20464_, _20117_, _25088_);
  nor _53497_ (_20465_, _20464_, _20463_);
  nor _53498_ (_10321_, _20465_, rst);
  nand _53499_ (_20466_, _26261_, _03356_);
  nor _53500_ (_20467_, _20466_, _24716_);
  not _53501_ (_20468_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand _53502_ (_20469_, _20466_, _20468_);
  nand _53503_ (_20470_, _20469_, _20117_);
  nor _53504_ (_20471_, _20470_, _20467_);
  nor _53505_ (_20472_, _20117_, _26096_);
  nor _53506_ (_20473_, _20472_, _20471_);
  nor _53507_ (_10323_, _20473_, rst);
  nand _53508_ (_20474_, _07670_, _28096_);
  nand _53509_ (_20475_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nand _53510_ (_10340_, _20475_, _20474_);
  nand _53511_ (_20476_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nand _53512_ (_20477_, _04601_, _25150_);
  nand _53513_ (_10342_, _20477_, _20476_);
  nor _53514_ (_20478_, _25051_, _24795_);
  not _53515_ (_20479_, _20478_);
  nand _53516_ (_20480_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nand _53517_ (_20481_, _20478_, _25203_);
  nand _53518_ (_10344_, _20481_, _20480_);
  nand _53519_ (_20482_, _00150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _53520_ (_20483_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  not _53521_ (_20484_, _00257_);
  not _53522_ (_20485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _53523_ (_20486_, _00204_, _20485_);
  nand _53524_ (_20487_, _20486_, _00169_);
  nor _53525_ (_20488_, _20487_, _20484_);
  nand _53526_ (_20489_, _00189_, _00169_);
  nor _53527_ (_20490_, _20489_, _00190_);
  not _53528_ (_20491_, _20490_);
  nand _53529_ (_20492_, _20489_, _00190_);
  nand _53530_ (_20493_, _20492_, _20491_);
  nand _53531_ (_20494_, _20493_, _00158_);
  nor _53532_ (_20495_, _20494_, _20488_);
  nor _53533_ (_20496_, _20495_, _20483_);
  nand _53534_ (_20497_, _20496_, _00240_);
  nand _53535_ (_20498_, _20497_, _20482_);
  nor _53536_ (_20499_, _00141_, _25088_);
  nor _53537_ (_20500_, _20499_, _20498_);
  nor _53538_ (_10347_, _20500_, rst);
  nand _53539_ (_20501_, _25061_, _25039_);
  nand _53540_ (_20502_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nand _53541_ (_10349_, _20502_, _20501_);
  nand _53542_ (_20503_, _18946_, _25150_);
  nand _53543_ (_20504_, _18948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nand _53544_ (_28328_, _20504_, _20503_);
  nor _53545_ (_20505_, _01000_, _25057_);
  nand _53546_ (_20506_, _20505_, _25203_);
  not _53547_ (_20507_, _20505_);
  nand _53548_ (_20508_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  nand _53549_ (_10358_, _20508_, _20506_);
  nand _53550_ (_20509_, _20505_, _24830_);
  nand _53551_ (_20510_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nand _53552_ (_10361_, _20510_, _20509_);
  nor _53553_ (_20511_, _01000_, _28080_);
  nand _53554_ (_20512_, _20511_, _24789_);
  not _53555_ (_20513_, _20511_);
  nand _53556_ (_20514_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  nand _53557_ (_10364_, _20514_, _20512_);
  nand _53558_ (_20515_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  nand _53559_ (_20516_, _20478_, _28096_);
  nand _53560_ (_10367_, _20516_, _20515_);
  nand _53561_ (_20517_, _20511_, _25203_);
  nand _53562_ (_20518_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nand _53563_ (_10371_, _20518_, _20517_);
  nand _53564_ (_20519_, _20511_, _25099_);
  nand _53565_ (_20520_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  nand _53566_ (_10373_, _20520_, _20519_);
  nor _53567_ (_20521_, _01000_, _28073_);
  nand _53568_ (_20522_, _20521_, _25039_);
  not _53569_ (_20523_, _20521_);
  nand _53570_ (_20524_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  nand _53571_ (_28343_, _20524_, _20522_);
  nand _53572_ (_20525_, _00150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _53573_ (_20526_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nand _53574_ (_20527_, _20491_, _00191_);
  nand _53575_ (_20528_, _20490_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _53576_ (_20529_, _20528_, _20527_);
  nand _53577_ (_20530_, _20529_, _00158_);
  not _53578_ (_20531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _53579_ (_20532_, _20243_, _20531_);
  nor _53580_ (_20533_, _20532_, _20530_);
  nor _53581_ (_20534_, _20533_, _20526_);
  nand _53582_ (_20535_, _20534_, _00240_);
  nand _53583_ (_20536_, _20535_, _20525_);
  nor _53584_ (_20537_, _00141_, _25703_);
  nor _53585_ (_20538_, _20537_, _20536_);
  nor _53586_ (_10379_, _20538_, rst);
  nand _53587_ (_20539_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  nand _53588_ (_20540_, _20478_, _25099_);
  nand _53589_ (_28303_, _20540_, _20539_);
  nand _53590_ (_20541_, _20521_, _28096_);
  nand _53591_ (_20542_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  nand _53592_ (_10385_, _20542_, _20541_);
  nor _53593_ (_20543_, _01000_, _00122_);
  nand _53594_ (_20544_, _20543_, _25039_);
  not _53595_ (_20545_, _20543_);
  nand _53596_ (_20546_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  nand _53597_ (_28342_, _20546_, _20544_);
  nand _53598_ (_20547_, _20543_, _28096_);
  nand _53599_ (_20548_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nand _53600_ (_10393_, _20548_, _20547_);
  nand _53601_ (_20549_, _18131_, _24830_);
  nand _53602_ (_20550_, _18133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  nand _53603_ (_10399_, _20550_, _20549_);
  nand _53604_ (_20551_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nand _53605_ (_20552_, _20478_, _24830_);
  nand _53606_ (_10401_, _20552_, _20551_);
  nand _53607_ (_20553_, _18545_, _24789_);
  nand _53608_ (_20554_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  nand _53609_ (_10403_, _20554_, _20553_);
  nor _53610_ (_20555_, _01000_, _25047_);
  nand _53611_ (_20556_, _20555_, _24927_);
  not _53612_ (_20557_, _20555_);
  nand _53613_ (_20558_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  nand _53614_ (_10405_, _20558_, _20556_);
  nand _53615_ (_20559_, _20555_, _25203_);
  nand _53616_ (_20560_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  nand _53617_ (_10407_, _20560_, _20559_);
  nand _53618_ (_20561_, _20555_, _24830_);
  nand _53619_ (_20562_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nand _53620_ (_10413_, _20562_, _20561_);
  nor _53621_ (_10419_, _04855_, rst);
  nor _53622_ (_20563_, _01000_, _00415_);
  nand _53623_ (_20564_, _20563_, _25150_);
  not _53624_ (_20565_, _20563_);
  nand _53625_ (_20566_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  nand _53626_ (_28340_, _20566_, _20564_);
  nor _53627_ (_10463_, _04753_, rst);
  nand _53628_ (_20567_, _07670_, _25203_);
  nand _53629_ (_20568_, _07674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  nand _53630_ (_10484_, _20568_, _20567_);
  not _53631_ (_20569_, _00315_);
  nand _53632_ (_20570_, _20569_, _00183_);
  nand _53633_ (_20571_, _00315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _53634_ (_20572_, _20571_, _20570_);
  nor _53635_ (_20573_, _20243_, _05946_);
  nor _53636_ (_20574_, _20573_, _00157_);
  nand _53637_ (_20575_, _20574_, _20572_);
  nand _53638_ (_20576_, _00157_, _05946_);
  nand _53639_ (_20577_, _20576_, _20575_);
  nor _53640_ (_20578_, _20577_, _00241_);
  nand _53641_ (_20579_, _00150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _53642_ (_20580_, _00140_, _24821_);
  nand _53643_ (_20581_, _20580_, _20579_);
  nor _53644_ (_20582_, _20581_, _20578_);
  nor _53645_ (_10488_, _20582_, rst);
  nor _53646_ (_10496_, _04808_, rst);
  nand _53647_ (_20583_, _20563_, _28096_);
  nand _53648_ (_20584_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  nand _53649_ (_10513_, _20584_, _20583_);
  nand _53650_ (_20585_, _12089_, _25099_);
  nand _53651_ (_20586_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  nand _53652_ (_10521_, _20586_, _20585_);
  nor _53653_ (_10523_, _04828_, rst);
  nor _53654_ (_10525_, _04811_, rst);
  nor _53655_ (_20587_, _01000_, _24882_);
  nand _53656_ (_20588_, _20587_, _25150_);
  not _53657_ (_20589_, _20587_);
  nand _53658_ (_20590_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  nand _53659_ (_10536_, _20590_, _20588_);
  nor _53660_ (_20591_, _01000_, _00629_);
  nand _53661_ (_20592_, _20591_, _25150_);
  not _53662_ (_20593_, _20591_);
  nand _53663_ (_20594_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  nand _53664_ (_10556_, _20594_, _20592_);
  nand _53665_ (_20595_, _20591_, _25039_);
  nand _53666_ (_20596_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  nand _53667_ (_10562_, _20596_, _20595_);
  nand _53668_ (_20597_, _04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  nand _53669_ (_20598_, _04601_, _24927_);
  nand _53670_ (_28296_, _20598_, _20597_);
  nand _53671_ (_20599_, _20170_, _25150_);
  nand _53672_ (_20600_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  nand _53673_ (_10587_, _20600_, _20599_);
  nand _53674_ (_20601_, _20591_, _24830_);
  nand _53675_ (_20602_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nand _53676_ (_10601_, _20602_, _20601_);
  nand _53677_ (_20603_, _01108_, _24789_);
  nand _53678_ (_20604_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  nand _53679_ (_10610_, _20604_, _20603_);
  nand _53680_ (_20606_, _01153_, _24830_);
  nand _53681_ (_20607_, _01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  nand _53682_ (_10614_, _20607_, _20606_);
  nand _53683_ (_20608_, _18519_, _25203_);
  nand _53684_ (_20609_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  nand _53685_ (_10618_, _20609_, _20608_);
  nor _53686_ (_20610_, _01000_, _00954_);
  nand _53687_ (_20611_, _20610_, _25039_);
  not _53688_ (_20612_, _20610_);
  nand _53689_ (_20613_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  nand _53690_ (_10634_, _20613_, _20611_);
  nand _53691_ (_20614_, _08806_, _24927_);
  nand _53692_ (_20615_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  nand _53693_ (_10637_, _20615_, _20614_);
  nor _53694_ (_10640_, _04698_, rst);
  nand _53695_ (_20616_, _18519_, _24927_);
  nand _53696_ (_20617_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  nand _53697_ (_10647_, _20617_, _20616_);
  nor _53698_ (_20618_, _01000_, _00393_);
  nand _53699_ (_20619_, _20618_, _24927_);
  not _53700_ (_20620_, _20618_);
  nand _53701_ (_20621_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  nand _53702_ (_28338_, _20621_, _20619_);
  nand _53703_ (_20622_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  nand _53704_ (_20623_, _20478_, _24789_);
  nand _53705_ (_28305_, _20623_, _20622_);
  nor _53706_ (_10656_, _04682_, rst);
  nand _53707_ (_20624_, _01116_, _25099_);
  nand _53708_ (_20625_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nand _53709_ (_10660_, _20625_, _20624_);
  nand _53710_ (_20626_, _01182_, _25150_);
  nand _53711_ (_20627_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  nand _53712_ (_10670_, _20627_, _20626_);
  nor _53713_ (_20628_, _00302_, _25140_);
  nor _53714_ (_20629_, _00308_, _00170_);
  nor _53715_ (_20630_, _20629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _53716_ (_20631_, _20630_, _00311_);
  not _53717_ (_20632_, _20323_);
  nor _53718_ (_20633_, _00170_, _13092_);
  nand _53719_ (_20634_, _20633_, _20632_);
  nand _53720_ (_20635_, _20634_, _00158_);
  nor _53721_ (_20636_, _20635_, _20631_);
  nor _53722_ (_20637_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _53723_ (_20638_, _20637_, _20636_);
  nand _53724_ (_20639_, _20638_, _00240_);
  nand _53725_ (_20640_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _53726_ (_20641_, _20640_, _20639_);
  nor _53727_ (_20642_, _20641_, _20628_);
  nor _53728_ (_10676_, _20642_, rst);
  nand _53729_ (_20643_, _20511_, _24927_);
  nand _53730_ (_20644_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  nand _53731_ (_10678_, _20644_, _20643_);
  nand _53732_ (_20645_, _20521_, _25150_);
  nand _53733_ (_20646_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nand _53734_ (_10685_, _20646_, _20645_);
  nand _53735_ (_20647_, _20543_, _25150_);
  nand _53736_ (_20648_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  nand _53737_ (_10691_, _20648_, _20647_);
  nand _53738_ (_20649_, _04111_, _28096_);
  nand _53739_ (_20650_, _04113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand _53740_ (_28376_, _20650_, _20649_);
  nand _53741_ (_20651_, _20555_, _24789_);
  nand _53742_ (_20652_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  nand _53743_ (_10695_, _20652_, _20651_);
  nor _53744_ (_20653_, _00302_, _25029_);
  nand _53745_ (_20654_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _53746_ (_20655_, _00307_, _00169_);
  nor _53747_ (_20656_, _00306_, _00170_);
  not _53748_ (_20657_, _20656_);
  nand _53749_ (_20658_, _20657_, _00172_);
  nand _53750_ (_20659_, _20658_, _20655_);
  nand _53751_ (_20660_, _20659_, _00158_);
  nand _53752_ (_20661_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor _53753_ (_20662_, _20661_, _20323_);
  nor _53754_ (_20663_, _20662_, _20660_);
  nor _53755_ (_20664_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor _53756_ (_20665_, _20664_, _20663_);
  nand _53757_ (_20666_, _20665_, _00240_);
  nand _53758_ (_20667_, _20666_, _20654_);
  nor _53759_ (_20668_, _20667_, _20653_);
  nor _53760_ (_10701_, _20668_, rst);
  nor _53761_ (_20669_, _00302_, _26096_);
  nor _53762_ (_20670_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  not _53763_ (_20671_, _20629_);
  nand _53764_ (_20672_, _20655_, _00173_);
  nand _53765_ (_20673_, _20672_, _20671_);
  nand _53766_ (_20674_, _20673_, _00158_);
  not _53767_ (_20675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _53768_ (_20676_, _20243_, _20675_);
  nor _53769_ (_20677_, _20676_, _20674_);
  nor _53770_ (_20678_, _20677_, _20670_);
  nand _53771_ (_20679_, _20678_, _00240_);
  nand _53772_ (_20680_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand _53773_ (_20681_, _20680_, _20679_);
  nor _53774_ (_20682_, _20681_, _20669_);
  nor _53775_ (_10705_, _20682_, rst);
  nand _53776_ (_20683_, _18286_, _25039_);
  nand _53777_ (_20684_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  nand _53778_ (_10709_, _20684_, _20683_);
  nor _53779_ (_20685_, _00302_, _25195_);
  nand _53780_ (_20686_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _53781_ (_20687_, _00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand _53782_ (_20688_, _12437_, _00181_);
  nand _53783_ (_20689_, _20688_, _20657_);
  nand _53784_ (_20690_, _20689_, _00158_);
  nand _53785_ (_20691_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor _53786_ (_20692_, _20691_, _20323_);
  nor _53787_ (_20693_, _20692_, _20690_);
  nor _53788_ (_20694_, _20693_, _20687_);
  nand _53789_ (_20695_, _20694_, _00240_);
  nand _53790_ (_20696_, _20695_, _20686_);
  nor _53791_ (_20697_, _20696_, _20685_);
  nor _53792_ (_10713_, _20697_, rst);
  nand _53793_ (_20698_, _20618_, _25099_);
  nand _53794_ (_20699_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  nand _53795_ (_10724_, _20699_, _20698_);
  nand _53796_ (_20700_, _20587_, _25203_);
  nand _53797_ (_20701_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  nand _53798_ (_10727_, _20701_, _20700_);
  nand _53799_ (_20702_, _07908_, _25039_);
  nand _53800_ (_20703_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nand _53801_ (_10730_, _20703_, _20702_);
  nand _53802_ (_20704_, _01182_, _24927_);
  nand _53803_ (_20705_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  nand _53804_ (_10732_, _20705_, _20704_);
  nand _53805_ (_20706_, _08653_, _25203_);
  nand _53806_ (_20707_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  nand _53807_ (_28293_, _20707_, _20706_);
  nand _53808_ (_20708_, _20610_, _25150_);
  nand _53809_ (_20709_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  nand _53810_ (_10739_, _20709_, _20708_);
  nand _53811_ (_20710_, _12089_, _24830_);
  nand _53812_ (_20711_, _12092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  nand _53813_ (_10744_, _20711_, _20710_);
  nand _53814_ (_20712_, _20505_, _25039_);
  nand _53815_ (_20713_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  nand _53816_ (_28344_, _20713_, _20712_);
  nand _53817_ (_20714_, _20587_, _24830_);
  nand _53818_ (_20715_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  nand _53819_ (_10757_, _20715_, _20714_);
  nand _53820_ (_20716_, _20610_, _24830_);
  nand _53821_ (_20717_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  nand _53822_ (_10766_, _20717_, _20716_);
  nand _53823_ (_20718_, _20543_, _24789_);
  nand _53824_ (_20719_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  nand _53825_ (_10773_, _20719_, _20718_);
  nand _53826_ (_20720_, _18286_, _25150_);
  nand _53827_ (_20721_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nand _53828_ (_10779_, _20721_, _20720_);
  nor _53829_ (_20722_, _00122_, _24984_);
  nand _53830_ (_20723_, _20722_, _25039_);
  not _53831_ (_20724_, _20722_);
  nand _53832_ (_20725_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  nand _53833_ (_10792_, _20725_, _20723_);
  nor _53834_ (_20726_, _25047_, _24984_);
  nand _53835_ (_20727_, _20726_, _25150_);
  not _53836_ (_20728_, _20726_);
  nand _53837_ (_20729_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  nand _53838_ (_10799_, _20729_, _20727_);
  nand _53839_ (_20730_, _18286_, _24927_);
  nand _53840_ (_20731_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  nand _53841_ (_10802_, _20731_, _20730_);
  nor _53842_ (_20732_, _03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _53843_ (_28236_, _20732_, _04340_);
  nand _53844_ (_20733_, _20726_, _25099_);
  nand _53845_ (_20734_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nand _53846_ (_10807_, _20734_, _20733_);
  nor _53847_ (_20735_, _00415_, _24984_);
  nand _53848_ (_20736_, _20735_, _24789_);
  not _53849_ (_20737_, _20735_);
  nand _53850_ (_20738_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  nand _53851_ (_10810_, _20738_, _20736_);
  nand _53852_ (_20739_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  nand _53853_ (_20740_, _20478_, _25150_);
  nand _53854_ (_28304_, _20740_, _20739_);
  nand _53855_ (_20741_, _28081_, _24789_);
  nand _53856_ (_20742_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  nand _53857_ (_10823_, _20742_, _20741_);
  nand _53858_ (_20743_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  nand _53859_ (_20744_, _20478_, _24927_);
  nand _53860_ (_10825_, _20744_, _20743_);
  nor _53861_ (_20745_, _00954_, _24984_);
  nand _53862_ (_20746_, _20745_, _25150_);
  not _53863_ (_20747_, _20745_);
  nand _53864_ (_20748_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  nand _53865_ (_10829_, _20748_, _20746_);
  nand _53866_ (_20749_, _20745_, _25203_);
  nand _53867_ (_20750_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nand _53868_ (_10832_, _20750_, _20749_);
  nor _53869_ (_20751_, _00393_, _24984_);
  nand _53870_ (_20752_, _20751_, _25039_);
  not _53871_ (_20753_, _20751_);
  nand _53872_ (_20754_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nand _53873_ (_10842_, _20754_, _20752_);
  nand _53874_ (_20755_, _25150_, _24985_);
  nand _53875_ (_20756_, _24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nand _53876_ (_10845_, _20756_, _20755_);
  nor _53877_ (_20757_, _24984_, _24882_);
  nand _53878_ (_20758_, _20757_, _24927_);
  not _53879_ (_20759_, _20757_);
  nand _53880_ (_20760_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  nand _53881_ (_10854_, _20760_, _20758_);
  nand _53882_ (_20761_, _20757_, _24830_);
  nand _53883_ (_20762_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  nand _53884_ (_10861_, _20762_, _20761_);
  nor _53885_ (_20763_, _00629_, _24984_);
  nand _53886_ (_20764_, _20763_, _25150_);
  not _53887_ (_20765_, _20763_);
  nand _53888_ (_20766_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  nand _53889_ (_10869_, _20766_, _20764_);
  nor _53890_ (_20767_, _01913_, _00227_);
  nand _53891_ (_20768_, _20767_, _24717_);
  nor _53892_ (_20769_, _20767_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor _53893_ (_20770_, _20769_, _26245_);
  nand _53894_ (_20771_, _20770_, _20768_);
  nand _53895_ (_20772_, _01919_, _25625_);
  nor _53896_ (_20773_, _01919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor _53897_ (_20774_, _20773_, _25631_);
  nand _53898_ (_20775_, _20774_, _20772_);
  nand _53899_ (_20776_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nand _53900_ (_20777_, _20776_, _20775_);
  nor _53901_ (_20778_, _20777_, rst);
  nand _53902_ (_10878_, _20778_, _20771_);
  nand _53903_ (_20779_, _20763_, _25099_);
  nand _53904_ (_20780_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  nand _53905_ (_10885_, _20780_, _20779_);
  nand _53906_ (_20781_, _17060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _53907_ (_20782_, _07987_, _18324_);
  nand _53908_ (_20783_, _20782_, _07983_);
  nand _53909_ (_20784_, _20783_, _20781_);
  nor _53910_ (_20785_, _17050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _53911_ (_20786_, _20785_, _17052_);
  nand _53912_ (_20787_, _20786_, _17059_);
  nand _53913_ (_20788_, _20787_, _07942_);
  nor _53914_ (_20789_, _20788_, _20784_);
  nand _53915_ (_20790_, _07941_, _25088_);
  nand _53916_ (_20791_, _20790_, _26487_);
  nor _53917_ (_10891_, _20791_, _20789_);
  nor _53918_ (_20792_, _01000_, _24795_);
  nand _53919_ (_20793_, _20792_, _25150_);
  not _53920_ (_20794_, _20792_);
  nand _53921_ (_20795_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  nand _53922_ (_28355_, _20795_, _20793_);
  nand _53923_ (_20796_, _12096_, _25150_);
  nand _53924_ (_20797_, _12098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  nand _53925_ (_10898_, _20797_, _20796_);
  nand _53926_ (_20798_, _20792_, _24830_);
  nand _53927_ (_20799_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  nand _53928_ (_10900_, _20799_, _20798_);
  nor _53929_ (_20800_, _01000_, _24059_);
  nand _53930_ (_20801_, _20800_, _24927_);
  not _53931_ (_20802_, _20800_);
  nand _53932_ (_20803_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  nand _53933_ (_10904_, _20803_, _20801_);
  nand _53934_ (_20804_, _20800_, _25099_);
  nand _53935_ (_20805_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nand _53936_ (_10908_, _20805_, _20804_);
  nand _53937_ (_20806_, _20479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  nand _53938_ (_20807_, _20478_, _25039_);
  nand _53939_ (_10914_, _20807_, _20806_);
  nor _53940_ (_20808_, _00114_, _24984_);
  nand _53941_ (_20809_, _20808_, _24927_);
  not _53942_ (_20810_, _20808_);
  nand _53943_ (_20811_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  nand _53944_ (_10917_, _20811_, _20809_);
  nand _53945_ (_20812_, _20808_, _25203_);
  nand _53946_ (_20813_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  nand _53947_ (_10919_, _20813_, _20812_);
  nor _53948_ (_20814_, _01000_, _00926_);
  nand _53949_ (_20815_, _20814_, _24789_);
  not _53950_ (_20816_, _20814_);
  nand _53951_ (_20817_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  nand _53952_ (_10921_, _20817_, _20815_);
  nand _53953_ (_20818_, _20722_, _25099_);
  nand _53954_ (_20819_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nand _53955_ (_10924_, _20819_, _20818_);
  nand _53956_ (_20820_, _20726_, _25203_);
  nand _53957_ (_20821_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nand _53958_ (_28365_, _20821_, _20820_);
  nand _53959_ (_20822_, _20735_, _28096_);
  nand _53960_ (_20823_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nand _53961_ (_10930_, _20823_, _20822_);
  nand _53962_ (_20824_, _20745_, _24830_);
  nand _53963_ (_20825_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  nand _53964_ (_10938_, _20825_, _20824_);
  nand _53965_ (_20826_, _20751_, _25099_);
  nand _53966_ (_20827_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nand _53967_ (_10941_, _20827_, _20826_);
  nand _53968_ (_20828_, _20757_, _28096_);
  nand _53969_ (_20829_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  nand _53970_ (_10943_, _20829_, _20828_);
  nand _53971_ (_20830_, _08653_, _24927_);
  nand _53972_ (_20831_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  nand _53973_ (_10945_, _20831_, _20830_);
  nand _53974_ (_20832_, _20763_, _25203_);
  nand _53975_ (_20833_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nand _53976_ (_10947_, _20833_, _20832_);
  nand _53977_ (_20834_, _04251_, _25203_);
  nand _53978_ (_20835_, _04253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nand _53979_ (_10949_, _20835_, _20834_);
  nand _53980_ (_20836_, _28063_, _25203_);
  nand _53981_ (_20837_, _28065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nand _53982_ (_10954_, _20837_, _20836_);
  nor _53983_ (_20838_, _00227_, _03254_);
  nand _53984_ (_20839_, _20838_, _24717_);
  nor _53985_ (_20840_, _20838_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor _53986_ (_20841_, _20840_, _26245_);
  nand _53987_ (_20842_, _20841_, _20839_);
  nand _53988_ (_20843_, _03260_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand _53989_ (_20844_, _03094_, _24782_);
  nand _53990_ (_20845_, _20844_, _20843_);
  nand _53991_ (_20846_, _20845_, _25630_);
  nand _53992_ (_20847_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand _53993_ (_20848_, _20847_, _20846_);
  nor _53994_ (_20849_, _20848_, rst);
  nand _53995_ (_10960_, _20849_, _20842_);
  nand _53996_ (_20850_, _20792_, _28096_);
  nand _53997_ (_20851_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  nand _53998_ (_10963_, _20851_, _20850_);
  nand _53999_ (_20852_, _20800_, _24789_);
  nand _54000_ (_20853_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  nand _54001_ (_28352_, _20853_, _20852_);
  nand _54002_ (_20854_, _20808_, _24789_);
  nand _54003_ (_20855_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  nand _54004_ (_10968_, _20855_, _20854_);
  nand _54005_ (_20856_, _20722_, _24927_);
  nand _54006_ (_20857_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  nand _54007_ (_10972_, _20857_, _20856_);
  nand _54008_ (_20858_, _19068_, _25099_);
  nand _54009_ (_20859_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  nand _54010_ (_10976_, _20859_, _20858_);
  nand _54011_ (_20860_, _20745_, _25039_);
  nand _54012_ (_20861_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  nand _54013_ (_10981_, _20861_, _20860_);
  nand _54014_ (_20862_, _20751_, _24927_);
  nand _54015_ (_20863_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  nand _54016_ (_10982_, _20863_, _20862_);
  nand _54017_ (_20864_, _20763_, _24789_);
  nand _54018_ (_20865_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  nand _54019_ (_10985_, _20865_, _20864_);
  nand _54020_ (_20866_, _20808_, _24830_);
  nand _54021_ (_20867_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nand _54022_ (_10993_, _20867_, _20866_);
  nand _54023_ (_20868_, _18545_, _25099_);
  nand _54024_ (_20869_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  nand _54025_ (_10997_, _20869_, _20868_);
  nand _54026_ (_20870_, _18545_, _24830_);
  nand _54027_ (_20871_, _18547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nand _54028_ (_10999_, _20871_, _20870_);
  nand _54029_ (_20872_, _20757_, _25150_);
  nand _54030_ (_20874_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nand _54031_ (_11001_, _20874_, _20872_);
  nand _54032_ (_20875_, _20792_, _25203_);
  nand _54033_ (_20876_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  nand _54034_ (_28353_, _20876_, _20875_);
  nand _54035_ (_20877_, _18173_, _25039_);
  nand _54036_ (_20878_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nand _54037_ (_11005_, _20878_, _20877_);
  nand _54038_ (_20879_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nand _54039_ (_20880_, _08329_, _28096_);
  nand _54040_ (_28302_, _20880_, _20879_);
  nand _54041_ (_20881_, _20618_, _24789_);
  nand _54042_ (_20882_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  nand _54043_ (_28339_, _20882_, _20881_);
  nand _54044_ (_20883_, _00927_, _25150_);
  nand _54045_ (_20884_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  nand _54046_ (_11013_, _20884_, _20883_);
  nand _54047_ (_20885_, _07941_, _24820_);
  nand _54048_ (_20886_, _20885_, _26487_);
  nor _54049_ (_20887_, _17059_, _17049_);
  nand _54050_ (_20888_, _07960_, _17049_);
  nor _54051_ (_20889_, _17058_, _17050_);
  nand _54052_ (_20890_, _20889_, _20888_);
  not _54053_ (_20891_, _07945_);
  nor _54054_ (_20892_, _18318_, _20891_);
  nand _54055_ (_20893_, _20892_, _18311_);
  nand _54056_ (_20894_, _20893_, _20890_);
  nand _54057_ (_20895_, _20894_, _07983_);
  nand _54058_ (_20896_, _20895_, _18306_);
  nor _54059_ (_20897_, _20896_, _20887_);
  nor _54060_ (_11019_, _20897_, _20886_);
  nand _54061_ (_20899_, _20814_, _24927_);
  nand _54062_ (_20900_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  nand _54063_ (_11022_, _20900_, _20899_);
  nand _54064_ (_20901_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nand _54065_ (_20902_, _08329_, _25099_);
  nand _54066_ (_11024_, _20902_, _20901_);
  nand _54067_ (_20903_, _20618_, _25039_);
  nand _54068_ (_20904_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  nand _54069_ (_11026_, _20904_, _20903_);
  nand _54070_ (_20905_, _25152_, _25150_);
  nand _54071_ (_20906_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  nand _54072_ (_11028_, _20906_, _20905_);
  nand _54073_ (_20907_, _20618_, _25150_);
  nand _54074_ (_20908_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nand _54075_ (_11030_, _20908_, _20907_);
  nand _54076_ (_20909_, _20814_, _25150_);
  nand _54077_ (_20910_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nand _54078_ (_11032_, _20910_, _20909_);
  nand _54079_ (_20911_, _18537_, _24927_);
  nand _54080_ (_20912_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nand _54081_ (_11034_, _20912_, _20911_);
  nand _54082_ (_20913_, _00927_, _25099_);
  nand _54083_ (_20914_, _00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nand _54084_ (_11036_, _20914_, _20913_);
  nand _54085_ (_20915_, _20808_, _25099_);
  nand _54086_ (_20916_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  nand _54087_ (_28359_, _20916_, _20915_);
  nand _54088_ (_20917_, _20610_, _25099_);
  nand _54089_ (_20918_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nand _54090_ (_11039_, _20918_, _20917_);
  nand _54091_ (_20919_, _00735_, _28096_);
  nand _54092_ (_20920_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  nand _54093_ (_11041_, _20920_, _20919_);
  nand _54094_ (_20921_, _00735_, _24830_);
  nand _54095_ (_20922_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  nand _54096_ (_11043_, _20922_, _20921_);
  nand _54097_ (_20923_, _18173_, _25203_);
  nand _54098_ (_20924_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  nand _54099_ (_11045_, _20924_, _20923_);
  nand _54100_ (_20925_, _20610_, _28096_);
  nand _54101_ (_20926_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  nand _54102_ (_11047_, _20926_, _20925_);
  nand _54103_ (_20927_, _20808_, _28096_);
  nand _54104_ (_20928_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nand _54105_ (_11052_, _20928_, _20927_);
  nand _54106_ (_20929_, _00735_, _25203_);
  nand _54107_ (_20930_, _00737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nand _54108_ (_11053_, _20930_, _20929_);
  nand _54109_ (_20931_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  nand _54110_ (_20932_, _25150_, _24796_);
  nand _54111_ (_11056_, _20932_, _20931_);
  nand _54112_ (_20933_, _20808_, _25039_);
  nand _54113_ (_20934_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nand _54114_ (_28360_, _20934_, _20933_);
  nor _54115_ (_20935_, _01542_, _00227_);
  nand _54116_ (_20936_, _20935_, _24717_);
  nor _54117_ (_20937_, _20935_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor _54118_ (_20938_, _20937_, _26245_);
  nand _54119_ (_20939_, _20938_, _20936_);
  nand _54120_ (_20940_, _01552_, _25625_);
  nor _54121_ (_20941_, _01552_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor _54122_ (_20942_, _20941_, _25631_);
  nand _54123_ (_20943_, _20942_, _20940_);
  nand _54124_ (_20944_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nand _54125_ (_20945_, _20944_, _20943_);
  nor _54126_ (_20946_, _20945_, rst);
  nand _54127_ (_11060_, _20946_, _20939_);
  nand _54128_ (_20947_, _18537_, _25150_);
  nand _54129_ (_20948_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  nand _54130_ (_28263_, _20948_, _20947_);
  nand _54131_ (_20949_, _20610_, _25203_);
  nand _54132_ (_20950_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  nand _54133_ (_11066_, _20950_, _20949_);
  nor _54134_ (_20951_, _00269_, _25139_);
  nor _54135_ (_20952_, _00280_, _20242_);
  nor _54136_ (_20953_, _00282_, _00242_);
  nor _54137_ (_20954_, _20953_, _20952_);
  nand _54138_ (_20955_, _20954_, _00269_);
  nand _54139_ (_20956_, _20955_, _26487_);
  nor _54140_ (_11068_, _20956_, _20951_);
  nand _54141_ (_20957_, _20808_, _25150_);
  nand _54142_ (_20958_, _20810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  nand _54143_ (_11070_, _20958_, _20957_);
  nand _54144_ (_20959_, _20610_, _24927_);
  nand _54145_ (_20960_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  nand _54146_ (_11072_, _20960_, _20959_);
  nand _54147_ (_20961_, _00632_, _25203_);
  nand _54148_ (_20962_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nand _54149_ (_11074_, _20962_, _20961_);
  nand _54150_ (_20963_, _00632_, _28096_);
  nand _54151_ (_20964_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nand _54152_ (_11077_, _20964_, _20963_);
  nand _54153_ (_20965_, _01108_, _24927_);
  nand _54154_ (_20966_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nand _54155_ (_11080_, _20966_, _20965_);
  nand _54156_ (_20967_, _00416_, _25203_);
  nand _54157_ (_20968_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nand _54158_ (_11082_, _20968_, _20967_);
  nor _54159_ (_20969_, _01714_, _00227_);
  nand _54160_ (_20970_, _20969_, _24717_);
  nor _54161_ (_20971_, _20969_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor _54162_ (_20972_, _20971_, _26245_);
  nand _54163_ (_20973_, _20972_, _20970_);
  nand _54164_ (_20974_, _01720_, _25625_);
  nor _54165_ (_20975_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor _54166_ (_20976_, _20975_, _25631_);
  nand _54167_ (_20977_, _20976_, _20974_);
  nand _54168_ (_20978_, _26243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nand _54169_ (_20979_, _20978_, _20977_);
  nor _54170_ (_20980_, _20979_, rst);
  nand _54171_ (_11084_, _20980_, _20973_);
  nand _54172_ (_20981_, _01001_, _24789_);
  nand _54173_ (_20982_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  nand _54174_ (_28349_, _20982_, _20981_);
  nand _54175_ (_20983_, _00416_, _25099_);
  nand _54176_ (_20984_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  nand _54177_ (_11090_, _20984_, _20983_);
  nand _54178_ (_20985_, _20800_, _24830_);
  nand _54179_ (_20986_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nand _54180_ (_28350_, _20986_, _20985_);
  nand _54181_ (_20987_, _01108_, _25150_);
  nand _54182_ (_20988_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  nand _54183_ (_11095_, _20988_, _20987_);
  nand _54184_ (_20989_, _00416_, _24927_);
  nand _54185_ (_20990_, _00418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  nand _54186_ (_11097_, _20990_, _20989_);
  nand _54187_ (_20991_, _20800_, _28096_);
  nand _54188_ (_20992_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  nand _54189_ (_11099_, _20992_, _20991_);
  nand _54190_ (_20993_, _03540_, _25039_);
  nand _54191_ (_20994_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  nand _54192_ (_11103_, _20994_, _20993_);
  nand _54193_ (_20995_, _19068_, _28096_);
  nand _54194_ (_20996_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  nand _54195_ (_11106_, _20996_, _20995_);
  nand _54196_ (_20997_, _00356_, _25099_);
  nand _54197_ (_20998_, _00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nand _54198_ (_11108_, _20998_, _20997_);
  nand _54199_ (_20999_, _20800_, _25203_);
  nand _54200_ (_21001_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nand _54201_ (_11110_, _21001_, _20999_);
  nand _54202_ (_21002_, _20591_, _25099_);
  nand _54203_ (_21003_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  nand _54204_ (_11112_, _21003_, _21002_);
  nand _54205_ (_21004_, _08387_, _25203_);
  nand _54206_ (_21005_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  nand _54207_ (_11115_, _21005_, _21004_);
  nand _54208_ (_21006_, _03894_, _24830_);
  nand _54209_ (_21007_, _03896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nand _54210_ (_11117_, _21007_, _21006_);
  nand _54211_ (_21008_, _20800_, _25039_);
  nand _54212_ (_21009_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  nand _54213_ (_28351_, _21009_, _21008_);
  nand _54214_ (_21010_, _20591_, _28096_);
  nand _54215_ (_21011_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nand _54216_ (_11120_, _21011_, _21010_);
  nand _54217_ (_21012_, _00123_, _25203_);
  nand _54218_ (_21013_, _00125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nand _54219_ (_11121_, _21013_, _21012_);
  nand _54220_ (_21014_, _20800_, _25150_);
  nand _54221_ (_21015_, _20802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nand _54222_ (_11123_, _21015_, _21014_);
  nand _54223_ (_21016_, _28099_, _25099_);
  nand _54224_ (_21017_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nand _54225_ (_28312_, _21017_, _21016_);
  nand _54226_ (_21018_, _20591_, _25203_);
  nand _54227_ (_21019_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nand _54228_ (_11128_, _21019_, _21018_);
  nand _54229_ (_21020_, _28099_, _24927_);
  nand _54230_ (_21021_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  nand _54231_ (_11133_, _21021_, _21020_);
  nand _54232_ (_21022_, _20591_, _24927_);
  nand _54233_ (_21023_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  nand _54234_ (_11136_, _21023_, _21022_);
  nor _54235_ (_21024_, _00269_, _25028_);
  nor _54236_ (_21025_, _00280_, _20270_);
  nor _54237_ (_21026_, _00282_, _00162_);
  nor _54238_ (_21027_, _21026_, _21025_);
  nand _54239_ (_21028_, _21027_, _00269_);
  nand _54240_ (_21029_, _21028_, _26487_);
  nor _54241_ (_11138_, _21029_, _21024_);
  nand _54242_ (_21030_, _28099_, _25039_);
  nand _54243_ (_21031_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  nand _54244_ (_11140_, _21031_, _21030_);
  nand _54245_ (_21032_, _20792_, _25099_);
  nand _54246_ (_21033_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  nand _54247_ (_11142_, _21033_, _21032_);
  nand _54248_ (_21034_, _20591_, _24789_);
  nand _54249_ (_21035_, _20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  nand _54250_ (_11146_, _21035_, _21034_);
  nand _54251_ (_21037_, _07810_, _24789_);
  nand _54252_ (_21038_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  nand _54253_ (_11149_, _21038_, _21037_);
  nand _54254_ (_21039_, _18537_, _24789_);
  nand _54255_ (_21040_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  nand _54256_ (_11151_, _21040_, _21039_);
  nand _54257_ (_21041_, _20792_, _25039_);
  nand _54258_ (_21042_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nand _54259_ (_28354_, _21042_, _21041_);
  nand _54260_ (_21043_, _20587_, _25099_);
  nand _54261_ (_21044_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nand _54262_ (_11154_, _21044_, _21043_);
  not _54263_ (_21045_, _04598_);
  nand _54264_ (_21046_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nand _54265_ (_11157_, _21046_, _21045_);
  nand _54266_ (_21047_, _03442_, _24830_);
  nand _54267_ (_21048_, _03444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  nand _54268_ (_11159_, _21048_, _21047_);
  nand _54269_ (_21049_, _25099_, _24890_);
  nand _54270_ (_21050_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nand _54271_ (_11161_, _21050_, _21049_);
  nand _54272_ (_21051_, _00991_, _24927_);
  nand _54273_ (_21052_, _00993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  nand _54274_ (_11164_, _21052_, _21051_);
  nand _54275_ (_21053_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  nand _54276_ (_21054_, _08329_, _24927_);
  nand _54277_ (_11169_, _21054_, _21053_);
  nand _54278_ (_21055_, _04312_, _28096_);
  nand _54279_ (_21056_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  nand _54280_ (_11171_, _21056_, _21055_);
  nand _54281_ (_21057_, _20792_, _24927_);
  nand _54282_ (_21058_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  nand _54283_ (_11173_, _21058_, _21057_);
  nand _54284_ (_21059_, _18286_, _25099_);
  nand _54285_ (_21060_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  nand _54286_ (_28264_, _21060_, _21059_);
  nand _54287_ (_21061_, _20587_, _28096_);
  nand _54288_ (_21062_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  nand _54289_ (_28335_, _21062_, _21061_);
  nand _54290_ (_21063_, _18286_, _24830_);
  nand _54291_ (_21064_, _18288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nand _54292_ (_11179_, _21064_, _21063_);
  nand _54293_ (_21065_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nand _54294_ (_21066_, _08329_, _25039_);
  nand _54295_ (_11181_, _21066_, _21065_);
  nand _54296_ (_21067_, _08331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  nand _54297_ (_21068_, _08329_, _25203_);
  nand _54298_ (_11183_, _21068_, _21067_);
  nor _54299_ (_21069_, _00269_, _24920_);
  nor _54300_ (_21070_, _00280_, _20255_);
  nor _54301_ (_21071_, _00282_, _00161_);
  nor _54302_ (_21072_, _21071_, _21070_);
  nand _54303_ (_21073_, _21072_, _00269_);
  nand _54304_ (_21074_, _21073_, _26487_);
  nor _54305_ (_11185_, _21074_, _21069_);
  nand _54306_ (_21075_, _04312_, _24830_);
  nand _54307_ (_21076_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  nand _54308_ (_11187_, _21076_, _21075_);
  nand _54309_ (_21077_, _20792_, _24789_);
  nand _54310_ (_21078_, _20794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  nand _54311_ (_11189_, _21078_, _21077_);
  nand _54312_ (_21079_, _20587_, _25039_);
  nand _54313_ (_21080_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nand _54314_ (_28336_, _21080_, _21079_);
  nand _54315_ (_21081_, _01182_, _24789_);
  nand _54316_ (_21082_, _01185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  nand _54317_ (_11193_, _21082_, _21081_);
  nand _54318_ (_21083_, _04312_, _24927_);
  nand _54319_ (_21084_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  nand _54320_ (_11196_, _21084_, _21083_);
  nand _54321_ (_21085_, _20814_, _24830_);
  nand _54322_ (_21086_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  nand _54323_ (_28356_, _21086_, _21085_);
  nand _54324_ (_21087_, _25000_, _24927_);
  nand _54325_ (_21088_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  nand _54326_ (_11203_, _21088_, _21087_);
  nand _54327_ (_21089_, _20587_, _24927_);
  nand _54328_ (_21090_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  nand _54329_ (_11208_, _21090_, _21089_);
  nand _54330_ (_21092_, _28096_, _25000_);
  nand _54331_ (_21093_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  nand _54332_ (_11210_, _21093_, _21092_);
  nand _54333_ (_21094_, _20814_, _25099_);
  nand _54334_ (_21095_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nand _54335_ (_11212_, _21095_, _21094_);
  nor _54336_ (_21096_, _00269_, _25194_);
  nor _54337_ (_21097_, _00280_, _20322_);
  nor _54338_ (_21098_, _00282_, _00171_);
  nor _54339_ (_21099_, _21098_, _21097_);
  nand _54340_ (_21100_, _21099_, _00269_);
  nand _54341_ (_21101_, _21100_, _26487_);
  nor _54342_ (_11214_, _21101_, _21096_);
  nand _54343_ (_21102_, _00479_, _25203_);
  nand _54344_ (_21103_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  nand _54345_ (_11218_, _21103_, _21102_);
  nand _54346_ (_21104_, _20587_, _24789_);
  nand _54347_ (_21105_, _20589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  nand _54348_ (_11221_, _21105_, _21104_);
  nand _54349_ (_21106_, _20814_, _28096_);
  nand _54350_ (_21107_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  nand _54351_ (_11223_, _21107_, _21106_);
  nor _54352_ (_21108_, _07942_, _25028_);
  nand _54353_ (_21109_, _07975_, _07961_);
  nand _54354_ (_21110_, _21109_, _07977_);
  nor _54355_ (_21111_, _21110_, _17060_);
  nand _54356_ (_21112_, _17060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _54357_ (_21113_, _20892_, _18671_);
  nor _54358_ (_21114_, _21113_, _18554_);
  nand _54359_ (_21115_, _21114_, _07983_);
  nand _54360_ (_21116_, _21115_, _21112_);
  nor _54361_ (_21117_, _21116_, _21111_);
  nand _54362_ (_21118_, _21117_, _07942_);
  nand _54363_ (_21119_, _21118_, _26487_);
  nor _54364_ (_11226_, _21119_, _21108_);
  nand _54365_ (_21120_, _20618_, _24830_);
  nand _54366_ (_21121_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nand _54367_ (_28337_, _21121_, _21120_);
  nand _54368_ (_21122_, _18533_, _24789_);
  nand _54369_ (_21123_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  nand _54370_ (_11228_, _21123_, _21122_);
  nand _54371_ (_21124_, _20814_, _25203_);
  nand _54372_ (_21125_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nand _54373_ (_28357_, _21125_, _21124_);
  nand _54374_ (_21126_, _20618_, _28096_);
  nand _54375_ (_21127_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nand _54376_ (_11231_, _21127_, _21126_);
  nand _54377_ (_21128_, _24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  nand _54378_ (_21129_, _25203_, _24796_);
  nand _54379_ (_11233_, _21129_, _21128_);
  nand _54380_ (_21131_, _19068_, _25203_);
  nand _54381_ (_21132_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nand _54382_ (_11238_, _21132_, _21131_);
  nand _54383_ (_21133_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  nand _54384_ (_21134_, _08549_, _25203_);
  nand _54385_ (_11240_, _21134_, _21133_);
  not _54386_ (_21135_, _04587_);
  nand _54387_ (_21136_, _24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nand _54388_ (_11244_, _21136_, _21135_);
  nand _54389_ (_21137_, _18533_, _25150_);
  nand _54390_ (_21138_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nand _54391_ (_11247_, _21138_, _21137_);
  nand _54392_ (_21139_, _18533_, _24927_);
  nand _54393_ (_21140_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  nand _54394_ (_11249_, _21140_, _21139_);
  nand _54395_ (_21141_, _20814_, _25039_);
  nand _54396_ (_21142_, _20816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  nand _54397_ (_28358_, _21142_, _21141_);
  nand _54398_ (_21143_, _20618_, _25203_);
  nand _54399_ (_21144_, _20620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  nand _54400_ (_11252_, _21144_, _21143_);
  nand _54401_ (_21145_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  nand _54402_ (_21146_, _08549_, _24927_);
  nand _54403_ (_28301_, _21146_, _21145_);
  nand _54404_ (_21147_, _25152_, _25099_);
  nand _54405_ (_21148_, _25154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nand _54406_ (_11257_, _21148_, _21147_);
  nand _54407_ (_21149_, _18157_, _24789_);
  nand _54408_ (_21150_, _18159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  nand _54409_ (_11262_, _21150_, _21149_);
  nand _54410_ (_21151_, _20763_, _24830_);
  nand _54411_ (_21152_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nand _54412_ (_11266_, _21152_, _21151_);
  nand _54413_ (_21153_, _20610_, _24789_);
  nand _54414_ (_21154_, _20612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  nand _54415_ (_11268_, _21154_, _21153_);
  nand _54416_ (_21155_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  nand _54417_ (_21156_, _08549_, _25039_);
  nand _54418_ (_11270_, _21156_, _21155_);
  nand _54419_ (_21157_, _00632_, _24789_);
  nand _54420_ (_21158_, _00634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  nand _54421_ (_11272_, _21158_, _21157_);
  nand _54422_ (_21159_, _20763_, _28096_);
  nand _54423_ (_21160_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nand _54424_ (_11274_, _21160_, _21159_);
  nand _54425_ (_21161_, _20563_, _24830_);
  nand _54426_ (_21162_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  nand _54427_ (_11277_, _21162_, _21161_);
  nand _54428_ (_21163_, _03840_, _25150_);
  nand _54429_ (_21164_, _03842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nand _54430_ (_28316_, _21164_, _21163_);
  nand _54431_ (_21165_, _18173_, _24830_);
  nand _54432_ (_21166_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  nand _54433_ (_11280_, _21166_, _21165_);
  nand _54434_ (_21167_, _18537_, _25099_);
  nand _54435_ (_21168_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nand _54436_ (_11282_, _21168_, _21167_);
  nand _54437_ (_21169_, _08387_, _28096_);
  nand _54438_ (_21170_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nand _54439_ (_28285_, _21170_, _21169_);
  nor _54440_ (_21171_, _07942_, _25139_);
  nor _54441_ (_21172_, _07949_, _07951_);
  nor _54442_ (_21173_, _07987_, _18569_);
  nand _54443_ (_21174_, _07971_, _07951_);
  nand _54444_ (_21175_, _21174_, _07985_);
  nor _54445_ (_21176_, _21175_, _07947_);
  nor _54446_ (_21177_, _21176_, _21173_);
  nor _54447_ (_21178_, _21177_, _07948_);
  nor _54448_ (_21179_, _21178_, _21172_);
  nand _54449_ (_21180_, _21179_, _07942_);
  nand _54450_ (_21181_, _21180_, _26487_);
  nor _54451_ (_11285_, _21181_, _21171_);
  nand _54452_ (_21182_, _03868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  nand _54453_ (_21183_, _03867_, _28096_);
  nand _54454_ (_11287_, _21183_, _21182_);
  nand _54455_ (_21184_, _19024_, _25203_);
  nand _54456_ (_21185_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nand _54457_ (_11292_, _21185_, _21184_);
  nand _54458_ (_21186_, _20763_, _25039_);
  nand _54459_ (_21187_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  nand _54460_ (_11294_, _21187_, _21186_);
  nor _54461_ (_21188_, _07942_, _24920_);
  nor _54462_ (_21189_, _07949_, _07952_);
  not _54463_ (_21190_, _07947_);
  nand _54464_ (_21191_, _07969_, _07952_);
  nand _54465_ (_21192_, _21191_, _21190_);
  nor _54466_ (_21193_, _21192_, _07970_);
  nor _54467_ (_21194_, _17064_, _18552_);
  nor _54468_ (_21195_, _21194_, _21193_);
  nor _54469_ (_21196_, _21195_, _07948_);
  nor _54470_ (_21197_, _21196_, _21189_);
  nand _54471_ (_21198_, _21197_, _07942_);
  nand _54472_ (_21199_, _21198_, _26487_);
  nor _54473_ (_11295_, _21199_, _21188_);
  nand _54474_ (_21200_, _20563_, _25099_);
  nand _54475_ (_21201_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  nand _54476_ (_11298_, _21201_, _21200_);
  nand _54477_ (_21202_, _20563_, _25203_);
  nand _54478_ (_21203_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nand _54479_ (_11300_, _21203_, _21202_);
  nand _54480_ (_21204_, _18816_, _24830_);
  nand _54481_ (_21205_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  nand _54482_ (_11302_, _21205_, _21204_);
  nand _54483_ (_21206_, _20763_, _24927_);
  nand _54484_ (_21207_, _20765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  nand _54485_ (_28361_, _21207_, _21206_);
  nand _54486_ (_21208_, _18537_, _25203_);
  nand _54487_ (_21209_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  nand _54488_ (_11305_, _21209_, _21208_);
  nand _54489_ (_21210_, _20563_, _25039_);
  nand _54490_ (_21211_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  nand _54491_ (_11308_, _21211_, _21210_);
  nand _54492_ (_21212_, _18537_, _28096_);
  nand _54493_ (_21213_, _18539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nand _54494_ (_11310_, _21213_, _21212_);
  nand _54495_ (_21214_, _18816_, _25039_);
  nand _54496_ (_21215_, _18818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nand _54497_ (_11313_, _21215_, _21214_);
  nand _54498_ (_21216_, _20757_, _25099_);
  nand _54499_ (_21217_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nand _54500_ (_11315_, _21217_, _21216_);
  nand _54501_ (_21218_, _18519_, _25099_);
  nand _54502_ (_21219_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nand _54503_ (_11317_, _21219_, _21218_);
  nand _54504_ (_21220_, _20563_, _24927_);
  nand _54505_ (_21221_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  nand _54506_ (_11321_, _21221_, _21220_);
  nand _54507_ (_21222_, _20757_, _25203_);
  nand _54508_ (_21223_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  nand _54509_ (_11324_, _21223_, _21222_);
  nand _54510_ (_21224_, _25150_, _24890_);
  nand _54511_ (_21225_, _24929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  nand _54512_ (_11326_, _21225_, _21224_);
  nand _54513_ (_21226_, _20563_, _24789_);
  nand _54514_ (_21227_, _20565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  nand _54515_ (_11328_, _21227_, _21226_);
  nand _54516_ (_21228_, _18871_, _28096_);
  nand _54517_ (_21229_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nand _54518_ (_11330_, _21229_, _21228_);
  nand _54519_ (_21230_, _19068_, _24927_);
  nand _54520_ (_21231_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  nand _54521_ (_28369_, _21231_, _21230_);
  nand _54522_ (_21232_, _18871_, _24830_);
  nand _54523_ (_21233_, _18873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nand _54524_ (_11332_, _21233_, _21232_);
  nand _54525_ (_21234_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  nand _54526_ (_21235_, _08549_, _24789_);
  nand _54527_ (_11335_, _21235_, _21234_);
  nand _54528_ (_21236_, _20757_, _25039_);
  nand _54529_ (_21237_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nand _54530_ (_11340_, _21237_, _21236_);
  nand _54531_ (_21238_, _00282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nand _54532_ (_21239_, _00280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _54533_ (_21240_, _21239_, _21238_);
  nor _54534_ (_21241_, _21240_, _00268_);
  nand _54535_ (_21242_, _00268_, _25088_);
  nand _54536_ (_21243_, _21242_, _26487_);
  nor _54537_ (_11343_, _21243_, _21241_);
  nor _54538_ (_21244_, _00269_, _25680_);
  nor _54539_ (_21245_, _00280_, _20531_);
  nor _54540_ (_21246_, _00282_, _00191_);
  nor _54541_ (_21247_, _21246_, _21245_);
  nand _54542_ (_21248_, _21247_, _00269_);
  nand _54543_ (_21249_, _21248_, _26487_);
  nor _54544_ (_11346_, _21249_, _21244_);
  nand _54545_ (_21250_, _18533_, _24830_);
  nand _54546_ (_21251_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nand _54547_ (_11348_, _21251_, _21250_);
  nand _54548_ (_21252_, _00280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _54549_ (_21253_, _00282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _54550_ (_21254_, _21253_, _21252_);
  nor _54551_ (_21255_, _21254_, _00268_);
  nand _54552_ (_21256_, _00268_, _24820_);
  nand _54553_ (_21257_, _21256_, _26487_);
  nor _54554_ (_11351_, _21257_, _21255_);
  nand _54555_ (_21258_, _03446_, _24927_);
  nand _54556_ (_21259_, _03449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand _54557_ (_11353_, _21259_, _21258_);
  nand _54558_ (_21260_, _20757_, _24789_);
  nand _54559_ (_21261_, _20759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  nand _54560_ (_11355_, _21261_, _21260_);
  nand _54561_ (_21262_, _20555_, _25099_);
  nand _54562_ (_21263_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nand _54563_ (_28341_, _21263_, _21262_);
  nand _54564_ (_21264_, _19024_, _25039_);
  nand _54565_ (_21265_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  nand _54566_ (_11362_, _21265_, _21264_);
  nand _54567_ (_21266_, _20751_, _24830_);
  nand _54568_ (_21267_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nand _54569_ (_11364_, _21267_, _21266_);
  nand _54570_ (_21269_, _03858_, _25150_);
  nand _54571_ (_21270_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  nand _54572_ (_11365_, _21270_, _21269_);
  nand _54573_ (_21271_, _20555_, _28096_);
  nand _54574_ (_21272_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nand _54575_ (_11367_, _21272_, _21271_);
  nand _54576_ (_21273_, _03858_, _28096_);
  nand _54577_ (_21274_, _03861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nand _54578_ (_11369_, _21274_, _21273_);
  nand _54579_ (_21275_, _20751_, _28096_);
  nand _54580_ (_21276_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nand _54581_ (_11371_, _21276_, _21275_);
  nand _54582_ (_21277_, _20555_, _25039_);
  nand _54583_ (_21278_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  nand _54584_ (_11377_, _21278_, _21277_);
  nand _54585_ (_21279_, _07908_, _28096_);
  nand _54586_ (_21280_, _07910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  nand _54587_ (_28325_, _21280_, _21279_);
  nand _54588_ (_21281_, _20555_, _25150_);
  nand _54589_ (_21282_, _20557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nand _54590_ (_11380_, _21282_, _21281_);
  nand _54591_ (_21284_, _04308_, _25039_);
  nand _54592_ (_21285_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  nand _54593_ (_11384_, _21285_, _21284_);
  nand _54594_ (_21286_, _20751_, _25203_);
  nand _54595_ (_21287_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  nand _54596_ (_28362_, _21287_, _21286_);
  nand _54597_ (_21288_, _04308_, _25099_);
  nand _54598_ (_21289_, _04310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  nand _54599_ (_11396_, _21289_, _21288_);
  nand _54600_ (_21290_, _20751_, _25150_);
  nand _54601_ (_21291_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nand _54602_ (_11399_, _21291_, _21290_);
  nand _54603_ (_21292_, _20543_, _24830_);
  nand _54604_ (_21293_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  nand _54605_ (_11403_, _21293_, _21292_);
  nand _54606_ (_21294_, _18135_, _24789_);
  nand _54607_ (_21295_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  nand _54608_ (_11415_, _21295_, _21294_);
  nand _54609_ (_21296_, _03822_, _25099_);
  nand _54610_ (_21297_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nand _54611_ (_11417_, _21297_, _21296_);
  nand _54612_ (_21298_, _03822_, _24789_);
  nand _54613_ (_21299_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  nand _54614_ (_11420_, _21299_, _21298_);
  nand _54615_ (_21300_, _20170_, _25099_);
  nand _54616_ (_21301_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  nand _54617_ (_11422_, _21301_, _21300_);
  nand _54618_ (_21302_, _20751_, _24789_);
  nand _54619_ (_21303_, _20753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  nand _54620_ (_11425_, _21303_, _21302_);
  nand _54621_ (_21305_, _20543_, _25099_);
  nand _54622_ (_21306_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  nand _54623_ (_11428_, _21306_, _21305_);
  nand _54624_ (_21307_, _20745_, _25099_);
  nand _54625_ (_21308_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  nand _54626_ (_28363_, _21308_, _21307_);
  nand _54627_ (_21309_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nand _54628_ (_21310_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand _54629_ (_21311_, _21310_, _21309_);
  nand _54630_ (_21312_, _21311_, _06717_);
  nand _54631_ (_21313_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nand _54632_ (_21314_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand _54633_ (_21315_, _21314_, _21313_);
  nand _54634_ (_21316_, _21315_, _06716_);
  nand _54635_ (_21317_, _21316_, _21312_);
  nand _54636_ (_21318_, _21317_, _06748_);
  nand _54637_ (_21319_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nand _54638_ (_21320_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand _54639_ (_21321_, _21320_, _21319_);
  nand _54640_ (_21322_, _21321_, _06717_);
  nand _54641_ (_21323_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nand _54642_ (_21324_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand _54643_ (_21325_, _21324_, _21323_);
  nand _54644_ (_21326_, _21325_, _06716_);
  nand _54645_ (_21327_, _21326_, _21322_);
  nand _54646_ (_21328_, _21327_, _06751_);
  nand _54647_ (_21329_, _21328_, _21318_);
  nand _54648_ (_21330_, _21329_, _06761_);
  nor _54649_ (_21331_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _54650_ (_21332_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _54651_ (_21333_, _21332_, _21331_);
  nand _54652_ (_21334_, _21333_, _06716_);
  nand _54653_ (_21335_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand _54654_ (_21336_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nand _54655_ (_21337_, _21336_, _21335_);
  nand _54656_ (_21338_, _21337_, _06717_);
  nand _54657_ (_21339_, _21338_, _21334_);
  nand _54658_ (_21340_, _21339_, _06748_);
  nor _54659_ (_21341_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _54660_ (_21342_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor _54661_ (_21343_, _21342_, _21341_);
  nand _54662_ (_21344_, _21343_, _06716_);
  nand _54663_ (_21345_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand _54664_ (_21346_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nand _54665_ (_21347_, _21346_, _21345_);
  nand _54666_ (_21348_, _21347_, _06717_);
  nand _54667_ (_21349_, _21348_, _21344_);
  nand _54668_ (_21350_, _21349_, _06751_);
  nand _54669_ (_21351_, _21350_, _21340_);
  nand _54670_ (_21352_, _21351_, _06760_);
  nand _54671_ (_21353_, _21352_, _21330_);
  nand _54672_ (_21354_, _21353_, _06780_);
  nand _54673_ (_21355_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  nand _54674_ (_21356_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  nand _54675_ (_21357_, _21356_, _21355_);
  nand _54676_ (_21358_, _21357_, _06717_);
  nand _54677_ (_21359_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  nand _54678_ (_21360_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  nand _54679_ (_21361_, _21360_, _21359_);
  nand _54680_ (_21362_, _21361_, _06716_);
  nand _54681_ (_21363_, _21362_, _21358_);
  nand _54682_ (_21364_, _21363_, _06748_);
  nand _54683_ (_21365_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  nand _54684_ (_21366_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  nand _54685_ (_21367_, _21366_, _21365_);
  nand _54686_ (_21368_, _21367_, _06717_);
  nand _54687_ (_21369_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nand _54688_ (_21370_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  nand _54689_ (_21371_, _21370_, _21369_);
  nand _54690_ (_21372_, _21371_, _06716_);
  nand _54691_ (_21373_, _21372_, _21368_);
  nand _54692_ (_21374_, _21373_, _06751_);
  nand _54693_ (_21375_, _21374_, _21364_);
  nand _54694_ (_21376_, _21375_, _06761_);
  nor _54695_ (_21377_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  nor _54696_ (_21378_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nor _54697_ (_21379_, _21378_, _21377_);
  nand _54698_ (_21380_, _21379_, _06717_);
  nor _54699_ (_21381_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  nor _54700_ (_21382_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  nor _54701_ (_21383_, _21382_, _21381_);
  nand _54702_ (_21384_, _21383_, _06716_);
  nand _54703_ (_21385_, _21384_, _21380_);
  nand _54704_ (_21386_, _21385_, _06748_);
  nor _54705_ (_21387_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  nor _54706_ (_21388_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nor _54707_ (_21389_, _21388_, _21387_);
  nand _54708_ (_21390_, _21389_, _06717_);
  nor _54709_ (_21391_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  nor _54710_ (_21392_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  nor _54711_ (_21393_, _21392_, _21391_);
  nand _54712_ (_21394_, _21393_, _06716_);
  nand _54713_ (_21395_, _21394_, _21390_);
  nand _54714_ (_21396_, _21395_, _06751_);
  nand _54715_ (_21397_, _21396_, _21386_);
  nand _54716_ (_21398_, _21397_, _06760_);
  nand _54717_ (_21399_, _21398_, _21376_);
  nand _54718_ (_21400_, _21399_, _06731_);
  nand _54719_ (_21401_, _21400_, _21354_);
  nand _54720_ (_21402_, _21401_, _06733_);
  nand _54721_ (_21403_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  nand _54722_ (_21404_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  nand _54723_ (_21405_, _21404_, _21403_);
  nand _54724_ (_21406_, _21405_, _06717_);
  nand _54725_ (_21407_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  nand _54726_ (_21408_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  nand _54727_ (_21409_, _21408_, _21407_);
  nand _54728_ (_21410_, _21409_, _06716_);
  nand _54729_ (_21411_, _21410_, _21406_);
  nand _54730_ (_21412_, _21411_, _06748_);
  nand _54731_ (_21413_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  nand _54732_ (_21414_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  nand _54733_ (_21415_, _21414_, _21413_);
  nand _54734_ (_21416_, _21415_, _06717_);
  nand _54735_ (_21417_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nand _54736_ (_21418_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  nand _54737_ (_21419_, _21418_, _21417_);
  nand _54738_ (_21420_, _21419_, _06716_);
  nand _54739_ (_21421_, _21420_, _21416_);
  nand _54740_ (_21422_, _21421_, _06751_);
  nand _54741_ (_21423_, _21422_, _21412_);
  nand _54742_ (_21424_, _21423_, _06761_);
  nor _54743_ (_21425_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  nor _54744_ (_21426_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  nor _54745_ (_21427_, _21426_, _21425_);
  nand _54746_ (_21428_, _21427_, _06717_);
  nor _54747_ (_21429_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  nor _54748_ (_21430_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  nor _54749_ (_21431_, _21430_, _21429_);
  nand _54750_ (_21432_, _21431_, _06716_);
  nand _54751_ (_21433_, _21432_, _21428_);
  nand _54752_ (_21434_, _21433_, _06748_);
  nor _54753_ (_21435_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  nor _54754_ (_21436_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nor _54755_ (_21437_, _21436_, _21435_);
  nand _54756_ (_21438_, _21437_, _06717_);
  nor _54757_ (_21439_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  nor _54758_ (_21440_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  nor _54759_ (_21441_, _21440_, _21439_);
  nand _54760_ (_21442_, _21441_, _06716_);
  nand _54761_ (_21443_, _21442_, _21438_);
  nand _54762_ (_21444_, _21443_, _06751_);
  nand _54763_ (_21445_, _21444_, _21434_);
  nand _54764_ (_21446_, _21445_, _06760_);
  nand _54765_ (_21447_, _21446_, _21424_);
  nand _54766_ (_21448_, _21447_, _06731_);
  nand _54767_ (_21449_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  nand _54768_ (_21450_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  nand _54769_ (_21451_, _21450_, _21449_);
  nand _54770_ (_21452_, _21451_, _06717_);
  nand _54771_ (_21453_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  nand _54772_ (_21454_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  nand _54773_ (_21455_, _21454_, _21453_);
  nand _54774_ (_21456_, _21455_, _06716_);
  nand _54775_ (_21457_, _21456_, _21452_);
  nand _54776_ (_21458_, _21457_, _06748_);
  nand _54777_ (_21459_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  nand _54778_ (_21460_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  nand _54779_ (_21461_, _21460_, _21459_);
  nand _54780_ (_21462_, _21461_, _06717_);
  nand _54781_ (_21463_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  nand _54782_ (_21464_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  nand _54783_ (_21465_, _21464_, _21463_);
  nand _54784_ (_21466_, _21465_, _06716_);
  nand _54785_ (_21467_, _21466_, _21462_);
  nand _54786_ (_21468_, _21467_, _06751_);
  nand _54787_ (_21469_, _21468_, _21458_);
  nand _54788_ (_21470_, _21469_, _06761_);
  nor _54789_ (_21471_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  nor _54790_ (_21472_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  nor _54791_ (_21473_, _21472_, _21471_);
  nand _54792_ (_21474_, _21473_, _06716_);
  nand _54793_ (_21475_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  nand _54794_ (_21476_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  nand _54795_ (_21477_, _21476_, _21475_);
  nand _54796_ (_21478_, _21477_, _06717_);
  nand _54797_ (_21479_, _21478_, _21474_);
  nand _54798_ (_21480_, _21479_, _06748_);
  nor _54799_ (_21481_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  nor _54800_ (_21482_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  nor _54801_ (_21483_, _21482_, _21481_);
  nand _54802_ (_21484_, _21483_, _06716_);
  nand _54803_ (_21485_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  nand _54804_ (_21486_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  nand _54805_ (_21487_, _21486_, _21485_);
  nand _54806_ (_21488_, _21487_, _06717_);
  nand _54807_ (_21489_, _21488_, _21484_);
  nand _54808_ (_21490_, _21489_, _06751_);
  nand _54809_ (_21491_, _21490_, _21480_);
  nand _54810_ (_21492_, _21491_, _06760_);
  nand _54811_ (_21493_, _21492_, _21470_);
  nand _54812_ (_21494_, _21493_, _06780_);
  nand _54813_ (_21495_, _21494_, _21448_);
  nand _54814_ (_21496_, _21495_, _06734_);
  nand _54815_ (_21497_, _21496_, _21402_);
  nand _54816_ (_21498_, _21497_, _13106_);
  nor _54817_ (_21499_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  nor _54818_ (_21500_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  nor _54819_ (_21501_, _21500_, _21499_);
  nand _54820_ (_21502_, _21501_, _06717_);
  nor _54821_ (_21503_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  nor _54822_ (_21504_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  nor _54823_ (_21505_, _21504_, _21503_);
  nand _54824_ (_21506_, _21505_, _06716_);
  nand _54825_ (_21507_, _21506_, _21502_);
  nand _54826_ (_21508_, _21507_, _06751_);
  nor _54827_ (_21509_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  nor _54828_ (_21510_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  nor _54829_ (_21511_, _21510_, _21509_);
  nand _54830_ (_21512_, _21511_, _06717_);
  nor _54831_ (_21513_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  nor _54832_ (_21514_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  nor _54833_ (_21515_, _21514_, _21513_);
  nand _54834_ (_21516_, _21515_, _06716_);
  nand _54835_ (_21517_, _21516_, _21512_);
  nand _54836_ (_21518_, _21517_, _06748_);
  nand _54837_ (_21519_, _21518_, _21508_);
  nand _54838_ (_21520_, _21519_, _06760_);
  nand _54839_ (_21521_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  nand _54840_ (_21522_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  nand _54841_ (_21523_, _21522_, _21521_);
  nand _54842_ (_21524_, _21523_, _06717_);
  nand _54843_ (_21525_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  nand _54844_ (_21526_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  nand _54845_ (_21527_, _21526_, _21525_);
  nand _54846_ (_21528_, _21527_, _06716_);
  nand _54847_ (_21529_, _21528_, _21524_);
  nand _54848_ (_21530_, _21529_, _06751_);
  nand _54849_ (_21531_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  nand _54850_ (_21532_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  nand _54851_ (_21533_, _21532_, _21531_);
  nand _54852_ (_21534_, _21533_, _06717_);
  nand _54853_ (_21535_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  nand _54854_ (_21536_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  nand _54855_ (_21537_, _21536_, _21535_);
  nand _54856_ (_21538_, _21537_, _06716_);
  nand _54857_ (_21539_, _21538_, _21534_);
  nand _54858_ (_21540_, _21539_, _06748_);
  nand _54859_ (_21541_, _21540_, _21530_);
  nand _54860_ (_21542_, _21541_, _06761_);
  nand _54861_ (_21543_, _21542_, _21520_);
  nand _54862_ (_21544_, _21543_, _06731_);
  nor _54863_ (_21545_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  nor _54864_ (_21546_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  nor _54865_ (_21547_, _21546_, _21545_);
  nand _54866_ (_21548_, _21547_, _06716_);
  nand _54867_ (_21549_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  nand _54868_ (_21550_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  nand _54869_ (_21551_, _21550_, _21549_);
  nand _54870_ (_21552_, _21551_, _06717_);
  nand _54871_ (_21553_, _21552_, _21548_);
  nand _54872_ (_21554_, _21553_, _06751_);
  nor _54873_ (_21555_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  nor _54874_ (_21556_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  nor _54875_ (_21557_, _21556_, _21555_);
  nand _54876_ (_21558_, _21557_, _06716_);
  nand _54877_ (_21559_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  nand _54878_ (_21560_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  nand _54879_ (_21561_, _21560_, _21559_);
  nand _54880_ (_21562_, _21561_, _06717_);
  nand _54881_ (_21563_, _21562_, _21558_);
  nand _54882_ (_21564_, _21563_, _06748_);
  nand _54883_ (_21565_, _21564_, _21554_);
  nand _54884_ (_21566_, _21565_, _06760_);
  nand _54885_ (_21567_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  nand _54886_ (_21568_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  nand _54887_ (_21569_, _21568_, _21567_);
  nand _54888_ (_21570_, _21569_, _06717_);
  nand _54889_ (_21571_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  nand _54890_ (_21573_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  nand _54891_ (_21574_, _21573_, _21571_);
  nand _54892_ (_21575_, _21574_, _06716_);
  nand _54893_ (_21576_, _21575_, _21570_);
  nand _54894_ (_21577_, _21576_, _06751_);
  nand _54895_ (_21578_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  nand _54896_ (_21579_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nand _54897_ (_21580_, _21579_, _21578_);
  nand _54898_ (_21581_, _21580_, _06717_);
  nand _54899_ (_21582_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  nand _54900_ (_21583_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  nand _54901_ (_21584_, _21583_, _21582_);
  nand _54902_ (_21585_, _21584_, _06716_);
  nand _54903_ (_21586_, _21585_, _21581_);
  nand _54904_ (_21587_, _21586_, _06748_);
  nand _54905_ (_21588_, _21587_, _21577_);
  nand _54906_ (_21589_, _21588_, _06761_);
  nand _54907_ (_21590_, _21589_, _21566_);
  nand _54908_ (_21591_, _21590_, _06780_);
  nand _54909_ (_21592_, _21591_, _21544_);
  nand _54910_ (_21593_, _21592_, _06733_);
  nand _54911_ (_21594_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  nand _54912_ (_21595_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  nand _54913_ (_21596_, _21595_, _21594_);
  nand _54914_ (_21597_, _21596_, _06717_);
  nand _54915_ (_21598_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  nand _54916_ (_21599_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  nand _54917_ (_21600_, _21599_, _21598_);
  nand _54918_ (_21601_, _21600_, _06716_);
  nand _54919_ (_21602_, _21601_, _21597_);
  nand _54920_ (_21603_, _21602_, _06748_);
  nand _54921_ (_21604_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  nand _54922_ (_21605_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  nand _54923_ (_21606_, _21605_, _21604_);
  nand _54924_ (_21607_, _21606_, _06717_);
  nand _54925_ (_21608_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  nand _54926_ (_21609_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  nand _54927_ (_21610_, _21609_, _21608_);
  nand _54928_ (_21611_, _21610_, _06716_);
  nand _54929_ (_21612_, _21611_, _21607_);
  nand _54930_ (_21613_, _21612_, _06751_);
  nand _54931_ (_21614_, _21613_, _21603_);
  nand _54932_ (_21615_, _21614_, _06761_);
  nor _54933_ (_21616_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  nor _54934_ (_21617_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  nor _54935_ (_21618_, _21617_, _21616_);
  nand _54936_ (_21619_, _21618_, _06716_);
  nand _54937_ (_21620_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  nand _54938_ (_21621_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  nand _54939_ (_21622_, _21621_, _21620_);
  nand _54940_ (_21624_, _21622_, _06717_);
  nand _54941_ (_21625_, _21624_, _21619_);
  nand _54942_ (_21626_, _21625_, _06748_);
  nor _54943_ (_21627_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  nor _54944_ (_21628_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nor _54945_ (_21629_, _21628_, _21627_);
  nand _54946_ (_21630_, _21629_, _06716_);
  nand _54947_ (_21631_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  nand _54948_ (_21632_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  nand _54949_ (_21633_, _21632_, _21631_);
  nand _54950_ (_21634_, _21633_, _06717_);
  nand _54951_ (_21635_, _21634_, _21630_);
  nand _54952_ (_21636_, _21635_, _06751_);
  nand _54953_ (_21637_, _21636_, _21626_);
  nand _54954_ (_21638_, _21637_, _06760_);
  nand _54955_ (_21639_, _21638_, _21615_);
  nand _54956_ (_21640_, _21639_, _06780_);
  nand _54957_ (_21641_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  nand _54958_ (_21642_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  nand _54959_ (_21643_, _21642_, _21641_);
  nand _54960_ (_21644_, _21643_, _06717_);
  nand _54961_ (_21645_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  nand _54962_ (_21646_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  nand _54963_ (_21647_, _21646_, _21645_);
  nand _54964_ (_21648_, _21647_, _06716_);
  nand _54965_ (_21649_, _21648_, _21644_);
  nand _54966_ (_21650_, _21649_, _06748_);
  nand _54967_ (_21651_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  nand _54968_ (_21652_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  nand _54969_ (_21653_, _21652_, _21651_);
  nand _54970_ (_21655_, _21653_, _06717_);
  nand _54971_ (_21656_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  nand _54972_ (_21657_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  nand _54973_ (_21658_, _21657_, _21656_);
  nand _54974_ (_21659_, _21658_, _06716_);
  nand _54975_ (_21660_, _21659_, _21655_);
  nand _54976_ (_21661_, _21660_, _06751_);
  nand _54977_ (_21662_, _21661_, _21650_);
  nand _54978_ (_21663_, _21662_, _06761_);
  nor _54979_ (_21664_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  nor _54980_ (_21665_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nor _54981_ (_21666_, _21665_, _21664_);
  nand _54982_ (_21667_, _21666_, _06717_);
  nor _54983_ (_21668_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  nor _54984_ (_21669_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  nor _54985_ (_21670_, _21669_, _21668_);
  nand _54986_ (_21671_, _21670_, _06716_);
  nand _54987_ (_21672_, _21671_, _21667_);
  nand _54988_ (_21673_, _21672_, _06748_);
  nor _54989_ (_21674_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  nor _54990_ (_21675_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  nor _54991_ (_21676_, _21675_, _21674_);
  nand _54992_ (_21677_, _21676_, _06717_);
  nor _54993_ (_21678_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  nor _54994_ (_21679_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nor _54995_ (_21680_, _21679_, _21678_);
  nand _54996_ (_21681_, _21680_, _06716_);
  nand _54997_ (_21682_, _21681_, _21677_);
  nand _54998_ (_21683_, _21682_, _06751_);
  nand _54999_ (_21684_, _21683_, _21673_);
  nand _55000_ (_21685_, _21684_, _06760_);
  nand _55001_ (_21686_, _21685_, _21663_);
  nand _55002_ (_21687_, _21686_, _06731_);
  nand _55003_ (_21688_, _21687_, _21640_);
  nand _55004_ (_21689_, _21688_, _06734_);
  nand _55005_ (_21690_, _21689_, _21593_);
  nand _55006_ (_21691_, _21690_, _06723_);
  nand _55007_ (_21692_, _21691_, _21498_);
  nor _55008_ (_21693_, _21692_, _25929_);
  nand _55009_ (_21694_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  nand _55010_ (_21695_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  nand _55011_ (_21696_, _21695_, _21694_);
  nand _55012_ (_21697_, _21696_, _06716_);
  nand _55013_ (_21698_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  nand _55014_ (_21699_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  nand _55015_ (_21700_, _21699_, _21698_);
  nand _55016_ (_21701_, _21700_, _06717_);
  nand _55017_ (_21702_, _21701_, _21697_);
  nand _55018_ (_21703_, _21702_, _06748_);
  nand _55019_ (_21704_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  nand _55020_ (_21705_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  nand _55021_ (_21706_, _21705_, _21704_);
  nand _55022_ (_21707_, _21706_, _06716_);
  nand _55023_ (_21708_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  nand _55024_ (_21709_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  nand _55025_ (_21710_, _21709_, _21708_);
  nand _55026_ (_21711_, _21710_, _06717_);
  nand _55027_ (_21712_, _21711_, _21707_);
  nand _55028_ (_21713_, _21712_, _06751_);
  nand _55029_ (_21714_, _21713_, _21703_);
  nand _55030_ (_21715_, _21714_, _06761_);
  nand _55031_ (_21716_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  nand _55032_ (_21717_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  nand _55033_ (_21718_, _21717_, _21716_);
  nand _55034_ (_21719_, _21718_, _06717_);
  nor _55035_ (_21720_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  nor _55036_ (_21721_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  nor _55037_ (_21722_, _21721_, _21720_);
  nand _55038_ (_21723_, _21722_, _06716_);
  nand _55039_ (_21724_, _21723_, _21719_);
  nand _55040_ (_21725_, _21724_, _06748_);
  nand _55041_ (_21726_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  nand _55042_ (_21727_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  nand _55043_ (_21728_, _21727_, _21726_);
  nand _55044_ (_21729_, _21728_, _06717_);
  nor _55045_ (_21730_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  nor _55046_ (_21731_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  nor _55047_ (_21732_, _21731_, _21730_);
  nand _55048_ (_21733_, _21732_, _06716_);
  nand _55049_ (_21734_, _21733_, _21729_);
  nand _55050_ (_21735_, _21734_, _06751_);
  nand _55051_ (_21736_, _21735_, _21725_);
  nand _55052_ (_21737_, _21736_, _06760_);
  nand _55053_ (_21738_, _21737_, _21715_);
  nand _55054_ (_21739_, _21738_, _06780_);
  nand _55055_ (_21740_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  nand _55056_ (_21741_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  nand _55057_ (_21742_, _21741_, _21740_);
  nand _55058_ (_21743_, _21742_, _06717_);
  nand _55059_ (_21744_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  nand _55060_ (_21745_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  nand _55061_ (_21746_, _21745_, _21744_);
  nand _55062_ (_21747_, _21746_, _06716_);
  nand _55063_ (_21748_, _21747_, _21743_);
  nand _55064_ (_21749_, _21748_, _06748_);
  nand _55065_ (_21750_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  nand _55066_ (_21751_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  nand _55067_ (_21752_, _21751_, _21750_);
  nand _55068_ (_21753_, _21752_, _06717_);
  nand _55069_ (_21754_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  nand _55070_ (_21755_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  nand _55071_ (_21756_, _21755_, _21754_);
  nand _55072_ (_21757_, _21756_, _06716_);
  nand _55073_ (_21758_, _21757_, _21753_);
  nand _55074_ (_21759_, _21758_, _06751_);
  nand _55075_ (_21760_, _21759_, _21749_);
  nand _55076_ (_21761_, _21760_, _06761_);
  nor _55077_ (_21762_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  nor _55078_ (_21763_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  nor _55079_ (_21764_, _21763_, _21762_);
  nand _55080_ (_21765_, _21764_, _06717_);
  nor _55081_ (_21766_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  nor _55082_ (_21767_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  nor _55083_ (_21768_, _21767_, _21766_);
  nand _55084_ (_21769_, _21768_, _06716_);
  nand _55085_ (_21770_, _21769_, _21765_);
  nand _55086_ (_21771_, _21770_, _06748_);
  nor _55087_ (_21772_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  nor _55088_ (_21773_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  nor _55089_ (_21774_, _21773_, _21772_);
  nor _55090_ (_21775_, _21774_, _06716_);
  nor _55091_ (_21776_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  nor _55092_ (_21777_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  nor _55093_ (_21778_, _21777_, _21776_);
  nor _55094_ (_21779_, _21778_, _06717_);
  nor _55095_ (_21780_, _21779_, _21775_);
  nand _55096_ (_21781_, _21780_, _06751_);
  nand _55097_ (_21782_, _21781_, _21771_);
  nand _55098_ (_21783_, _21782_, _06760_);
  nand _55099_ (_21784_, _21783_, _21761_);
  nand _55100_ (_21785_, _21784_, _06731_);
  nand _55101_ (_21786_, _21785_, _21739_);
  nand _55102_ (_21787_, _21786_, _06734_);
  nand _55103_ (_21788_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  nand _55104_ (_21789_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  nand _55105_ (_21790_, _21789_, _21788_);
  nand _55106_ (_21791_, _21790_, _06717_);
  nand _55107_ (_21792_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  nand _55108_ (_21793_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nand _55109_ (_21794_, _21793_, _21792_);
  nand _55110_ (_21795_, _21794_, _06716_);
  nand _55111_ (_21796_, _21795_, _21791_);
  nand _55112_ (_21797_, _21796_, _06748_);
  nand _55113_ (_21798_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  nand _55114_ (_21799_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  nand _55115_ (_21800_, _21799_, _21798_);
  nand _55116_ (_21801_, _21800_, _06717_);
  nand _55117_ (_21802_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  nand _55118_ (_21803_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  nand _55119_ (_21804_, _21803_, _21802_);
  nand _55120_ (_21805_, _21804_, _06716_);
  nand _55121_ (_21806_, _21805_, _21801_);
  nand _55122_ (_21807_, _21806_, _06751_);
  nand _55123_ (_21808_, _21807_, _21797_);
  nand _55124_ (_21809_, _21808_, _06761_);
  nor _55125_ (_21810_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  nor _55126_ (_21811_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  nor _55127_ (_21812_, _21811_, _21810_);
  nand _55128_ (_21813_, _21812_, _06717_);
  nor _55129_ (_21814_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  nor _55130_ (_21815_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  nor _55131_ (_21816_, _21815_, _21814_);
  nand _55132_ (_21817_, _21816_, _06716_);
  nand _55133_ (_21818_, _21817_, _21813_);
  nand _55134_ (_21819_, _21818_, _06748_);
  nor _55135_ (_21820_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  nor _55136_ (_21821_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  nor _55137_ (_21822_, _21821_, _21820_);
  nand _55138_ (_21823_, _21822_, _06717_);
  nor _55139_ (_21824_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  nor _55140_ (_21825_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  nor _55141_ (_21826_, _21825_, _21824_);
  nand _55142_ (_21827_, _21826_, _06716_);
  nand _55143_ (_21828_, _21827_, _21823_);
  nand _55144_ (_21829_, _21828_, _06751_);
  nand _55145_ (_21830_, _21829_, _21819_);
  nand _55146_ (_21831_, _21830_, _06760_);
  nand _55147_ (_21832_, _21831_, _21809_);
  nand _55148_ (_21833_, _21832_, _06780_);
  nand _55149_ (_21834_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  nand _55150_ (_21835_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  nand _55151_ (_21836_, _21835_, _21834_);
  nand _55152_ (_21837_, _21836_, _06717_);
  nand _55153_ (_21838_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  nand _55154_ (_21839_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  nand _55155_ (_21840_, _21839_, _21838_);
  nand _55156_ (_21841_, _21840_, _06716_);
  nand _55157_ (_21842_, _21841_, _21837_);
  nand _55158_ (_21843_, _21842_, _06748_);
  nand _55159_ (_21844_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  nand _55160_ (_21846_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  nand _55161_ (_21847_, _21846_, _21844_);
  nand _55162_ (_21848_, _21847_, _06717_);
  nand _55163_ (_21849_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  nand _55164_ (_21850_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  nand _55165_ (_21851_, _21850_, _21849_);
  nand _55166_ (_21852_, _21851_, _06716_);
  nand _55167_ (_21853_, _21852_, _21848_);
  nand _55168_ (_21854_, _21853_, _06751_);
  nand _55169_ (_21855_, _21854_, _21843_);
  nand _55170_ (_21856_, _21855_, _06761_);
  nor _55171_ (_21857_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  nor _55172_ (_21858_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  nor _55173_ (_21859_, _21858_, _21857_);
  nand _55174_ (_21860_, _21859_, _06717_);
  nor _55175_ (_21861_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  nor _55176_ (_21862_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  nor _55177_ (_21863_, _21862_, _21861_);
  nand _55178_ (_21864_, _21863_, _06716_);
  nand _55179_ (_21865_, _21864_, _21860_);
  nand _55180_ (_21866_, _21865_, _06748_);
  nor _55181_ (_21867_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  nor _55182_ (_21868_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  nor _55183_ (_21869_, _21868_, _21867_);
  nand _55184_ (_21870_, _21869_, _06717_);
  nor _55185_ (_21871_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nor _55186_ (_21872_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  nor _55187_ (_21873_, _21872_, _21871_);
  nand _55188_ (_21874_, _21873_, _06716_);
  nand _55189_ (_21875_, _21874_, _21870_);
  nand _55190_ (_21876_, _21875_, _06751_);
  nand _55191_ (_21877_, _21876_, _21866_);
  nand _55192_ (_21878_, _21877_, _06760_);
  nand _55193_ (_21879_, _21878_, _21856_);
  nand _55194_ (_21880_, _21879_, _06731_);
  nand _55195_ (_21881_, _21880_, _21833_);
  nand _55196_ (_21882_, _21881_, _06733_);
  nand _55197_ (_21883_, _21882_, _21787_);
  nand _55198_ (_21884_, _21883_, _13106_);
  nand _55199_ (_21885_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  nand _55200_ (_21886_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  nand _55201_ (_21887_, _21886_, _21885_);
  nand _55202_ (_21888_, _21887_, _06716_);
  nand _55203_ (_21889_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nand _55204_ (_21890_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  nand _55205_ (_21891_, _21890_, _21889_);
  nand _55206_ (_21892_, _21891_, _06717_);
  nand _55207_ (_21893_, _21892_, _21888_);
  nand _55208_ (_21894_, _21893_, _06748_);
  nand _55209_ (_21895_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  nand _55210_ (_21896_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  nand _55211_ (_21897_, _21896_, _21895_);
  nand _55212_ (_21898_, _21897_, _06716_);
  nand _55213_ (_21899_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  nand _55214_ (_21900_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  nand _55215_ (_21901_, _21900_, _21899_);
  nand _55216_ (_21902_, _21901_, _06717_);
  nand _55217_ (_21903_, _21902_, _21898_);
  nand _55218_ (_21904_, _21903_, _06751_);
  nand _55219_ (_21905_, _21904_, _21894_);
  nand _55220_ (_21906_, _21905_, _06761_);
  nand _55221_ (_21907_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  nand _55222_ (_21908_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  nand _55223_ (_21909_, _21908_, _21907_);
  nand _55224_ (_21910_, _21909_, _06717_);
  nor _55225_ (_21911_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  nor _55226_ (_21912_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  nor _55227_ (_21913_, _21912_, _21911_);
  nand _55228_ (_21914_, _21913_, _06716_);
  nand _55229_ (_21915_, _21914_, _21910_);
  nand _55230_ (_21916_, _21915_, _06748_);
  nand _55231_ (_21917_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  nand _55232_ (_21918_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  nand _55233_ (_21919_, _21918_, _21917_);
  nand _55234_ (_21920_, _21919_, _06717_);
  nor _55235_ (_21921_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  nor _55236_ (_21922_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  nor _55237_ (_21923_, _21922_, _21921_);
  nand _55238_ (_21924_, _21923_, _06716_);
  nand _55239_ (_21925_, _21924_, _21920_);
  nand _55240_ (_21926_, _21925_, _06751_);
  nand _55241_ (_21927_, _21926_, _21916_);
  nand _55242_ (_21928_, _21927_, _06760_);
  nand _55243_ (_21929_, _21928_, _21906_);
  nand _55244_ (_21930_, _21929_, _06780_);
  nand _55245_ (_21931_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  nand _55246_ (_21932_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  nand _55247_ (_21933_, _21932_, _21931_);
  nand _55248_ (_21934_, _21933_, _06717_);
  nand _55249_ (_21935_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  nand _55250_ (_21936_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nand _55251_ (_21937_, _21936_, _21935_);
  nand _55252_ (_21938_, _21937_, _06716_);
  nand _55253_ (_21939_, _21938_, _21934_);
  nand _55254_ (_21940_, _21939_, _06748_);
  nand _55255_ (_21941_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  nand _55256_ (_21942_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  nand _55257_ (_21943_, _21942_, _21941_);
  nand _55258_ (_21944_, _21943_, _06717_);
  nand _55259_ (_21945_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  nand _55260_ (_21946_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  nand _55261_ (_21947_, _21946_, _21945_);
  nand _55262_ (_21948_, _21947_, _06716_);
  nand _55263_ (_21949_, _21948_, _21944_);
  nand _55264_ (_21950_, _21949_, _06751_);
  nand _55265_ (_21951_, _21950_, _21940_);
  nand _55266_ (_21952_, _21951_, _06761_);
  nor _55267_ (_21953_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  nor _55268_ (_21954_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  nor _55269_ (_21955_, _21954_, _21953_);
  nand _55270_ (_21956_, _21955_, _06717_);
  nor _55271_ (_21957_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  nor _55272_ (_21958_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  nor _55273_ (_21959_, _21958_, _21957_);
  nand _55274_ (_21960_, _21959_, _06716_);
  nand _55275_ (_21961_, _21960_, _21956_);
  nand _55276_ (_21962_, _21961_, _06748_);
  nor _55277_ (_21963_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nor _55278_ (_21964_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  nor _55279_ (_21965_, _21964_, _21963_);
  nor _55280_ (_21966_, _21965_, _06716_);
  nor _55281_ (_21967_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  nor _55282_ (_21968_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  nor _55283_ (_21969_, _21968_, _21967_);
  nor _55284_ (_21970_, _21969_, _06717_);
  nor _55285_ (_21971_, _21970_, _21966_);
  nand _55286_ (_21972_, _21971_, _06751_);
  nand _55287_ (_21973_, _21972_, _21962_);
  nand _55288_ (_21974_, _21973_, _06760_);
  nand _55289_ (_21975_, _21974_, _21952_);
  nand _55290_ (_21976_, _21975_, _06731_);
  nand _55291_ (_21977_, _21976_, _21930_);
  nand _55292_ (_21978_, _21977_, _06734_);
  nand _55293_ (_21979_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  nand _55294_ (_21980_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  nand _55295_ (_21981_, _21980_, _21979_);
  nand _55296_ (_21982_, _21981_, _06717_);
  nand _55297_ (_21983_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nand _55298_ (_21984_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  nand _55299_ (_21985_, _21984_, _21983_);
  nand _55300_ (_21986_, _21985_, _06716_);
  nand _55301_ (_21987_, _21986_, _21982_);
  nand _55302_ (_21988_, _21987_, _06748_);
  nand _55303_ (_21989_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  nand _55304_ (_21990_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  nand _55305_ (_21991_, _21990_, _21989_);
  nand _55306_ (_21992_, _21991_, _06717_);
  nand _55307_ (_21993_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  nand _55308_ (_21994_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  nand _55309_ (_21995_, _21994_, _21993_);
  nand _55310_ (_21996_, _21995_, _06716_);
  nand _55311_ (_21997_, _21996_, _21992_);
  nand _55312_ (_21998_, _21997_, _06751_);
  nand _55313_ (_21999_, _21998_, _21988_);
  nand _55314_ (_22000_, _21999_, _06761_);
  nor _55315_ (_22001_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  nor _55316_ (_22002_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  nor _55317_ (_22003_, _22002_, _22001_);
  nand _55318_ (_22004_, _22003_, _06717_);
  nor _55319_ (_22005_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  nor _55320_ (_22006_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  nor _55321_ (_22007_, _22006_, _22005_);
  nand _55322_ (_22008_, _22007_, _06716_);
  nand _55323_ (_22009_, _22008_, _22004_);
  nand _55324_ (_22010_, _22009_, _06748_);
  nor _55325_ (_22011_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  nor _55326_ (_22012_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  nor _55327_ (_22013_, _22012_, _22011_);
  nand _55328_ (_22014_, _22013_, _06717_);
  nor _55329_ (_22015_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  nor _55330_ (_22017_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  nor _55331_ (_22018_, _22017_, _22015_);
  nand _55332_ (_22019_, _22018_, _06716_);
  nand _55333_ (_22020_, _22019_, _22014_);
  nand _55334_ (_22021_, _22020_, _06751_);
  nand _55335_ (_22022_, _22021_, _22010_);
  nand _55336_ (_22023_, _22022_, _06760_);
  nand _55337_ (_22024_, _22023_, _22000_);
  nand _55338_ (_22025_, _22024_, _06731_);
  nand _55339_ (_22026_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  nand _55340_ (_22027_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  nand _55341_ (_22028_, _22027_, _22026_);
  nand _55342_ (_22029_, _22028_, _06717_);
  nand _55343_ (_22030_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  nand _55344_ (_22031_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  nand _55345_ (_22032_, _22031_, _22030_);
  nand _55346_ (_22033_, _22032_, _06716_);
  nand _55347_ (_22034_, _22033_, _22029_);
  nand _55348_ (_22035_, _22034_, _06748_);
  nand _55349_ (_22036_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  nand _55350_ (_22037_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  nand _55351_ (_22038_, _22037_, _22036_);
  nand _55352_ (_22039_, _22038_, _06717_);
  nand _55353_ (_22040_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  nand _55354_ (_22041_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  nand _55355_ (_22042_, _22041_, _22040_);
  nand _55356_ (_22043_, _22042_, _06716_);
  nand _55357_ (_22044_, _22043_, _22039_);
  nand _55358_ (_22045_, _22044_, _06751_);
  nand _55359_ (_22046_, _22045_, _22035_);
  nand _55360_ (_22047_, _22046_, _06761_);
  nor _55361_ (_22048_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  nor _55362_ (_22049_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  nor _55363_ (_22050_, _22049_, _22048_);
  nand _55364_ (_22051_, _22050_, _06717_);
  nor _55365_ (_22052_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  nor _55366_ (_22053_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  nor _55367_ (_22054_, _22053_, _22052_);
  nand _55368_ (_22055_, _22054_, _06716_);
  nand _55369_ (_22056_, _22055_, _22051_);
  nand _55370_ (_22057_, _22056_, _06748_);
  nor _55371_ (_22058_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  nor _55372_ (_22059_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  nor _55373_ (_22060_, _22059_, _22058_);
  nand _55374_ (_22061_, _22060_, _06717_);
  nor _55375_ (_22062_, _06771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  nor _55376_ (_22063_, _06774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  nor _55377_ (_22064_, _22063_, _22062_);
  nand _55378_ (_22065_, _22064_, _06716_);
  nand _55379_ (_22066_, _22065_, _22061_);
  nand _55380_ (_22067_, _22066_, _06751_);
  nand _55381_ (_22068_, _22067_, _22057_);
  nand _55382_ (_22069_, _22068_, _06760_);
  nand _55383_ (_22070_, _22069_, _22047_);
  nand _55384_ (_22071_, _22070_, _06780_);
  nand _55385_ (_22072_, _22071_, _22025_);
  nand _55386_ (_22073_, _22072_, _06733_);
  nand _55387_ (_22074_, _22073_, _21978_);
  nand _55388_ (_22075_, _22074_, _06723_);
  nand _55389_ (_22076_, _22075_, _21884_);
  nor _55390_ (_22077_, _22076_, _25843_);
  nor _55391_ (_22078_, _22077_, _21693_);
  nor _55392_ (_22079_, _22078_, _13105_);
  nand _55393_ (_22080_, _13105_, _24180_);
  nand _55394_ (_22081_, _22080_, _26487_);
  nor _55395_ (_11433_, _22081_, _22079_);
  nand _55396_ (_22082_, _20543_, _25203_);
  nand _55397_ (_22083_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  nand _55398_ (_11442_, _22083_, _22082_);
  nand _55399_ (_22084_, _20170_, _24927_);
  nand _55400_ (_22085_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  nand _55401_ (_11444_, _22085_, _22084_);
  nor _55402_ (_28219_[7], _26523_, rst);
  nand _55403_ (_22086_, _20543_, _24927_);
  nand _55404_ (_22087_, _20545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  nand _55405_ (_11451_, _22087_, _22086_);
  nand _55406_ (_22088_, _20745_, _28096_);
  nand _55407_ (_22089_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  nand _55408_ (_11453_, _22089_, _22088_);
  nand _55409_ (_22090_, _20521_, _24830_);
  nand _55410_ (_22091_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nand _55411_ (_11459_, _22091_, _22090_);
  nand _55412_ (_22092_, _18058_, _25039_);
  nand _55413_ (_22093_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nand _55414_ (_11461_, _22093_, _22092_);
  nand _55415_ (_22094_, _20745_, _24927_);
  nand _55416_ (_22095_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  nand _55417_ (_11463_, _22095_, _22094_);
  nand _55418_ (_22096_, _18058_, _25099_);
  nand _55419_ (_22097_, _18060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  nand _55420_ (_11466_, _22097_, _22096_);
  nand _55421_ (_22098_, _20745_, _24789_);
  nand _55422_ (_22099_, _20747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  nand _55423_ (_28364_, _22099_, _22098_);
  nand _55424_ (_22100_, _20521_, _25099_);
  nand _55425_ (_22101_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nand _55426_ (_11472_, _22101_, _22100_);
  nand _55427_ (_22102_, _20735_, _24830_);
  nand _55428_ (_22103_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nand _55429_ (_11478_, _22103_, _22102_);
  nand _55430_ (_22104_, _20521_, _25203_);
  nand _55431_ (_22105_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nand _55432_ (_11481_, _22105_, _22104_);
  nand _55433_ (_22106_, _11827_, _24927_);
  nand _55434_ (_22107_, _11829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  nand _55435_ (_11483_, _22107_, _22106_);
  nand _55436_ (_22108_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nand _55437_ (_22109_, _08334_, _25150_);
  nand _55438_ (_11487_, _22109_, _22108_);
  nand _55439_ (_22110_, _20521_, _24927_);
  nand _55440_ (_22111_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  nand _55441_ (_11489_, _22111_, _22110_);
  nand _55442_ (_22112_, _04624_, _24927_);
  nand _55443_ (_22113_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  nand _55444_ (_11493_, _22113_, _22112_);
  nand _55445_ (_22114_, _20735_, _25099_);
  nand _55446_ (_22115_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  nand _55447_ (_11495_, _22115_, _22114_);
  nand _55448_ (_22116_, _04624_, _28096_);
  nand _55449_ (_22117_, _04626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nand _55450_ (_11497_, _22117_, _22116_);
  nand _55451_ (_22118_, _20735_, _25203_);
  nand _55452_ (_22119_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  nand _55453_ (_11499_, _22119_, _22118_);
  nand _55454_ (_22120_, _03834_, _24927_);
  nand _55455_ (_22121_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  nand _55456_ (_11501_, _22121_, _22120_);
  nand _55457_ (_22122_, _20521_, _24789_);
  nand _55458_ (_22123_, _20523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  nand _55459_ (_11504_, _22123_, _22122_);
  nand _55460_ (_22124_, _20735_, _25039_);
  nand _55461_ (_22125_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  nand _55462_ (_11507_, _22125_, _22124_);
  nand _55463_ (_22126_, _20511_, _24830_);
  nand _55464_ (_22127_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  nand _55465_ (_11509_, _22127_, _22126_);
  nand _55466_ (_22128_, _20735_, _24927_);
  nand _55467_ (_22129_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  nand _55468_ (_11514_, _22129_, _22128_);
  nand _55469_ (_22130_, _20511_, _28096_);
  nand _55470_ (_22131_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  nand _55471_ (_11515_, _22131_, _22130_);
  nor _55472_ (_28218_[7], _25837_, rst);
  nand _55473_ (_22132_, _20511_, _25039_);
  nand _55474_ (_22133_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  nand _55475_ (_11519_, _22133_, _22132_);
  nand _55476_ (_22134_, _20735_, _25150_);
  nand _55477_ (_22135_, _20737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nand _55478_ (_11521_, _22135_, _22134_);
  nand _55479_ (_22136_, _19094_, _24830_);
  nand _55480_ (_22137_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nand _55481_ (_11523_, _22137_, _22136_);
  nand _55482_ (_22138_, _20726_, _24830_);
  nand _55483_ (_22139_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  nand _55484_ (_11525_, _22139_, _22138_);
  nand _55485_ (_22140_, _20511_, _25150_);
  nand _55486_ (_22141_, _20513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  nand _55487_ (_11527_, _22141_, _22140_);
  nand _55488_ (_22142_, _20726_, _28096_);
  nand _55489_ (_22143_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  nand _55490_ (_11529_, _22143_, _22142_);
  nand _55491_ (_22144_, _19068_, _24789_);
  nand _55492_ (_22145_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  nand _55493_ (_11532_, _22145_, _22144_);
  nand _55494_ (_22146_, _19094_, _25039_);
  nand _55495_ (_22147_, _19096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  nand _55496_ (_11536_, _22147_, _22146_);
  nand _55497_ (_22148_, _18533_, _25203_);
  nand _55498_ (_22149_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nand _55499_ (_11538_, _22149_, _22148_);
  nand _55500_ (_22150_, _20726_, _25039_);
  nand _55501_ (_22151_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nand _55502_ (_11539_, _22151_, _22150_);
  nand _55503_ (_22152_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  nand _55504_ (_22153_, _08334_, _24927_);
  nand _55505_ (_28300_, _22153_, _22152_);
  nand _55506_ (_22154_, _18533_, _28096_);
  nand _55507_ (_22155_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  nand _55508_ (_28261_, _22155_, _22154_);
  nand _55509_ (_22156_, _18533_, _25099_);
  nand _55510_ (_22157_, _18535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  nand _55511_ (_11544_, _22157_, _22156_);
  nand _55512_ (_22158_, _20505_, _25099_);
  nand _55513_ (_22159_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nand _55514_ (_11546_, _22159_, _22158_);
  nand _55515_ (_22160_, _07882_, _25039_);
  nand _55516_ (_22161_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nand _55517_ (_11548_, _22161_, _22160_);
  nand _55518_ (_22162_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  nand _55519_ (_22163_, _08334_, _25039_);
  nand _55520_ (_11550_, _22163_, _22162_);
  nand _55521_ (_22164_, _07882_, _25099_);
  nand _55522_ (_22165_, _07884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  nand _55523_ (_11552_, _22165_, _22164_);
  nand _55524_ (_22166_, _20726_, _24927_);
  nand _55525_ (_22167_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  nand _55526_ (_11553_, _22167_, _22166_);
  nand _55527_ (_22168_, _20505_, _28096_);
  nand _55528_ (_22169_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nand _55529_ (_11555_, _22169_, _22168_);
  nand _55530_ (_22170_, _07423_, _24830_);
  nand _55531_ (_22171_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  nand _55532_ (_11557_, _22171_, _22170_);
  nand _55533_ (_22172_, _20505_, _24927_);
  nand _55534_ (_22173_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  nand _55535_ (_28345_, _22173_, _22172_);
  nand _55536_ (_22174_, _20726_, _24789_);
  nand _55537_ (_22175_, _20728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  nand _55538_ (_11559_, _22175_, _22174_);
  nand _55539_ (_22176_, _20505_, _25150_);
  nand _55540_ (_22177_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nand _55541_ (_11561_, _22177_, _22176_);
  nand _55542_ (_22178_, _20722_, _24830_);
  nand _55543_ (_22179_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nand _55544_ (_11563_, _22179_, _22178_);
  nand _55545_ (_22180_, _20722_, _28096_);
  nand _55546_ (_22181_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  nand _55547_ (_11567_, _22181_, _22180_);
  nand _55548_ (_22182_, _20505_, _24789_);
  nand _55549_ (_22183_, _20507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  nand _55550_ (_11569_, _22183_, _22182_);
  nand _55551_ (_22184_, _28096_, _28081_);
  nand _55552_ (_22185_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  nand _55553_ (_11574_, _22185_, _22184_);
  nand _55554_ (_22186_, _01116_, _24830_);
  nand _55555_ (_22187_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  nand _55556_ (_11576_, _22187_, _22186_);
  nand _55557_ (_22188_, _28096_, _25061_);
  nand _55558_ (_22189_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  nand _55559_ (_11578_, _22189_, _22188_);
  nand _55560_ (_22190_, _20722_, _25203_);
  nand _55561_ (_22191_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  nand _55562_ (_11580_, _22191_, _22190_);
  nand _55563_ (_22192_, _18135_, _25099_);
  nand _55564_ (_22193_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  nand _55565_ (_11587_, _22193_, _22192_);
  nand _55566_ (_22194_, _18135_, _25203_);
  nand _55567_ (_22195_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  nand _55568_ (_28258_, _22195_, _22194_);
  nand _55569_ (_22196_, _03822_, _25150_);
  nand _55570_ (_22197_, _03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  nand _55571_ (_11592_, _22197_, _22196_);
  nand _55572_ (_22198_, _18135_, _28096_);
  nand _55573_ (_22199_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nand _55574_ (_11593_, _22199_, _22198_);
  nor _55575_ (_22200_, _21113_, _18553_);
  nand _55576_ (_22201_, _22200_, _07983_);
  not _55577_ (_22202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand _55578_ (_22203_, _17053_, _22202_);
  nand _55579_ (_22204_, _22203_, _07975_);
  nand _55580_ (_22205_, _22204_, _17059_);
  nand _55581_ (_22206_, _17060_, _22202_);
  nand _55582_ (_22207_, _22206_, _22205_);
  nand _55583_ (_22208_, _22207_, _22201_);
  nand _55584_ (_22209_, _22208_, _18328_);
  nand _55585_ (_22210_, _18307_, _25194_);
  nand _55586_ (_11598_, _22210_, _22209_);
  nand _55587_ (_22211_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  nand _55588_ (_22212_, _28074_, _25099_);
  nand _55589_ (_11600_, _22212_, _22211_);
  nand _55590_ (_22213_, _18334_, _25039_);
  nand _55591_ (_22214_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  nand _55592_ (_11602_, _22214_, _22213_);
  nand _55593_ (_22215_, _00979_, _25039_);
  nand _55594_ (_22216_, _00981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nand _55595_ (_11603_, _22216_, _22215_);
  nand _55596_ (_22217_, _08653_, _25099_);
  nand _55597_ (_22218_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  nand _55598_ (_11605_, _22218_, _22217_);
  nand _55599_ (_22219_, _01905_, _24830_);
  nand _55600_ (_22220_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand _55601_ (_28315_, _22220_, _22219_);
  nand _55602_ (_22221_, _01905_, _25150_);
  nand _55603_ (_22222_, _01907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nand _55604_ (_11608_, _22222_, _22221_);
  nand _55605_ (_22223_, _28081_, _25150_);
  nand _55606_ (_22224_, _28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nand _55607_ (_11610_, _22224_, _22223_);
  nand _55608_ (_22225_, _08387_, _25099_);
  nand _55609_ (_22226_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nand _55610_ (_11613_, _22226_, _22225_);
  nand _55611_ (_22227_, _18519_, _25039_);
  nand _55612_ (_22228_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nand _55613_ (_11614_, _22228_, _22227_);
  nand _55614_ (_22229_, _25099_, _25000_);
  nand _55615_ (_22230_, _25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  nand _55616_ (_11617_, _22230_, _22229_);
  nand _55617_ (_22231_, _08653_, _24830_);
  nand _55618_ (_22232_, _08655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  nand _55619_ (_11618_, _22232_, _22231_);
  nand _55620_ (_22233_, _08387_, _24830_);
  nand _55621_ (_22234_, _08390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  nand _55622_ (_11620_, _22234_, _22233_);
  nor _55623_ (_22235_, _00271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor _55624_ (_22236_, _00272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _55625_ (_22237_, _22236_, _22235_);
  nor _55626_ (_22238_, _22237_, _00279_);
  nor _55627_ (_22239_, _00287_, _24821_);
  nor _55628_ (_22240_, _22239_, _22238_);
  nor _55629_ (_22241_, _22240_, _03944_);
  nand _55630_ (_22243_, _03944_, _05904_);
  nand _55631_ (_22244_, _22243_, _26487_);
  nor _55632_ (_11622_, _22244_, _22241_);
  nor _55633_ (_22245_, _00287_, _25680_);
  nand _55634_ (_22246_, _00272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand _55635_ (_22247_, _00271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand _55636_ (_22248_, _22247_, _22246_);
  nor _55637_ (_22249_, _22248_, _00279_);
  nor _55638_ (_22250_, _22249_, _22245_);
  nor _55639_ (_22251_, _22250_, _03944_);
  not _55640_ (_22252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand _55641_ (_22253_, _03944_, _22252_);
  nand _55642_ (_22254_, _22253_, _26487_);
  nor _55643_ (_11624_, _22254_, _22251_);
  nor _55644_ (_22255_, _00287_, _25089_);
  nand _55645_ (_22256_, _00272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand _55646_ (_22257_, _00271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _55647_ (_22258_, _22257_, _22256_);
  nor _55648_ (_22259_, _22258_, _00279_);
  nor _55649_ (_22260_, _22259_, _22255_);
  nor _55650_ (_22261_, _22260_, _03944_);
  nand _55651_ (_22262_, _03944_, _12426_);
  nand _55652_ (_22263_, _22262_, _26487_);
  nor _55653_ (_11626_, _22263_, _22261_);
  nor _55654_ (_22264_, _00287_, _24920_);
  nor _55655_ (_22265_, _00271_, _20675_);
  nor _55656_ (_22266_, _00272_, _00173_);
  nor _55657_ (_22267_, _22266_, _22265_);
  nand _55658_ (_22268_, _22267_, _00287_);
  nand _55659_ (_22269_, _22268_, _00269_);
  nor _55660_ (_22270_, _22269_, _22264_);
  nor _55661_ (_22271_, _00297_, _20675_);
  nor _55662_ (_22272_, _22271_, _22270_);
  nor _55663_ (_11630_, _22272_, rst);
  nor _55664_ (_22273_, _00287_, _25028_);
  nand _55665_ (_22274_, _00272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _55666_ (_22275_, _00271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _55667_ (_22276_, _22275_, _22274_);
  nor _55668_ (_22277_, _22276_, _00279_);
  nor _55669_ (_22278_, _22277_, _22273_);
  nor _55670_ (_22279_, _22278_, _03944_);
  not _55671_ (_22280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _55672_ (_22281_, _03944_, _22280_);
  nand _55673_ (_22282_, _22281_, _26487_);
  nor _55674_ (_11632_, _22282_, _22279_);
  nand _55675_ (_22283_, _13080_, _24927_);
  nand _55676_ (_22284_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  nand _55677_ (_11635_, _22284_, _22283_);
  nand _55678_ (_22285_, _00995_, _25203_);
  nand _55679_ (_22286_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  nand _55680_ (_28366_, _22286_, _22285_);
  nand _55681_ (_22287_, _01009_, _25039_);
  nand _55682_ (_22288_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  nand _55683_ (_11641_, _22288_, _22287_);
  nand _55684_ (_22289_, _03911_, _25099_);
  nand _55685_ (_22290_, _03913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  nand _55686_ (_28284_, _22290_, _22289_);
  nand _55687_ (_22291_, _19024_, _28096_);
  nand _55688_ (_22292_, _19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  nand _55689_ (_11645_, _22292_, _22291_);
  nand _55690_ (_22293_, _18334_, _24927_);
  nand _55691_ (_22294_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nand _55692_ (_11650_, _22294_, _22293_);
  nand _55693_ (_22295_, _03540_, _24830_);
  nand _55694_ (_22296_, _03542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nand _55695_ (_11651_, _22296_, _22295_);
  nand _55696_ (_22297_, _01001_, _24830_);
  nand _55697_ (_22298_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  nand _55698_ (_11653_, _22298_, _22297_);
  nand _55699_ (_22299_, _01120_, _24927_);
  nand _55700_ (_22300_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  nand _55701_ (_11655_, _22300_, _22299_);
  nand _55702_ (_22301_, _01120_, _25203_);
  nand _55703_ (_22302_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nand _55704_ (_11656_, _22302_, _22301_);
  nand _55705_ (_22303_, _08806_, _25150_);
  nand _55706_ (_22304_, _08808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  nand _55707_ (_11664_, _22304_, _22303_);
  nand _55708_ (_22305_, _00985_, _24927_);
  nand _55709_ (_22306_, _00987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nand _55710_ (_11667_, _22306_, _22305_);
  nand _55711_ (_22308_, _01001_, _25099_);
  nand _55712_ (_22309_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  nand _55713_ (_28348_, _22309_, _22308_);
  nand _55714_ (_22310_, _01120_, _25039_);
  nand _55715_ (_22311_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nand _55716_ (_11689_, _22311_, _22310_);
  nand _55717_ (_22312_, _01009_, _24830_);
  nand _55718_ (_22313_, _01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nand _55719_ (_11691_, _22313_, _22312_);
  nand _55720_ (_22314_, _08344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nand _55721_ (_22315_, _08343_, _25150_);
  nand _55722_ (_11704_, _22315_, _22314_);
  nand _55723_ (_22316_, _01104_, _25099_);
  nand _55724_ (_22317_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nand _55725_ (_11707_, _22317_, _22316_);
  nand _55726_ (_22318_, _28099_, _25150_);
  nand _55727_ (_22319_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  nand _55728_ (_11709_, _22319_, _22318_);
  nand _55729_ (_22320_, _01108_, _25203_);
  nand _55730_ (_22321_, _01110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  nand _55731_ (_11710_, _22321_, _22320_);
  nand _55732_ (_22322_, _01140_, _25150_);
  nand _55733_ (_22323_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nand _55734_ (_11712_, _22323_, _22322_);
  nand _55735_ (_22324_, _08551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  nand _55736_ (_22325_, _08549_, _24830_);
  nand _55737_ (_11714_, _22325_, _22324_);
  nand _55738_ (_22326_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  nand _55739_ (_22327_, _08334_, _24789_);
  nand _55740_ (_11715_, _22327_, _22326_);
  nand _55741_ (_22328_, _01001_, _25039_);
  nand _55742_ (_22329_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nand _55743_ (_11717_, _22329_, _22328_);
  nand _55744_ (_22330_, _01001_, _25150_);
  nand _55745_ (_22331_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  nand _55746_ (_11719_, _22331_, _22330_);
  nand _55747_ (_22332_, _18135_, _24927_);
  nand _55748_ (_22333_, _18137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  nand _55749_ (_28259_, _22333_, _22332_);
  nand _55750_ (_22335_, _07810_, _25203_);
  nand _55751_ (_22336_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nand _55752_ (_11721_, _22336_, _22335_);
  nand _55753_ (_22337_, _00995_, _25099_);
  nand _55754_ (_22338_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  nand _55755_ (_11723_, _22338_, _22337_);
  nand _55756_ (_22339_, _01120_, _25150_);
  nand _55757_ (_22340_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  nand _55758_ (_11725_, _22340_, _22339_);
  nand _55759_ (_22341_, _01120_, _24789_);
  nand _55760_ (_22342_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nand _55761_ (_11727_, _22342_, _22341_);
  nand _55762_ (_22343_, _18334_, _24830_);
  nand _55763_ (_22344_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nand _55764_ (_11728_, _22344_, _22343_);
  nand _55765_ (_22345_, _01001_, _25203_);
  nand _55766_ (_22346_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nand _55767_ (_11730_, _22346_, _22345_);
  nand _55768_ (_22347_, _01140_, _28096_);
  nand _55769_ (_22348_, _01142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nand _55770_ (_11732_, _22348_, _22347_);
  nor _55771_ (_11733_, _02581_, rst);
  nor _55772_ (_11735_, _02638_, rst);
  nor _55773_ (_11737_, _02707_, rst);
  nand _55774_ (_22349_, _00995_, _24830_);
  nand _55775_ (_22350_, _00997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  nand _55776_ (_11740_, _22350_, _22349_);
  nand _55777_ (_22351_, _01001_, _24927_);
  nand _55778_ (_22352_, _01003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  nand _55779_ (_11743_, _22352_, _22351_);
  nor _55780_ (_11752_, _02841_, rst);
  nor _55781_ (_22353_, _24770_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  nand _55782_ (_22354_, _24770_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  nand _55783_ (_22355_, _22354_, _26487_);
  nor _55784_ (_11754_, _22355_, _22353_);
  nor _55785_ (_11757_, _01953_, rst);
  nor _55786_ (_11760_, _02067_, rst);
  nor _55787_ (_11763_, _20428_, rst);
  not _55788_ (_22356_, _02269_);
  nor _55789_ (_11766_, _22356_, rst);
  nand _55790_ (_22357_, _01104_, _24927_);
  nand _55791_ (_22358_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  nand _55792_ (_11768_, _22358_, _22357_);
  nand _55793_ (_22359_, _19068_, _24830_);
  nand _55794_ (_22360_, _19070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  nand _55795_ (_28368_, _22360_, _22359_);
  nand _55796_ (_22361_, _01104_, _24789_);
  nand _55797_ (_22362_, _01106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  nand _55798_ (_28367_, _22362_, _22361_);
  nand _55799_ (_22363_, _01208_, _25099_);
  nand _55800_ (_22364_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nand _55801_ (_11773_, _22364_, _22363_);
  nand _55802_ (_22365_, _01533_, _25150_);
  nand _55803_ (_22366_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nand _55804_ (_11775_, _22366_, _22365_);
  nand _55805_ (_22367_, _01533_, _24830_);
  nand _55806_ (_22368_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  nand _55807_ (_11777_, _22368_, _22367_);
  nand _55808_ (_22369_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  nand _55809_ (_22370_, _08339_, _25150_);
  nand _55810_ (_11779_, _22370_, _22369_);
  nand _55811_ (_22371_, _19119_, _24830_);
  nand _55812_ (_22372_, _19121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  nand _55813_ (_11780_, _22372_, _22371_);
  nand _55814_ (_22373_, _01116_, _25203_);
  nand _55815_ (_22374_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  nand _55816_ (_28346_, _22374_, _22373_);
  nand _55817_ (_22375_, _06437_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor _55818_ (_22376_, _25509_, _25563_);
  nand _55819_ (_22377_, _06605_, _06488_);
  nor _55820_ (_22378_, _22377_, _22376_);
  nor _55821_ (_22379_, _25574_, _25532_);
  nor _55822_ (_22380_, _06613_, _25584_);
  nand _55823_ (_22381_, _22380_, _22379_);
  nand _55824_ (_22382_, _01061_, _25411_);
  nor _55825_ (_22383_, _01050_, _25467_);
  nand _55826_ (_22384_, _22383_, _22382_);
  nor _55827_ (_22385_, _22384_, _22381_);
  nand _55828_ (_22386_, _22385_, _22378_);
  nand _55829_ (_22387_, _22386_, _00883_);
  nand _55830_ (_28192_[1], _22387_, _22375_);
  not _55831_ (_22388_, _02000_);
  nor _55832_ (_11799_, _22388_, rst);
  nor _55833_ (_11801_, _27511_, rst);
  nor _55834_ (_11803_, _02782_, rst);
  nand _55835_ (_22389_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  nand _55836_ (_22390_, _08339_, _24789_);
  nand _55837_ (_11804_, _22390_, _22389_);
  nor _55838_ (_11806_, _27272_, rst);
  nand _55839_ (_22391_, _01116_, _24927_);
  nand _55840_ (_22392_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  nand _55841_ (_11808_, _22392_, _22391_);
  nand _55842_ (_22393_, _18523_, _25039_);
  nand _55843_ (_22394_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  nand _55844_ (_11810_, _22394_, _22393_);
  nand _55845_ (_22395_, _18334_, _28096_);
  nand _55846_ (_22396_, _18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  nand _55847_ (_11812_, _22396_, _22395_);
  nand _55848_ (_22397_, _18523_, _25203_);
  nand _55849_ (_22398_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nand _55850_ (_11814_, _22398_, _22397_);
  nand _55851_ (_22399_, _01120_, _24830_);
  nand _55852_ (_22400_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  nand _55853_ (_11817_, _22400_, _22399_);
  nand _55854_ (_22401_, _01120_, _25099_);
  nand _55855_ (_22402_, _01123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  nand _55856_ (_11819_, _22402_, _22401_);
  nand _55857_ (_22403_, _01116_, _25150_);
  nand _55858_ (_22404_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nand _55859_ (_11821_, _22404_, _22403_);
  nand _55860_ (_22405_, _28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nand _55861_ (_22406_, _28074_, _24830_);
  nand _55862_ (_11823_, _22406_, _22405_);
  nand _55863_ (_22407_, _18523_, _28096_);
  nand _55864_ (_22408_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nand _55865_ (_11825_, _22408_, _22407_);
  nand _55866_ (_22409_, _06437_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _55867_ (_22410_, _18736_);
  nand _55868_ (_22411_, _01064_, _25428_);
  nand _55869_ (_22412_, _06524_, _04277_);
  nor _55870_ (_22414_, _22412_, _22411_);
  nand _55871_ (_22415_, _22414_, _22410_);
  nand _55872_ (_22416_, _22415_, _00883_);
  nand _55873_ (_28189_[1], _22416_, _22409_);
  nand _55874_ (_22417_, _01533_, _25203_);
  nand _55875_ (_22418_, _01535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  nand _55876_ (_11830_, _22418_, _22417_);
  nand _55877_ (_22419_, _28099_, _24789_);
  nand _55878_ (_22420_, _28101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  nand _55879_ (_11832_, _22420_, _22419_);
  nand _55880_ (_22421_, _20722_, _25150_);
  nand _55881_ (_22422_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nand _55882_ (_11833_, _22422_, _22421_);
  nand _55883_ (_22423_, _20170_, _24830_);
  nand _55884_ (_22424_, _20172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  nand _55885_ (_11838_, _22424_, _22423_);
  nand _55886_ (_22425_, _01116_, _28096_);
  nand _55887_ (_22426_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nand _55888_ (_11847_, _22426_, _22425_);
  nand _55889_ (_22427_, _25150_, _25061_);
  nand _55890_ (_22428_, _25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  nand _55891_ (_28334_, _22428_, _22427_);
  nand _55892_ (_22429_, _18519_, _24789_);
  nand _55893_ (_22430_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  nand _55894_ (_11851_, _22430_, _22429_);
  nand _55895_ (_22431_, _01116_, _25039_);
  nand _55896_ (_22432_, _01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  nand _55897_ (_28347_, _22432_, _22431_);
  nand _55898_ (_22433_, _20722_, _24789_);
  nand _55899_ (_22434_, _20724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  nand _55900_ (_11860_, _22434_, _22433_);
  nand _55901_ (_22435_, _03850_, _24830_);
  nand _55902_ (_22436_, _03852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nand _55903_ (_11866_, _22436_, _22435_);
  nand _55904_ (_22437_, _18523_, _25150_);
  nand _55905_ (_22438_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  nand _55906_ (_11878_, _22438_, _22437_);
  nand _55907_ (_22439_, _01208_, _25039_);
  nand _55908_ (_22440_, _01210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  nand _55909_ (_11881_, _22440_, _22439_);
  nand _55910_ (_22441_, _13080_, _25150_);
  nand _55911_ (_22442_, _13082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nand _55912_ (_11883_, _22442_, _22441_);
  nand _55913_ (_22443_, _18519_, _25150_);
  nand _55914_ (_22444_, _18521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  nand _55915_ (_11885_, _22444_, _22443_);
  nor _55916_ (_22445_, _24770_, _27099_);
  nor _55917_ (_22446_, _27104_, _27506_);
  nor _55918_ (_22447_, _22446_, _22445_);
  nor _55919_ (_11888_, _22447_, rst);
  nand _55920_ (_22448_, _00479_, _25099_);
  nand _55921_ (_22449_, _00481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nand _55922_ (_11890_, _22449_, _22448_);
  nor _55923_ (_11893_, _02529_, rst);
  not _55924_ (_22450_, _02132_);
  nor _55925_ (_11897_, _22450_, rst);
  nand _55926_ (_22451_, _18523_, _24789_);
  nand _55927_ (_22452_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  nand _55928_ (_11965_, _22452_, _22451_);
  nand _55929_ (_22453_, _24866_, first_instr);
  nand _55930_ (_00000_, _22453_, _26487_);
  nand _55931_ (_22454_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nand _55932_ (_22455_, _08334_, _28096_);
  nand _55933_ (_11970_, _22455_, _22454_);
  nor _55934_ (_22456_, _00059_, _00055_);
  nand _55935_ (_22457_, _22456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _55936_ (_22458_, _22457_, _00067_);
  not _55937_ (_22459_, _22458_);
  nor _55938_ (_22460_, _00051_, _00047_);
  not _55939_ (_22461_, _22460_);
  nor _55940_ (_22463_, _22461_, _00043_);
  not _55941_ (_22464_, _22463_);
  nor _55942_ (_22465_, _22464_, _22459_);
  not _55943_ (_22466_, _22465_);
  nor _55944_ (_22467_, _22466_, _00071_);
  not _55945_ (_22468_, _22467_);
  nor _55946_ (_22469_, _22468_, _00075_);
  nand _55947_ (_22470_, _22469_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _55948_ (_22471_, _22470_, _00083_);
  not _55949_ (_22472_, _22471_);
  nor _55950_ (_22473_, _22472_, _00087_);
  nand _55951_ (_22474_, _22473_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _55952_ (_22475_, _22474_, _00095_);
  nor _55953_ (_22476_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _55954_ (_22477_, _24873_, _24868_);
  nor _55955_ (_22478_, _22477_, _22476_);
  not _55956_ (_22479_, _22474_);
  nor _55957_ (_22480_, _22479_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _55958_ (_22481_, _22480_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _55959_ (_22482_, _22481_, _22478_);
  nor _55960_ (_22483_, _22482_, _22475_);
  nor _55961_ (_22484_, _00075_, _00071_);
  not _55962_ (_22485_, _22484_);
  nor _55963_ (_22486_, _22485_, _00079_);
  not _55964_ (_22487_, _22486_);
  nor _55965_ (_22488_, _22487_, _22466_);
  not _55966_ (_22489_, _22488_);
  nor _55967_ (_22490_, _22489_, _00083_);
  not _55968_ (_22491_, _22490_);
  nor _55969_ (_22492_, _22491_, _00087_);
  not _55970_ (_22493_, _22492_);
  nand _55971_ (_22494_, _22493_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nand _55972_ (_22495_, _22492_, _00091_);
  nand _55973_ (_22496_, _22495_, _22494_);
  nor _55974_ (_22497_, _22496_, _00031_);
  nand _55975_ (_22498_, _22496_, _00031_);
  not _55976_ (_22499_, _22478_);
  nand _55977_ (_22500_, _22499_, _22475_);
  nand _55978_ (_22501_, _22500_, _22498_);
  nor _55979_ (_22502_, _22501_, _22497_);
  nor _55980_ (_22503_, _22480_, _22475_);
  nor _55981_ (_22504_, _22503_, _00035_);
  nor _55982_ (_22505_, _22490_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _55983_ (_22506_, _22505_, _22492_);
  not _55984_ (_22507_, _22506_);
  nor _55985_ (_22508_, _22507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _55986_ (_22509_, _22506_, _00027_);
  nor _55987_ (_22510_, _22509_, _22508_);
  nor _55988_ (_22511_, _22464_, _00055_);
  nand _55989_ (_22512_, _00059_, _28131_);
  nand _55990_ (_22513_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _55991_ (_22514_, _22513_, _22512_);
  nor _55992_ (_22515_, _22514_, _22511_);
  nand _55993_ (_22516_, _22514_, _22511_);
  nor _55994_ (_22517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _55995_ (_22518_, _00055_, _28127_);
  nor _55996_ (_22519_, _22518_, _22517_);
  nor _55997_ (_22520_, _22519_, _22464_);
  nor _55998_ (_22521_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _28110_);
  nor _55999_ (_22522_, _00039_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _56000_ (_22523_, _22522_, _22521_);
  nand _56001_ (_22524_, _00043_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _56002_ (_22525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _28115_);
  nand _56003_ (_22526_, _22525_, _22524_);
  nand _56004_ (_22527_, _22526_, _22523_);
  nor _56005_ (_22528_, _22527_, _22520_);
  nand _56006_ (_22529_, _22528_, _22516_);
  nor _56007_ (_22530_, _22529_, _22515_);
  nor _56008_ (_22531_, _00047_, _00043_);
  not _56009_ (_22532_, _22531_);
  nor _56010_ (_22533_, _22532_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56011_ (_22534_, _22531_, _00051_);
  nor _56012_ (_22535_, _22534_, _22533_);
  not _56013_ (_22536_, _22535_);
  nor _56014_ (_22537_, _22536_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56015_ (_22538_, _22535_, _28123_);
  nor _56016_ (_22539_, _22538_, _22537_);
  nor _56017_ (_22540_, _00047_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _56018_ (_22541_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _00043_);
  nor _56019_ (_22542_, _22541_, _22540_);
  nand _56020_ (_22543_, _22542_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _56021_ (_22544_, _22542_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _56022_ (_22545_, _22519_);
  nor _56023_ (_22546_, _22545_, _22463_);
  nor _56024_ (_22547_, _22546_, _22544_);
  nand _56025_ (_22548_, _22547_, _22543_);
  nor _56026_ (_22549_, _22548_, _22539_);
  nand _56027_ (_22550_, _22549_, _22530_);
  nor _56028_ (_22551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _56029_ (_22552_, _00075_, _00014_);
  nor _56030_ (_22553_, _22552_, _22551_);
  nor _56031_ (_22554_, _22553_, _22468_);
  not _56032_ (_22555_, _22553_);
  nor _56033_ (_22556_, _22555_, _22467_);
  nor _56034_ (_22557_, _22556_, _22554_);
  nand _56035_ (_22558_, _22463_, _22456_);
  nor _56036_ (_22559_, _22558_, _00063_);
  not _56037_ (_22560_, _22559_);
  nor _56038_ (_22561_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _56039_ (_22562_, _00067_, _00006_);
  nor _56040_ (_22563_, _22562_, _22561_);
  nor _56041_ (_22564_, _22563_, _22560_);
  not _56042_ (_22565_, _22563_);
  nor _56043_ (_22566_, _22565_, _22559_);
  nor _56044_ (_22567_, _22566_, _22564_);
  nand _56045_ (_22568_, _22567_, _22557_);
  nor _56046_ (_22569_, _22568_, _22550_);
  nor _56047_ (_22570_, _22465_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _56048_ (_22571_, _22570_, _22467_);
  not _56049_ (_22572_, _22571_);
  nor _56050_ (_22573_, _22572_, _00010_);
  nor _56051_ (_22574_, _22571_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _56052_ (_22575_, _22574_, _22573_);
  not _56053_ (_22576_, _22558_);
  nor _56054_ (_22577_, _22576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _56055_ (_22578_, _22577_, _22559_);
  not _56056_ (_22579_, _22578_);
  nor _56057_ (_22580_, _22579_, _00001_);
  nor _56058_ (_22581_, _22578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _56059_ (_22582_, _22581_, _22580_);
  nor _56060_ (_22583_, _22582_, _22575_);
  nand _56061_ (_22584_, _22583_, _22569_);
  nor _56062_ (_22585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _56063_ (_22586_, _00083_, _00023_);
  nor _56064_ (_22587_, _22586_, _22585_);
  nor _56065_ (_22588_, _22587_, _22489_);
  not _56066_ (_22589_, _22587_);
  nor _56067_ (_22590_, _22589_, _22488_);
  nor _56068_ (_22591_, _22590_, _22588_);
  nor _56069_ (_22592_, _22469_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _56070_ (_22594_, _22592_, _22488_);
  not _56071_ (_22595_, _22594_);
  nor _56072_ (_22596_, _22595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _56073_ (_22597_, _22594_, _00018_);
  nor _56074_ (_22598_, _22597_, _22596_);
  nand _56075_ (_22599_, _22598_, _22591_);
  nor _56076_ (_22600_, _22599_, _22584_);
  nand _56077_ (_22601_, _22600_, _22510_);
  nor _56078_ (_22602_, _22601_, _22504_);
  nand _56079_ (_22603_, _22602_, _22502_);
  nor _56080_ (_22604_, _22603_, _22483_);
  nor _56081_ (_22605_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56082_ (_22606_, \oc8051_symbolic_cxrom1.regvalid [14], _00051_);
  nor _56083_ (_22607_, _22606_, _00047_);
  not _56084_ (_22608_, _22607_);
  nor _56085_ (_22609_, _22608_, _22605_);
  nor _56086_ (_22610_, _06935_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56087_ (_22611_, _06932_, _00051_);
  nor _56088_ (_22612_, _22611_, _22610_);
  nor _56089_ (_22613_, _22612_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56090_ (_22614_, _22613_, _22609_);
  nor _56091_ (_22615_, _22614_, _00043_);
  nor _56092_ (_22616_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56093_ (_22617_, \oc8051_symbolic_cxrom1.regvalid [8], _00051_);
  nor _56094_ (_22618_, _22617_, _22616_);
  nand _56095_ (_22619_, _22618_, _00047_);
  nor _56096_ (_22620_, \oc8051_symbolic_cxrom1.regvalid [12], _00051_);
  nor _56097_ (_22621_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56098_ (_22622_, _22621_, _22620_);
  nand _56099_ (_22623_, _22622_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nand _56100_ (_22624_, _22623_, _22619_);
  nand _56101_ (_22625_, _22624_, _00043_);
  not _56102_ (_22626_, _22625_);
  nor _56103_ (_22627_, _22626_, _22615_);
  nand _56104_ (_22628_, _22627_, _00039_);
  nor _56105_ (_22629_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56106_ (_22630_, \oc8051_symbolic_cxrom1.regvalid [15], _00051_);
  nor _56107_ (_22631_, _22630_, _00047_);
  not _56108_ (_22632_, _22631_);
  nor _56109_ (_22633_, _22632_, _22629_);
  nor _56110_ (_22634_, _06852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56111_ (_22635_, _06871_, _00051_);
  nor _56112_ (_22636_, _22635_, _22634_);
  nor _56113_ (_22637_, _22636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56114_ (_22638_, _22637_, _22633_);
  nor _56115_ (_22639_, _22638_, _00043_);
  nor _56116_ (_22640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _56117_ (_22641_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56118_ (_22642_, \oc8051_symbolic_cxrom1.regvalid [9], _00051_);
  nor _56119_ (_22643_, _22642_, _22641_);
  nand _56120_ (_22644_, _22643_, _22640_);
  nor _56121_ (_22645_, \oc8051_symbolic_cxrom1.regvalid [13], _00051_);
  nor _56122_ (_22646_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56123_ (_22647_, _22646_, _22645_);
  nand _56124_ (_22648_, _22647_, _22540_);
  nand _56125_ (_22649_, _22648_, _22644_);
  nor _56126_ (_22650_, _22649_, _22639_);
  nand _56127_ (_22651_, _22650_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand _56128_ (_22652_, _22651_, _22628_);
  nor _56129_ (_22653_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _00039_);
  nand _56130_ (_22654_, _22653_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  not _56131_ (_22655_, _22654_);
  nor _56132_ (_22656_, _22655_, _00047_);
  nor _56133_ (_22657_, _00043_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _56134_ (_22658_, _22657_);
  nor _56135_ (_22659_, _22658_, _09052_);
  nor _56136_ (_22660_, _00043_, _00039_);
  nand _56137_ (_22661_, _22660_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nor _56138_ (_22662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand _56139_ (_22663_, _22662_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _56140_ (_22664_, _22663_, _22661_);
  nor _56141_ (_22665_, _22664_, _22659_);
  nand _56142_ (_22666_, _22665_, _22656_);
  nand _56143_ (_22667_, _22657_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  not _56144_ (_22668_, _22667_);
  not _56145_ (_22669_, _22660_);
  nor _56146_ (_22670_, _22669_, _08635_);
  nor _56147_ (_22671_, _22670_, _22668_);
  not _56148_ (_22672_, _22653_);
  nor _56149_ (_22673_, _22672_, _08304_);
  not _56150_ (_22675_, _22662_);
  nor _56151_ (_22676_, _22675_, _08129_);
  nor _56152_ (_22677_, _22676_, _22673_);
  nand _56153_ (_22678_, _22677_, _22671_);
  nor _56154_ (_22679_, _22678_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56155_ (_22680_, _22679_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand _56156_ (_22681_, _22680_, _22666_);
  nor _56157_ (_22682_, _00051_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  not _56158_ (_22683_, _22682_);
  nand _56159_ (_22684_, _22660_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _56160_ (_22685_, _22662_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _56161_ (_22686_, _22685_, _22684_);
  nand _56162_ (_22687_, _22657_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _56163_ (_22688_, _22653_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _56164_ (_22689_, _22688_, _22687_);
  nor _56165_ (_22690_, _22689_, _22686_);
  nor _56166_ (_22691_, _22690_, _22683_);
  nor _56167_ (_22692_, _22669_, _07372_);
  nor _56168_ (_22693_, _22675_, _09788_);
  nor _56169_ (_22694_, _22693_, _22692_);
  not _56170_ (_22696_, _22694_);
  nand _56171_ (_22697_, _22657_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _56172_ (_22698_, _22653_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _56173_ (_22699_, _22698_, _22697_);
  nor _56174_ (_22700_, _22699_, _22696_);
  nor _56175_ (_22701_, _22700_, _22461_);
  nor _56176_ (_22702_, _22701_, _22691_);
  nand _56177_ (_22703_, _22702_, _22681_);
  not _56178_ (_22704_, _22703_);
  nor _56179_ (_22705_, _22704_, _22652_);
  not _56180_ (_22706_, _22705_);
  not _56181_ (_22707_, _22652_);
  nand _56182_ (_22708_, _22657_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nand _56183_ (_22709_, _22660_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nand _56184_ (_22710_, _22709_, _22708_);
  nand _56185_ (_22711_, _22653_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  not _56186_ (_22712_, _22711_);
  nor _56187_ (_22713_, _22675_, _08781_);
  nor _56188_ (_22714_, _22713_, _22712_);
  not _56189_ (_22715_, _22714_);
  nor _56190_ (_22716_, _22715_, _22710_);
  nand _56191_ (_22717_, _22716_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56192_ (_22718_, _22658_, _08459_);
  nor _56193_ (_22719_, _22669_, _08620_);
  nor _56194_ (_22720_, _22719_, _22718_);
  nor _56195_ (_22721_, _22672_, _08285_);
  nand _56196_ (_22722_, _22662_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  not _56197_ (_22723_, _22722_);
  nor _56198_ (_22724_, _22723_, _22721_);
  nand _56199_ (_22725_, _22724_, _22720_);
  nor _56200_ (_22726_, _22725_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56201_ (_22727_, _22726_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand _56202_ (_22728_, _22727_, _22717_);
  nor _56203_ (_22729_, _22669_, _09644_);
  not _56204_ (_22730_, _22729_);
  nand _56205_ (_22731_, _22657_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nand _56206_ (_22732_, _22731_, _22730_);
  nand _56207_ (_22733_, _22662_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nand _56208_ (_22734_, _22653_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nand _56209_ (_22735_, _22734_, _22733_);
  nor _56210_ (_22736_, _22735_, _22732_);
  nor _56211_ (_22737_, _22736_, _22683_);
  nand _56212_ (_22738_, _22660_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nand _56213_ (_22739_, _22662_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nand _56214_ (_22740_, _22739_, _22738_);
  nand _56215_ (_22741_, _22657_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nand _56216_ (_22742_, _22653_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nand _56217_ (_22743_, _22742_, _22741_);
  nor _56218_ (_22744_, _22743_, _22740_);
  nor _56219_ (_22745_, _22744_, _22461_);
  nor _56220_ (_22746_, _22745_, _22737_);
  nand _56221_ (_22747_, _22746_, _22728_);
  nand _56222_ (_22748_, _22747_, _22707_);
  nor _56223_ (_22749_, _22658_, _09008_);
  nor _56224_ (_22750_, _22669_, _10481_);
  nor _56225_ (_22751_, _22750_, _22749_);
  nor _56226_ (_22752_, _22672_, _08878_);
  nor _56227_ (_22753_, _22675_, _10477_);
  nor _56228_ (_22754_, _22753_, _22752_);
  nand _56229_ (_22755_, _22754_, _22751_);
  nor _56230_ (_22756_, _22755_, _00047_);
  nor _56231_ (_22757_, _22675_, _08086_);
  nor _56232_ (_22758_, _22757_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nand _56233_ (_22759_, _22660_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  not _56234_ (_22760_, _22759_);
  nand _56235_ (_22761_, _22657_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nand _56236_ (_22762_, _22653_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand _56237_ (_22763_, _22762_, _22761_);
  nor _56238_ (_22764_, _22763_, _22760_);
  nand _56239_ (_22765_, _22764_, _22758_);
  nand _56240_ (_22766_, _22765_, _00051_);
  nor _56241_ (_22767_, _22766_, _22756_);
  nor _56242_ (_22768_, _22669_, _10491_);
  nor _56243_ (_22769_, _22675_, _10500_);
  nor _56244_ (_22770_, _22769_, _22768_);
  nor _56245_ (_22771_, _22658_, _10493_);
  nor _56246_ (_22772_, _22672_, _10498_);
  nor _56247_ (_22773_, _22772_, _22771_);
  nand _56248_ (_22774_, _22773_, _22770_);
  nand _56249_ (_22775_, _22774_, _22682_);
  nor _56250_ (_22776_, _22669_, _10516_);
  nor _56251_ (_22777_, _22675_, _10509_);
  nor _56252_ (_22778_, _22777_, _22776_);
  nor _56253_ (_22779_, _22658_, _10518_);
  nor _56254_ (_22780_, _22672_, _10507_);
  nor _56255_ (_22781_, _22780_, _22779_);
  nand _56256_ (_22782_, _22781_, _22778_);
  nand _56257_ (_22783_, _22782_, _22460_);
  nand _56258_ (_22784_, _22783_, _22775_);
  nor _56259_ (_22785_, _22784_, _22767_);
  not _56260_ (_22787_, _22785_);
  nor _56261_ (_22788_, _22658_, _08996_);
  nand _56262_ (_22789_, _22660_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  not _56263_ (_22790_, _22789_);
  nor _56264_ (_22791_, _22790_, _22788_);
  nor _56265_ (_22792_, _22672_, _08864_);
  nor _56266_ (_22793_, _22675_, _08739_);
  nor _56267_ (_22794_, _22793_, _22792_);
  nand _56268_ (_22795_, _22794_, _22791_);
  nor _56269_ (_22796_, _22795_, _00047_);
  nor _56270_ (_22797_, _22658_, _08419_);
  nor _56271_ (_22798_, _22669_, _10442_);
  nor _56272_ (_22799_, _22798_, _22797_);
  nor _56273_ (_22800_, _22672_, _08237_);
  nor _56274_ (_22801_, _22675_, _10438_);
  nor _56275_ (_22802_, _22801_, _22800_);
  nand _56276_ (_22803_, _22802_, _22799_);
  nor _56277_ (_22804_, _22803_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56278_ (_22805_, _22804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _56279_ (_22806_, _22805_);
  nor _56280_ (_22807_, _22806_, _22796_);
  nand _56281_ (_22808_, _22660_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nand _56282_ (_22809_, _22657_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nand _56283_ (_22810_, _22809_, _22808_);
  nand _56284_ (_22811_, _22662_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _56285_ (_22812_, _22672_, _09365_);
  not _56286_ (_22813_, _22812_);
  nand _56287_ (_22814_, _22813_, _22811_);
  nor _56288_ (_22815_, _22814_, _22810_);
  nor _56289_ (_22816_, _22815_, _22683_);
  nor _56290_ (_22817_, _22669_, _10431_);
  nand _56291_ (_22818_, _22662_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  not _56292_ (_22819_, _22818_);
  nor _56293_ (_22820_, _22819_, _22817_);
  nor _56294_ (_22821_, _22658_, _10433_);
  nand _56295_ (_22822_, _22653_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  not _56296_ (_22823_, _22822_);
  nor _56297_ (_22824_, _22823_, _22821_);
  nand _56298_ (_22825_, _22824_, _22820_);
  nand _56299_ (_22826_, _22825_, _22460_);
  not _56300_ (_22827_, _22826_);
  nor _56301_ (_22828_, _22827_, _22816_);
  not _56302_ (_22829_, _22828_);
  nor _56303_ (_22830_, _22829_, _22807_);
  nor _56304_ (_22831_, _22830_, _22652_);
  nand _56305_ (_22832_, _22653_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  not _56306_ (_22833_, _22832_);
  nor _56307_ (_22834_, _22833_, _00047_);
  nor _56308_ (_22835_, _22658_, _08983_);
  nand _56309_ (_22836_, _22660_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand _56310_ (_22837_, _22662_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand _56311_ (_22838_, _22837_, _22836_);
  nor _56312_ (_22839_, _22838_, _22835_);
  nand _56313_ (_22840_, _22839_, _22834_);
  nor _56314_ (_22841_, _22658_, _08407_);
  nor _56315_ (_22842_, _22669_, _10384_);
  nor _56316_ (_22843_, _22842_, _22841_);
  nor _56317_ (_22844_, _22672_, _08216_);
  nor _56318_ (_22845_, _22675_, _08056_);
  nor _56319_ (_22846_, _22845_, _22844_);
  nand _56320_ (_22847_, _22846_, _22843_);
  nor _56321_ (_22848_, _22847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56322_ (_22849_, _22848_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand _56323_ (_22850_, _22849_, _22840_);
  nand _56324_ (_22851_, _22660_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nand _56325_ (_22852_, _22662_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nand _56326_ (_22853_, _22852_, _22851_);
  nand _56327_ (_22854_, _22657_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand _56328_ (_22855_, _22653_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand _56329_ (_22856_, _22855_, _22854_);
  nor _56330_ (_22857_, _22856_, _22853_);
  nor _56331_ (_22858_, _22857_, _22683_);
  nor _56332_ (_22859_, _22669_, _10372_);
  nand _56333_ (_22860_, _22662_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  not _56334_ (_22861_, _22860_);
  nor _56335_ (_22862_, _22861_, _22859_);
  nor _56336_ (_22863_, _22658_, _10375_);
  nand _56337_ (_22864_, _22653_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  not _56338_ (_22865_, _22864_);
  nor _56339_ (_22866_, _22865_, _22863_);
  nand _56340_ (_22867_, _22866_, _22862_);
  nand _56341_ (_22868_, _22867_, _22460_);
  not _56342_ (_22869_, _22868_);
  nor _56343_ (_22870_, _22869_, _22858_);
  nand _56344_ (_22871_, _22870_, _22850_);
  nand _56345_ (_22872_, _22871_, _22707_);
  nand _56346_ (_22873_, _22660_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nand _56347_ (_22874_, _22662_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nand _56348_ (_22875_, _22874_, _22873_);
  nand _56349_ (_22876_, _22657_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand _56350_ (_22877_, _22653_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nand _56351_ (_22878_, _22877_, _22876_);
  nor _56352_ (_22879_, _22878_, _22875_);
  nor _56353_ (_22880_, _22879_, _22683_);
  nor _56354_ (_22881_, _22658_, _08964_);
  nand _56355_ (_22882_, _22660_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  not _56356_ (_22883_, _22882_);
  nor _56357_ (_22884_, _22883_, _22881_);
  nor _56358_ (_22885_, _22672_, _08837_);
  nand _56359_ (_22886_, _22662_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  not _56360_ (_22887_, _22886_);
  nor _56361_ (_22888_, _22887_, _22885_);
  nand _56362_ (_22889_, _22888_, _22884_);
  nor _56363_ (_22890_, _22889_, _00047_);
  nor _56364_ (_22891_, _22658_, _08393_);
  nor _56365_ (_22892_, _22669_, _08533_);
  nor _56366_ (_22893_, _22892_, _22891_);
  nor _56367_ (_22894_, _22672_, _08198_);
  nor _56368_ (_22895_, _22675_, _08040_);
  nor _56369_ (_22896_, _22895_, _22894_);
  nand _56370_ (_22897_, _22896_, _22893_);
  nor _56371_ (_22898_, _22897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56372_ (_22899_, _22898_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _56373_ (_22900_, _22899_);
  nor _56374_ (_22901_, _22900_, _22890_);
  not _56375_ (_22902_, _22901_);
  nor _56376_ (_22903_, _22669_, _10313_);
  nand _56377_ (_22904_, _22662_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  not _56378_ (_22905_, _22904_);
  nor _56379_ (_22906_, _22905_, _22903_);
  nor _56380_ (_22907_, _22658_, _10315_);
  nand _56381_ (_22908_, _22653_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  not _56382_ (_22909_, _22908_);
  nor _56383_ (_22910_, _22909_, _22907_);
  nand _56384_ (_22911_, _22910_, _22906_);
  nand _56385_ (_22912_, _22911_, _22460_);
  nand _56386_ (_22913_, _22912_, _22902_);
  nor _56387_ (_22914_, _22913_, _22880_);
  nor _56388_ (_22915_, _22914_, _22872_);
  nor _56389_ (_22916_, _22915_, _22831_);
  nor _56390_ (_22917_, _22916_, _22787_);
  not _56391_ (_22918_, _22917_);
  nand _56392_ (_22919_, _22918_, _22748_);
  nor _56393_ (_22920_, _22914_, _22652_);
  nor _56394_ (_22921_, _22920_, _22872_);
  not _56395_ (_22922_, _22921_);
  nor _56396_ (_22923_, _22922_, _22831_);
  nor _56397_ (_22924_, _22785_, _22652_);
  not _56398_ (_22925_, _22924_);
  nor _56399_ (_22926_, _22658_, _09027_);
  nand _56400_ (_22927_, _22660_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  not _56401_ (_22928_, _22927_);
  nor _56402_ (_22929_, _22928_, _22926_);
  nand _56403_ (_22930_, _22653_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  not _56404_ (_22931_, _22930_);
  nor _56405_ (_22932_, _22675_, _08769_);
  nor _56406_ (_22933_, _22932_, _22931_);
  nand _56407_ (_22934_, _22933_, _22929_);
  nor _56408_ (_22935_, _22934_, _00047_);
  nor _56409_ (_22936_, _22658_, _08447_);
  nor _56410_ (_22937_, _22669_, _08604_);
  nor _56411_ (_22938_, _22937_, _22936_);
  nor _56412_ (_22939_, _22672_, _08269_);
  nor _56413_ (_22940_, _22675_, _08104_);
  nor _56414_ (_22941_, _22940_, _22939_);
  nand _56415_ (_22942_, _22941_, _22938_);
  nor _56416_ (_22943_, _22942_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56417_ (_22944_, _22943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _56418_ (_22945_, _22944_);
  nor _56419_ (_22946_, _22945_, _22935_);
  nand _56420_ (_22947_, _22660_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _56421_ (_22948_, _22658_, _09507_);
  not _56422_ (_22949_, _22948_);
  nand _56423_ (_22950_, _22949_, _22947_);
  nand _56424_ (_22951_, _22662_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nand _56425_ (_22952_, _22653_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nand _56426_ (_22953_, _22952_, _22951_);
  nor _56427_ (_22954_, _22953_, _22950_);
  nor _56428_ (_22955_, _22954_, _22683_);
  nor _56429_ (_22956_, _22669_, _10546_);
  nand _56430_ (_22957_, _22662_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  not _56431_ (_22958_, _22957_);
  nor _56432_ (_22959_, _22958_, _22956_);
  nor _56433_ (_22960_, _22658_, _10548_);
  nand _56434_ (_22961_, _22653_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  not _56435_ (_22962_, _22961_);
  nor _56436_ (_22963_, _22962_, _22960_);
  nand _56437_ (_22964_, _22963_, _22959_);
  nand _56438_ (_22965_, _22964_, _22460_);
  not _56439_ (_22966_, _22965_);
  nor _56440_ (_22967_, _22966_, _22955_);
  not _56441_ (_22968_, _22967_);
  nor _56442_ (_22969_, _22968_, _22946_);
  not _56443_ (_22970_, _22969_);
  nor _56444_ (_22971_, _22970_, _22925_);
  nand _56445_ (_22972_, _22971_, _22923_);
  nor _56446_ (_22973_, _22969_, _22652_);
  nor _56447_ (_22974_, _22658_, _08938_);
  nand _56448_ (_22975_, _22660_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  not _56449_ (_22976_, _22975_);
  nor _56450_ (_22977_, _22976_, _22974_);
  nor _56451_ (_22978_, _22672_, _08815_);
  nand _56452_ (_22979_, _22662_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  not _56453_ (_22980_, _22979_);
  nor _56454_ (_22981_, _22980_, _22978_);
  nand _56455_ (_22982_, _22981_, _22977_);
  nor _56456_ (_22983_, _22982_, _00047_);
  nand _56457_ (_22984_, _22660_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _56458_ (_22985_, _22657_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand _56459_ (_22986_, _22985_, _22984_);
  nand _56460_ (_22987_, _22662_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand _56461_ (_22988_, _22653_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _56462_ (_22989_, _22988_, _22987_);
  nor _56463_ (_22990_, _22989_, _22986_);
  nand _56464_ (_22991_, _22990_, _00047_);
  nand _56465_ (_22992_, _22991_, _00051_);
  nor _56466_ (_22993_, _22992_, _22983_);
  nand _56467_ (_22994_, _22660_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nand _56468_ (_22995_, _22657_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nand _56469_ (_22996_, _22995_, _22994_);
  nand _56470_ (_22997_, _22662_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _56471_ (_22998_, _22672_, _09300_);
  not _56472_ (_22999_, _22998_);
  nand _56473_ (_23000_, _22999_, _22997_);
  nor _56474_ (_23001_, _23000_, _22996_);
  nor _56475_ (_23002_, _23001_, _22683_);
  nand _56476_ (_23003_, _22660_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nand _56477_ (_23004_, _22662_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nand _56478_ (_23005_, _23004_, _23003_);
  nand _56479_ (_23006_, _22657_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nand _56480_ (_23007_, _22653_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nand _56481_ (_23008_, _23007_, _23006_);
  nor _56482_ (_23009_, _23008_, _23005_);
  nor _56483_ (_23010_, _23009_, _22461_);
  nor _56484_ (_23011_, _23010_, _23002_);
  not _56485_ (_23012_, _23011_);
  nor _56486_ (_23013_, _23012_, _22993_);
  nor _56487_ (_23014_, _23013_, _22652_);
  nor _56488_ (_23015_, _23014_, _22831_);
  nand _56489_ (_23016_, _23015_, _22872_);
  not _56490_ (_23017_, _23016_);
  nand _56491_ (_23018_, _23017_, _22973_);
  nand _56492_ (_23019_, _23018_, _22972_);
  nor _56493_ (_23020_, _23019_, _22919_);
  not _56494_ (_23021_, _22748_);
  nand _56495_ (_23022_, _23014_, _22830_);
  nor _56496_ (_23023_, _23022_, _22922_);
  not _56497_ (_23024_, _23023_);
  nor _56498_ (_23025_, _23024_, _22924_);
  not _56499_ (_23026_, _23025_);
  nand _56500_ (_23027_, _23026_, _23021_);
  not _56501_ (_23028_, _22973_);
  nor _56502_ (_23029_, _23024_, _23028_);
  not _56503_ (_23030_, _23029_);
  nand _56504_ (_23031_, _23017_, _23028_);
  nand _56505_ (_23032_, _23031_, _23030_);
  nor _56506_ (_23033_, _23032_, _23027_);
  nor _56507_ (_23034_, _23033_, _23020_);
  nand _56508_ (_23035_, _23017_, _22920_);
  nor _56509_ (_23036_, _23035_, _22973_);
  nor _56510_ (_23038_, _23036_, _23034_);
  nor _56511_ (_23039_, _23038_, _22706_);
  nor _56512_ (_23040_, _23024_, _22973_);
  not _56513_ (_23041_, _22923_);
  nor _56514_ (_23042_, _23028_, _23041_);
  nor _56515_ (_23043_, _23042_, _23021_);
  nand _56516_ (_23044_, _22924_, _22831_);
  nor _56517_ (_23045_, _23044_, _23028_);
  nand _56518_ (_23046_, _23015_, _22921_);
  nor _56519_ (_23047_, _22969_, _22925_);
  nand _56520_ (_23048_, _23047_, _22915_);
  nand _56521_ (_23049_, _23048_, _23046_);
  nor _56522_ (_23050_, _23049_, _23045_);
  nand _56523_ (_23051_, _23050_, _23035_);
  nor _56524_ (_23052_, _23051_, _23027_);
  nor _56525_ (_23053_, _23052_, _23043_);
  nor _56526_ (_23054_, _23053_, _23040_);
  nor _56527_ (_23055_, _23054_, _22705_);
  nor _56528_ (_23056_, _23055_, _23039_);
  nor _56529_ (_23057_, _23056_, _22604_);
  nand _56530_ (_23059_, _22831_, _22704_);
  not _56531_ (_23060_, _22831_);
  nand _56532_ (_23061_, _23060_, _22787_);
  nand _56533_ (_23062_, _23061_, _23059_);
  nor _56534_ (_23063_, _22973_, _22916_);
  nand _56535_ (_23064_, _23063_, _23062_);
  nor _56536_ (_23065_, _23014_, _22872_);
  nand _56537_ (_23066_, _23065_, _23060_);
  nor _56538_ (_23067_, _23022_, _22914_);
  not _56539_ (_23068_, _22830_);
  nor _56540_ (_23069_, _23013_, _23068_);
  nor _56541_ (_23070_, _23069_, _23028_);
  nor _56542_ (_23071_, _23070_, _23067_);
  nand _56543_ (_23072_, _23071_, _23066_);
  nand _56544_ (_23073_, _23072_, _22705_);
  nor _56545_ (_23074_, _22917_, _22748_);
  nand _56546_ (_23075_, _23074_, _23073_);
  not _56547_ (_23076_, _23065_);
  nor _56548_ (_23077_, _23014_, _22920_);
  nand _56549_ (_23078_, _23077_, _22925_);
  nand _56550_ (_23079_, _23078_, _23076_);
  nand _56551_ (_23080_, _23079_, _23028_);
  nand _56552_ (_23081_, _23080_, _22916_);
  nand _56553_ (_23082_, _23081_, _22706_);
  nand _56554_ (_23083_, _22923_, _22925_);
  nor _56555_ (_23084_, _23014_, _22973_);
  nor _56556_ (_23085_, _23028_, _22704_);
  nor _56557_ (_23086_, _23085_, _23084_);
  nor _56558_ (_23087_, _23086_, _23083_);
  nand _56559_ (_23088_, _23067_, _22872_);
  nor _56560_ (_23089_, _23044_, _22973_);
  nor _56561_ (_23090_, _23089_, _23021_);
  nand _56562_ (_23091_, _23090_, _23088_);
  nor _56563_ (_23092_, _23091_, _23087_);
  nand _56564_ (_23093_, _23092_, _23082_);
  nand _56565_ (_23094_, _23093_, _23075_);
  nand _56566_ (_23095_, _23094_, _23064_);
  nor _56567_ (_23096_, _00091_, _00087_);
  nor _56568_ (_23097_, _22487_, _00083_);
  not _56569_ (_23098_, _23097_);
  nor _56570_ (_23099_, _22669_, _22461_);
  not _56571_ (_23100_, _23099_);
  nor _56572_ (_23101_, _23100_, _22459_);
  not _56573_ (_23102_, _23101_);
  nor _56574_ (_23103_, _23102_, _23098_);
  nand _56575_ (_23104_, _23103_, _23096_);
  nor _56576_ (_23105_, _23104_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not _56577_ (_23106_, _23104_);
  nor _56578_ (_23107_, _23106_, _00095_);
  nor _56579_ (_23108_, _23107_, _23105_);
  not _56580_ (_23109_, _23108_);
  nand _56581_ (_23110_, _23109_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _56582_ (_23111_, _23108_, _00035_);
  nand _56583_ (_23112_, _23111_, _23110_);
  nand _56584_ (_23113_, _22496_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand _56585_ (_23114_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _00039_);
  nand _56586_ (_23115_, _23114_, _23113_);
  nand _56587_ (_23116_, _23115_, _00031_);
  nand _56588_ (_23117_, _23116_, _23112_);
  nor _56589_ (_23118_, _23102_, _22487_);
  not _56590_ (_23119_, _23118_);
  nand _56591_ (_23120_, _23119_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nand _56592_ (_23121_, _23118_, _00083_);
  nand _56593_ (_23122_, _23121_, _23120_);
  nand _56594_ (_23123_, _23122_, _00023_);
  nand _56595_ (_23124_, _00063_, _00039_);
  nor _56596_ (_23125_, _23100_, _22457_);
  nor _56597_ (_23126_, _23125_, _22577_);
  nand _56598_ (_23127_, _23126_, _23124_);
  nand _56599_ (_23128_, _23127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _56600_ (_23129_, _22558_, _00039_);
  nor _56601_ (_23130_, _23100_, _00055_);
  nor _56602_ (_23131_, _23130_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _56603_ (_23132_, _23131_, _23129_);
  nand _56604_ (_23133_, _23132_, _28131_);
  nand _56605_ (_23134_, _23133_, _23128_);
  nor _56606_ (_23135_, _23132_, _28131_);
  not _56607_ (_23136_, _22523_);
  nor _56608_ (_23137_, _22657_, _22653_);
  not _56609_ (_23138_, _23137_);
  nor _56610_ (_23139_, _23138_, _28115_);
  nor _56611_ (_23140_, _23137_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _56612_ (_23141_, _23140_, _23139_);
  nand _56613_ (_23142_, _23141_, _23136_);
  nor _56614_ (_23143_, _23142_, _23135_);
  nor _56615_ (_23144_, _22669_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _56616_ (_23145_, _22660_, _00047_);
  nor _56617_ (_23146_, _23145_, _23144_);
  not _56618_ (_23147_, _23146_);
  nand _56619_ (_23148_, _23147_, _28119_);
  nand _56620_ (_23149_, _23146_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _56621_ (_23150_, _23149_, _23148_);
  nor _56622_ (_23151_, _22669_, _00047_);
  nor _56623_ (_23152_, _23151_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56624_ (_23153_, _23152_, _23099_);
  not _56625_ (_23154_, _23153_);
  nand _56626_ (_23155_, _23154_, _28123_);
  nand _56627_ (_23156_, _23153_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56628_ (_23157_, _23156_, _23155_);
  nor _56629_ (_23158_, _23125_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _56630_ (_23159_, _23158_, _23101_);
  nor _56631_ (_23160_, _23159_, _00006_);
  nor _56632_ (_23161_, _23100_, _22545_);
  nor _56633_ (_23162_, _23099_, _22519_);
  nor _56634_ (_23163_, _23162_, _23161_);
  nor _56635_ (_23164_, _23163_, _23160_);
  nand _56636_ (_23165_, _23164_, _23157_);
  nor _56637_ (_23166_, _23165_, _23150_);
  nand _56638_ (_23167_, _23166_, _23143_);
  nor _56639_ (_23168_, _23167_, _23134_);
  nand _56640_ (_23169_, _23168_, _23123_);
  nor _56641_ (_23170_, _23169_, _23117_);
  nand _56642_ (_23171_, _00079_, _00039_);
  nor _56643_ (_23172_, _23118_, _22592_);
  nand _56644_ (_23173_, _23172_, _23171_);
  nor _56645_ (_23174_, _23173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _56646_ (_23175_, _23104_, _00095_);
  nor _56647_ (_23176_, _23175_, _24873_);
  nand _56648_ (_23177_, _23175_, _24873_);
  not _56649_ (_23178_, _23177_);
  nor _56650_ (_23179_, _23178_, _23176_);
  not _56651_ (_23180_, _23179_);
  nor _56652_ (_23181_, _23180_, _24868_);
  nor _56653_ (_23182_, _23181_, _23174_);
  nor _56654_ (_23183_, _23179_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _56655_ (_23184_, _22472_, _00039_);
  not _56656_ (_23185_, _23184_);
  nor _56657_ (_23186_, _23185_, _00087_);
  nor _56658_ (_23187_, _23184_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _56659_ (_23188_, _23187_, _23186_);
  not _56660_ (_23189_, _23188_);
  nand _56661_ (_23190_, _23189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _56662_ (_23191_, _23188_, _00027_);
  nand _56663_ (_23192_, _23191_, _23190_);
  nor _56664_ (_23193_, _23192_, _23183_);
  nand _56665_ (_23194_, _23193_, _23182_);
  nand _56666_ (_23195_, _23173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _56667_ (_23196_, _23159_, _00006_);
  nand _56668_ (_23197_, _23196_, _23195_);
  nor _56669_ (_23198_, _23102_, _00071_);
  not _56670_ (_23200_, _23198_);
  nor _56671_ (_23201_, _23200_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _56672_ (_23202_, _23198_, _00075_);
  nor _56673_ (_23203_, _23202_, _23201_);
  not _56674_ (_23204_, _23203_);
  nor _56675_ (_23205_, _23204_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _56676_ (_23206_, _23203_, _00014_);
  nor _56677_ (_23207_, _23206_, _23205_);
  nor _56678_ (_23208_, _23207_, _23197_);
  nor _56679_ (_23209_, _23115_, _00031_);
  nor _56680_ (_23210_, _23127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _56681_ (_23211_, _23122_, _00023_);
  nor _56682_ (_23212_, _23211_, _23210_);
  nor _56683_ (_23213_, _22468_, _00039_);
  nor _56684_ (_23214_, _23101_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _56685_ (_23215_, _23214_, _23213_);
  not _56686_ (_23216_, _23215_);
  nor _56687_ (_23217_, _23216_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _56688_ (_23218_, _23215_, _00010_);
  nor _56689_ (_23219_, _23218_, _23217_);
  nand _56690_ (_23220_, _23219_, _23212_);
  nor _56691_ (_23221_, _23220_, _23209_);
  nand _56692_ (_23222_, _23221_, _23208_);
  nor _56693_ (_23223_, _23222_, _23194_);
  nand _56694_ (_23224_, _23223_, _23170_);
  nand _56695_ (_23225_, _23224_, _23095_);
  nor _56696_ (_23226_, _22662_, _22461_);
  not _56697_ (_23227_, _23226_);
  nor _56698_ (_23228_, _23227_, _22459_);
  not _56699_ (_23229_, _23228_);
  nor _56700_ (_23230_, _23229_, _22487_);
  not _56701_ (_23231_, _23230_);
  nor _56702_ (_23232_, _23231_, _00083_);
  not _56703_ (_23233_, _23232_);
  nor _56704_ (_23234_, _23233_, _00087_);
  nor _56705_ (_23235_, _23232_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _56706_ (_23236_, _23235_, _23234_);
  nor _56707_ (_23237_, _23236_, _00027_);
  nand _56708_ (_23238_, _23236_, _00027_);
  nand _56709_ (_23239_, _23226_, _22456_);
  nor _56710_ (_23240_, _23239_, _00063_);
  nor _56711_ (_23241_, _23240_, _00067_);
  not _56712_ (_23242_, _23240_);
  nor _56713_ (_23243_, _23242_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _56714_ (_23244_, _23243_, _23241_);
  not _56715_ (_23245_, _23244_);
  nand _56716_ (_23246_, _23245_, _00006_);
  nand _56717_ (_23247_, _23244_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand _56718_ (_23248_, _23247_, _23246_);
  nor _56719_ (_23249_, _23229_, _00071_);
  nor _56720_ (_23250_, _23228_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _56721_ (_23251_, _23250_, _23249_);
  not _56722_ (_23252_, _23251_);
  nand _56723_ (_23253_, _23252_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _56724_ (_23254_, _23251_, _00010_);
  nand _56725_ (_23255_, _23254_, _23253_);
  nor _56726_ (_23256_, _23255_, _23248_);
  nand _56727_ (_23257_, _23256_, _23238_);
  nor _56728_ (_23258_, _23257_, _23237_);
  nand _56729_ (_23259_, _23231_, _00083_);
  nand _56730_ (_23260_, _23259_, _23233_);
  nand _56731_ (_23261_, _23260_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _56732_ (_23262_, _23260_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _56733_ (_23263_, _23249_);
  nor _56734_ (_23264_, _23263_, _00075_);
  nor _56735_ (_23265_, _23249_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _56736_ (_23266_, _23265_, _23264_);
  nor _56737_ (_23267_, _23266_, _00014_);
  nor _56738_ (_23268_, _23267_, _23262_);
  nand _56739_ (_23269_, _23268_, _23261_);
  nand _56740_ (_23270_, _23239_, _00063_);
  nand _56741_ (_23271_, _23270_, _23242_);
  nor _56742_ (_23272_, _23271_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _56743_ (_23273_, _23227_, _00055_);
  nor _56744_ (_23274_, _23273_, _22514_);
  nand _56745_ (_23275_, _23273_, _22514_);
  nor _56746_ (_23276_, _22519_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56747_ (_23277_, _23276_, _23226_);
  nor _56748_ (_23278_, _22662_, _00047_);
  nor _56749_ (_23279_, _23278_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _56750_ (_23280_, _23279_, _22519_);
  not _56751_ (_23281_, _23280_);
  nand _56752_ (_23282_, _23281_, _23277_);
  nand _56753_ (_23283_, _23282_, _23275_);
  nor _56754_ (_23284_, _23283_, _23274_);
  nor _56755_ (_23285_, _23280_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56756_ (_23286_, _23285_, _23277_);
  nor _56757_ (_23287_, _23141_, _22523_);
  nand _56758_ (_23288_, _22672_, _22640_);
  not _56759_ (_23289_, _23288_);
  nor _56760_ (_23290_, _23289_, _23278_);
  nor _56761_ (_23291_, _23290_, _28119_);
  not _56762_ (_23292_, _23290_);
  nor _56763_ (_23293_, _23292_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _56764_ (_23294_, _23293_, _23291_);
  nand _56765_ (_23295_, _23294_, _23287_);
  nor _56766_ (_23296_, _23295_, _23286_);
  nand _56767_ (_23297_, _23296_, _23284_);
  nor _56768_ (_23298_, _23297_, _23272_);
  not _56769_ (_23299_, _23266_);
  nor _56770_ (_23300_, _23299_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not _56771_ (_23301_, _23271_);
  nor _56772_ (_23302_, _23301_, _00001_);
  nor _56773_ (_23303_, _23302_, _23300_);
  nand _56774_ (_23304_, _23303_, _23298_);
  nor _56775_ (_23305_, _23304_, _23269_);
  nand _56776_ (_23306_, _23305_, _23258_);
  nand _56777_ (_23307_, _23234_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _56778_ (_23308_, _23307_, _00095_);
  not _56779_ (_23309_, _23307_);
  nor _56780_ (_23310_, _23309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _56781_ (_23311_, _23310_, _23308_);
  not _56782_ (_23312_, _23311_);
  nand _56783_ (_23313_, _23312_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _56784_ (_23314_, _23311_, _00035_);
  nand _56785_ (_23315_, _23314_, _23313_);
  nor _56786_ (_23316_, _23315_, _23306_);
  nor _56787_ (_23317_, _23308_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  not _56788_ (_23318_, _23308_);
  nor _56789_ (_23319_, _23318_, _24873_);
  nor _56790_ (_23320_, _23319_, _23317_);
  nor _56791_ (_23321_, _23320_, _24868_);
  nand _56792_ (_23322_, _23320_, _24868_);
  nor _56793_ (_23323_, _23234_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _56794_ (_23324_, _23323_, _23309_);
  nor _56795_ (_23325_, _23324_, _00031_);
  nand _56796_ (_23326_, _23324_, _00031_);
  nor _56797_ (_23327_, _23264_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _56798_ (_23328_, _23327_, _23230_);
  nor _56799_ (_23329_, _23328_, _00018_);
  not _56800_ (_23330_, _23328_);
  nor _56801_ (_23331_, _23330_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _56802_ (_23332_, _23331_, _23329_);
  nand _56803_ (_23333_, _23332_, _23326_);
  nor _56804_ (_23334_, _23333_, _23325_);
  nand _56805_ (_23335_, _23334_, _23322_);
  nor _56806_ (_23336_, _23335_, _23321_);
  nand _56807_ (_23337_, _23336_, _23316_);
  not _56808_ (_23338_, _23047_);
  not _56809_ (_23339_, _23088_);
  nand _56810_ (_23340_, _23339_, _23338_);
  nand _56811_ (_23341_, _23029_, _22924_);
  nand _56812_ (_23342_, _23341_, _23340_);
  nor _56813_ (_23343_, _22748_, _22703_);
  nand _56814_ (_23344_, _23343_, _23342_);
  not _56815_ (_23345_, _22920_);
  not _56816_ (_23346_, _22971_);
  nor _56817_ (_23347_, _23016_, _23346_);
  nand _56818_ (_23348_, _23347_, _23345_);
  nand _56819_ (_23349_, _23025_, _23028_);
  nand _56820_ (_23351_, _23349_, _23348_);
  nor _56821_ (_23352_, _22747_, _22706_);
  nand _56822_ (_23353_, _23352_, _23351_);
  nand _56823_ (_23354_, _23353_, _23344_);
  nand _56824_ (_23355_, _23354_, _23337_);
  nand _56825_ (_23356_, _23355_, _23225_);
  nor _56826_ (_23357_, _23356_, _23057_);
  nor _56827_ (_23358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _56828_ (_23359_, _23358_, _28119_);
  not _56829_ (_23360_, _23359_);
  nand _56830_ (_23361_, _23358_, _28119_);
  nand _56831_ (_23362_, _23361_, _23360_);
  nor _56832_ (_23363_, _23359_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56833_ (_23364_, _23360_, _28123_);
  nor _56834_ (_23365_, _23364_, _23363_);
  nor _56835_ (_23366_, _23365_, _06909_);
  not _56836_ (_23367_, _23365_);
  nor _56837_ (_23368_, _23367_, _06915_);
  nor _56838_ (_23369_, _23368_, _23366_);
  nand _56839_ (_23370_, _23369_, _23362_);
  nor _56840_ (_23371_, _07469_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _56841_ (_23372_, _23362_);
  nand _56842_ (_23373_, _23365_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand _56843_ (_23374_, _23373_, _23372_);
  nor _56844_ (_23375_, _23374_, _23371_);
  nor _56845_ (_23376_, _23375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _56846_ (_23377_, _23376_, _23370_);
  nand _56847_ (_23378_, _23365_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _56848_ (_23379_, _06928_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56849_ (_23380_, _23379_, _23362_);
  nand _56850_ (_23381_, _23380_, _23378_);
  nand _56851_ (_23382_, _23367_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _56852_ (_23383_, _23365_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _56853_ (_23384_, _23383_, _23382_);
  nor _56854_ (_23385_, _23384_, _23372_);
  nor _56855_ (_23386_, _23385_, _28115_);
  nand _56856_ (_23387_, _23386_, _23381_);
  nand _56857_ (_23388_, _23387_, _23377_);
  nor _56858_ (_23389_, _28119_, _28115_);
  not _56859_ (_23390_, _23389_);
  nor _56860_ (_23391_, _23390_, _28110_);
  nor _56861_ (_23392_, _28115_, _28110_);
  nor _56862_ (_23393_, _23392_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _56863_ (_23394_, _23393_, _23391_);
  not _56864_ (_23395_, _23394_);
  nor _56865_ (_23396_, _23391_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56866_ (_23397_, _23391_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _56867_ (_23398_, _23397_);
  nor _56868_ (_23399_, _23398_, _23396_);
  nor _56869_ (_23400_, _23399_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _56870_ (_23401_, \oc8051_symbolic_cxrom1.regvalid [14], _28123_);
  nor _56871_ (_23402_, _23401_, _23400_);
  nor _56872_ (_23403_, _23402_, _23395_);
  not _56873_ (_23404_, _23399_);
  nor _56874_ (_23405_, _23404_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _56875_ (_23406_, _23399_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _56876_ (_23407_, _23406_, _23405_);
  nor _56877_ (_23408_, _23407_, _23394_);
  nor _56878_ (_23409_, _23408_, _23403_);
  nor _56879_ (_23410_, _23409_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _56880_ (_23411_, _23399_, _06915_);
  nor _56881_ (_23412_, _23399_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _56882_ (_23413_, _23412_, _23394_);
  nand _56883_ (_23414_, _23413_, _23411_);
  nor _56884_ (_23415_, _23399_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand _56885_ (_23416_, _07886_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56886_ (_23417_, _23416_, _23394_);
  nor _56887_ (_23418_, _23417_, _23415_);
  nor _56888_ (_23419_, _23418_, _28115_);
  nand _56889_ (_23420_, _23419_, _23414_);
  not _56890_ (_23421_, _23392_);
  nand _56891_ (_23422_, _06876_, _28123_);
  nand _56892_ (_23423_, _06862_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56893_ (_23424_, _23423_, _23422_);
  nand _56894_ (_23425_, _23424_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _56895_ (_23426_, _06852_, _28123_);
  nand _56896_ (_23427_, _06871_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56897_ (_23428_, _23427_, _23426_);
  nand _56898_ (_23429_, _23428_, _28119_);
  nand _56899_ (_23430_, _23429_, _23425_);
  nor _56900_ (_23431_, _23430_, _23421_);
  nand _56901_ (_23432_, _28115_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _56902_ (_23433_, _06888_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56903_ (_23434_, _06891_, _28123_);
  nor _56904_ (_23435_, _23434_, _23433_);
  nand _56905_ (_23436_, _23435_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _56906_ (_23437_, _06897_, _28123_);
  nand _56907_ (_23438_, _06895_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56908_ (_23439_, _23438_, _23437_);
  nand _56909_ (_23440_, _23439_, _28119_);
  nand _56910_ (_23441_, _23440_, _23436_);
  nor _56911_ (_23442_, _23441_, _23432_);
  nor _56912_ (_23443_, _23442_, _23431_);
  nor _56913_ (_23444_, _23430_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _56914_ (_23445_, _23435_);
  nor _56915_ (_23446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], _28115_);
  nand _56916_ (_23447_, _23446_, _23445_);
  nand _56917_ (_23448_, _06895_, _28123_);
  nor _56918_ (_23449_, \oc8051_symbolic_cxrom1.regvalid [1], _28123_);
  nor _56919_ (_23450_, _23449_, _23390_);
  nand _56920_ (_23451_, _23450_, _23448_);
  nand _56921_ (_23452_, _23451_, _23447_);
  nor _56922_ (_23453_, _23452_, _23444_);
  nor _56923_ (_23454_, _23453_, _23443_);
  nand _56924_ (_23455_, _23454_, _23420_);
  nor _56925_ (_23456_, _23455_, _23410_);
  nand _56926_ (_23457_, _23456_, _23388_);
  nor _56927_ (_23458_, _23399_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _56928_ (_23459_, _23423_, _23394_);
  nor _56929_ (_23460_, _23459_, _23458_);
  nor _56930_ (_23461_, _23399_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _56931_ (_23462_, _23399_, _06871_);
  nand _56932_ (_23463_, _23462_, _23395_);
  nor _56933_ (_23464_, _23463_, _23461_);
  nor _56934_ (_23465_, _23464_, _23460_);
  nand _56935_ (_23466_, _23465_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _56936_ (_23467_, _23365_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _56937_ (_23468_, _06876_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56938_ (_23469_, _23468_, _23362_);
  nand _56939_ (_23470_, _23469_, _23467_);
  nand _56940_ (_23471_, _23470_, _28115_);
  nor _56941_ (_23472_, _23367_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _56942_ (_23473_, _23365_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _56943_ (_23474_, _23473_, _23472_);
  nor _56944_ (_23475_, _23474_, _23372_);
  nor _56945_ (_23476_, _23475_, _23471_);
  nor _56946_ (_23477_, _23476_, _23452_);
  nand _56947_ (_23478_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56948_ (_23479_, \oc8051_symbolic_cxrom1.regvalid [0], _28123_);
  nand _56949_ (_23480_, _23479_, _23478_);
  nand _56950_ (_23482_, _23480_, _28119_);
  not _56951_ (_23483_, _23371_);
  nand _56952_ (_23484_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56953_ (_23485_, _23484_, _23483_);
  nand _56954_ (_23486_, _23485_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _56955_ (_23487_, _23486_, _23482_);
  nand _56956_ (_23488_, _23487_, _28115_);
  nor _56957_ (_23489_, _07937_, _28123_);
  nor _56958_ (_23490_, _23379_, _28119_);
  not _56959_ (_23491_, _23490_);
  nor _56960_ (_23492_, _23491_, _23489_);
  nor _56961_ (_23493_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _56962_ (_23494_, \oc8051_symbolic_cxrom1.regvalid [10], _28123_);
  nor _56963_ (_23495_, _23494_, _23493_);
  nor _56964_ (_23496_, _23495_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _56965_ (_23497_, _23496_, _23492_);
  nand _56966_ (_23498_, _23497_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _56967_ (_23499_, _23498_, _23488_);
  nand _56968_ (_23500_, _23499_, _28110_);
  nand _56969_ (_23501_, _23485_, _23446_);
  nand _56970_ (_23502_, _06915_, _28123_);
  nor _56971_ (_23503_, \oc8051_symbolic_cxrom1.regvalid [0], _28123_);
  nor _56972_ (_23504_, _23503_, _23390_);
  nand _56973_ (_23505_, _23504_, _23502_);
  nand _56974_ (_23506_, _23505_, _23501_);
  not _56975_ (_23507_, _23497_);
  nor _56976_ (_23508_, _23507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _56977_ (_23509_, _23508_, _23506_);
  nor _56978_ (_23510_, _23509_, _23500_);
  nor _56979_ (_23511_, _23399_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand _56980_ (_23512_, _06891_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _56981_ (_23513_, _23512_, _23394_);
  nor _56982_ (_23514_, _23513_, _23511_);
  nor _56983_ (_23515_, _23399_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand _56984_ (_23516_, _23399_, _06895_);
  nand _56985_ (_23517_, _23516_, _23395_);
  nor _56986_ (_23518_, _23517_, _23515_);
  nor _56987_ (_23519_, _23518_, _23514_);
  nand _56988_ (_23520_, _23519_, _28115_);
  nand _56989_ (_23521_, _23520_, _23510_);
  nor _56990_ (_23522_, _23521_, _23477_);
  nand _56991_ (_23523_, _23522_, _23466_);
  nand _56992_ (_23524_, _23523_, _23457_);
  nand _56993_ (_23525_, _23154_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand _56994_ (_23526_, _23153_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nand _56995_ (_23527_, _23526_, _23525_);
  nand _56996_ (_23528_, _23527_, _23147_);
  nand _56997_ (_23529_, _23153_, _06895_);
  nor _56998_ (_23530_, _23153_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _56999_ (_23531_, _23530_, _23147_);
  nand _57000_ (_23532_, _23531_, _23529_);
  nand _57001_ (_23533_, _23532_, _23528_);
  nand _57002_ (_23534_, _23533_, _22662_);
  nand _57003_ (_23535_, _23154_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand _57004_ (_23536_, _23153_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nand _57005_ (_23537_, _23536_, _23535_);
  nand _57006_ (_23538_, _23537_, _23147_);
  nand _57007_ (_23539_, _23153_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _57008_ (_23540_, _23154_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _57009_ (_23541_, _23540_, _23539_);
  nand _57010_ (_23542_, _23541_, _23146_);
  nand _57011_ (_23543_, _23542_, _23538_);
  nand _57012_ (_23544_, _23543_, _22653_);
  nand _57013_ (_23545_, _23544_, _23534_);
  nand _57014_ (_23546_, _23153_, _07886_);
  nor _57015_ (_23547_, _23153_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _57016_ (_23548_, _23547_, _23146_);
  nand _57017_ (_23549_, _23548_, _23546_);
  nand _57018_ (_23550_, _23153_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _57019_ (_23551_, _23154_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand _57020_ (_23553_, _23551_, _23550_);
  nand _57021_ (_23554_, _23553_, _23146_);
  nand _57022_ (_23555_, _23554_, _23549_);
  nand _57023_ (_23556_, _23555_, _22660_);
  nand _57024_ (_23557_, _23154_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _57025_ (_23558_, _23153_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand _57026_ (_23559_, _23558_, _23557_);
  nand _57027_ (_23560_, _23559_, _23147_);
  nand _57028_ (_23561_, _23153_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand _57029_ (_23562_, _23154_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _57030_ (_23563_, _23562_, _23561_);
  nand _57031_ (_23564_, _23563_, _23146_);
  nand _57032_ (_23565_, _23564_, _23560_);
  nand _57033_ (_23566_, _23565_, _22657_);
  nand _57034_ (_23567_, _23566_, _23556_);
  nor _57035_ (_23568_, _23567_, _23545_);
  nor _57036_ (_23569_, _23279_, _23226_);
  not _57037_ (_23570_, _23569_);
  nor _57038_ (_23571_, _23570_, _06895_);
  nor _57039_ (_23572_, _23569_, _06897_);
  nor _57040_ (_23573_, _23572_, _23571_);
  nor _57041_ (_23574_, _23573_, _22658_);
  nor _57042_ (_23575_, _23574_, _23290_);
  nor _57043_ (_23576_, _23570_, _06932_);
  nor _57044_ (_23577_, _23569_, _06935_);
  nor _57045_ (_23578_, _23577_, _23576_);
  nor _57046_ (_23579_, _23578_, _22669_);
  nand _57047_ (_23580_, _23569_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand _57048_ (_23581_, _23570_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _57049_ (_23582_, _23581_, _23580_);
  nand _57050_ (_23583_, _23582_, _22662_);
  nand _57051_ (_23584_, _23569_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _57052_ (_23585_, _23570_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand _57053_ (_23586_, _23585_, _23584_);
  nand _57054_ (_23587_, _23586_, _22653_);
  nand _57055_ (_23588_, _23587_, _23583_);
  nor _57056_ (_23589_, _23588_, _23579_);
  nand _57057_ (_23590_, _23589_, _23575_);
  nand _57058_ (_23591_, _23570_, _06888_);
  nor _57059_ (_23592_, _22658_, _22645_);
  nand _57060_ (_23593_, _23592_, _23591_);
  nand _57061_ (_23594_, _23593_, _23290_);
  nand _57062_ (_23595_, _23570_, _06928_);
  nor _57063_ (_23596_, _22669_, _22606_);
  nand _57064_ (_23597_, _23596_, _23595_);
  nor _57065_ (_23598_, _23569_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _57066_ (_23599_, _22630_);
  nand _57067_ (_23600_, _22662_, _23599_);
  nor _57068_ (_23601_, _23600_, _23598_);
  nor _57069_ (_23602_, _23569_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not _57070_ (_23603_, _22620_);
  nand _57071_ (_23604_, _22653_, _23603_);
  nor _57072_ (_23605_, _23604_, _23602_);
  nor _57073_ (_23606_, _23605_, _23601_);
  nand _57074_ (_23607_, _23606_, _23597_);
  nor _57075_ (_23608_, _23607_, _23594_);
  not _57076_ (_23609_, _22614_);
  nand _57077_ (_23610_, _23609_, _00043_);
  not _57078_ (_23611_, _22541_);
  not _57079_ (_23612_, _22622_);
  nor _57080_ (_23613_, _23612_, _23611_);
  nand _57081_ (_23614_, _22533_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _57082_ (_23615_, _22463_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand _57083_ (_23616_, _23615_, _23614_);
  nor _57084_ (_23617_, _23616_, _23613_);
  nand _57085_ (_23618_, _23617_, _23610_);
  nand _57086_ (_23619_, _23618_, _00039_);
  nor _57087_ (_23620_, _22672_, _22638_);
  nand _57088_ (_23621_, \oc8051_symbolic_cxrom1.regvalid [9], _00051_);
  nand _57089_ (_23622_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand _57090_ (_23623_, _23622_, _23621_);
  nand _57091_ (_23624_, _23623_, _23151_);
  nand _57092_ (_23625_, _23144_, _22647_);
  nand _57093_ (_23626_, _23625_, _23624_);
  nor _57094_ (_23627_, _23626_, _23620_);
  nand _57095_ (_23628_, _23627_, _23619_);
  not _57096_ (_23629_, first_instr);
  nand _57097_ (_23630_, _24869_, _23629_);
  nor _57098_ (_23631_, _23630_, _22652_);
  nand _57099_ (_23632_, _23631_, _23628_);
  nor _57100_ (_23633_, _23632_, _23608_);
  nand _57101_ (_23634_, _23633_, _23590_);
  nor _57102_ (_23635_, _23634_, _23568_);
  nand _57103_ (_23636_, _23635_, _23524_);
  nor _57104_ (property_invalid, _23636_, _23357_);
  nand _57105_ (_23637_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  nand _57106_ (_23638_, _08334_, _25099_);
  nand _57107_ (_12007_, _23638_, _23637_);
  nand _57108_ (_23639_, _11542_, _24927_);
  nand _57109_ (_23640_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  nand _57110_ (_28257_, _23640_, _23639_);
  nand _57111_ (_23641_, _11542_, _24789_);
  nand _57112_ (_23642_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  nand _57113_ (_12026_, _23642_, _23641_);
  nand _57114_ (_23643_, _11542_, _25150_);
  nand _57115_ (_23644_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nand _57116_ (_12033_, _23644_, _23643_);
  nand _57117_ (_23645_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  nand _57118_ (_23646_, _08339_, _25099_);
  nand _57119_ (_28298_, _23646_, _23645_);
  nand _57120_ (_23647_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nand _57121_ (_23648_, _08339_, _24830_);
  nand _57122_ (_12065_, _23648_, _23647_);
  nand _57123_ (_23649_, _18523_, _25099_);
  nand _57124_ (_23650_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  nand _57125_ (_12071_, _23650_, _23649_);
  nand _57126_ (_23651_, _18523_, _24830_);
  nand _57127_ (_23652_, _18525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nand _57128_ (_12075_, _23652_, _23651_);
  nand _57129_ (_23653_, _03782_, _24927_);
  nand _57130_ (_23655_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  nand _57131_ (_12082_, _23655_, _23653_);
  nand _57132_ (_23656_, _03782_, _25203_);
  nand _57133_ (_23657_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  nand _57134_ (_12087_, _23657_, _23656_);
  nand _57135_ (_23658_, _07810_, _25039_);
  nand _57136_ (_23659_, _07812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nand _57137_ (_12091_, _23659_, _23658_);
  nand _57138_ (_23660_, _03704_, _25150_);
  nand _57139_ (_23661_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  nand _57140_ (_12106_, _23661_, _23660_);
  nand _57141_ (_23662_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nand _57142_ (_23663_, _08339_, _25203_);
  nand _57143_ (_28299_, _23663_, _23662_);
  nand _57144_ (_23664_, _12010_, _28096_);
  nand _57145_ (_23665_, _12012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nand _57146_ (_12111_, _23665_, _23664_);
  nand _57147_ (_23666_, _03704_, _25039_);
  nand _57148_ (_23667_, _03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nand _57149_ (_12113_, _23667_, _23666_);
  nand _57150_ (_23668_, _18173_, _24789_);
  nand _57151_ (_23669_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  nand _57152_ (_12115_, _23669_, _23668_);
  nand _57153_ (_23670_, _11542_, _24830_);
  nand _57154_ (_23671_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  nand _57155_ (_12119_, _23671_, _23670_);
  nand _57156_ (_23672_, _08340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  nand _57157_ (_23673_, _08339_, _28096_);
  nand _57158_ (_12121_, _23673_, _23672_);
  nand _57159_ (_23674_, _18173_, _25150_);
  nand _57160_ (_23675_, _18175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  nand _57161_ (_12126_, _23675_, _23674_);
  nand _57162_ (_23676_, _03571_, _25203_);
  nand _57163_ (_23677_, _03573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  nand _57164_ (_12130_, _23677_, _23676_);
  nand _57165_ (_23678_, _03561_, _25039_);
  nand _57166_ (_23679_, _03563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  nand _57167_ (_28281_, _23679_, _23678_);
  dff _57168_ (first_instr, _00000_, clk);
  dff _57169_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _28169_[0], clk);
  dff _57170_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _28169_[1], clk);
  dff _57171_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _28169_[2], clk);
  dff _57172_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _28169_[3], clk);
  dff _57173_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _28169_[4], clk);
  dff _57174_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _28169_[5], clk);
  dff _57175_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _28169_[6], clk);
  dff _57176_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _28169_[7], clk);
  dff _57177_ (\oc8051_symbolic_cxrom1.regvalid [0], _28181_, clk);
  dff _57178_ (\oc8051_symbolic_cxrom1.regvalid [1], _28135_[1], clk);
  dff _57179_ (\oc8051_symbolic_cxrom1.regvalid [2], _28135_[2], clk);
  dff _57180_ (\oc8051_symbolic_cxrom1.regvalid [3], _28135_[3], clk);
  dff _57181_ (\oc8051_symbolic_cxrom1.regvalid [4], _28135_[4], clk);
  dff _57182_ (\oc8051_symbolic_cxrom1.regvalid [5], _28135_[5], clk);
  dff _57183_ (\oc8051_symbolic_cxrom1.regvalid [6], _28135_[6], clk);
  dff _57184_ (\oc8051_symbolic_cxrom1.regvalid [7], _28135_[7], clk);
  dff _57185_ (\oc8051_symbolic_cxrom1.regvalid [8], _28135_[8], clk);
  dff _57186_ (\oc8051_symbolic_cxrom1.regvalid [9], _28135_[9], clk);
  dff _57187_ (\oc8051_symbolic_cxrom1.regvalid [10], _28135_[10], clk);
  dff _57188_ (\oc8051_symbolic_cxrom1.regvalid [11], _28135_[11], clk);
  dff _57189_ (\oc8051_symbolic_cxrom1.regvalid [12], _28135_[12], clk);
  dff _57190_ (\oc8051_symbolic_cxrom1.regvalid [13], _28135_[13], clk);
  dff _57191_ (\oc8051_symbolic_cxrom1.regvalid [14], _28135_[14], clk);
  dff _57192_ (\oc8051_symbolic_cxrom1.regvalid [15], _28135_[15], clk);
  dff _57193_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _28174_[0], clk);
  dff _57194_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _28174_[1], clk);
  dff _57195_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _28174_[2], clk);
  dff _57196_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _28174_[3], clk);
  dff _57197_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _28174_[4], clk);
  dff _57198_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _28174_[5], clk);
  dff _57199_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _28174_[6], clk);
  dff _57200_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _28174_[7], clk);
  dff _57201_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _28152_, clk);
  dff _57202_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _28153_, clk);
  dff _57203_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _28154_, clk);
  dff _57204_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _28155_, clk);
  dff _57205_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _28156_, clk);
  dff _57206_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _28157_, clk);
  dff _57207_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _28158_, clk);
  dff _57208_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _28159_, clk);
  dff _57209_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _28175_[0], clk);
  dff _57210_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _28175_[1], clk);
  dff _57211_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _28175_[2], clk);
  dff _57212_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _28175_[3], clk);
  dff _57213_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _28175_[4], clk);
  dff _57214_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _28160_, clk);
  dff _57215_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _28175_[6], clk);
  dff _57216_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _28175_[7], clk);
  dff _57217_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _28176_[0], clk);
  dff _57218_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _28176_[1], clk);
  dff _57219_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _28176_[2], clk);
  dff _57220_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _28176_[3], clk);
  dff _57221_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _28176_[4], clk);
  dff _57222_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _28176_[5], clk);
  dff _57223_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _28176_[6], clk);
  dff _57224_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _28176_[7], clk);
  dff _57225_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _28177_[0], clk);
  dff _57226_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _28177_[1], clk);
  dff _57227_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _28177_[2], clk);
  dff _57228_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _28177_[3], clk);
  dff _57229_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _28177_[4], clk);
  dff _57230_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _28177_[5], clk);
  dff _57231_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _28177_[6], clk);
  dff _57232_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _28177_[7], clk);
  dff _57233_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _28178_[0], clk);
  dff _57234_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _28178_[1], clk);
  dff _57235_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _28178_[2], clk);
  dff _57236_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _28178_[3], clk);
  dff _57237_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _28178_[4], clk);
  dff _57238_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _28178_[5], clk);
  dff _57239_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _28178_[6], clk);
  dff _57240_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _28178_[7], clk);
  dff _57241_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _28179_[0], clk);
  dff _57242_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _28179_[1], clk);
  dff _57243_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _28179_[2], clk);
  dff _57244_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _28179_[3], clk);
  dff _57245_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _28179_[4], clk);
  dff _57246_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _28179_[5], clk);
  dff _57247_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _28179_[6], clk);
  dff _57248_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _28179_[7], clk);
  dff _57249_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _28161_, clk);
  dff _57250_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _28162_, clk);
  dff _57251_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _28163_, clk);
  dff _57252_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _28164_, clk);
  dff _57253_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _28165_, clk);
  dff _57254_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _28166_, clk);
  dff _57255_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _28167_, clk);
  dff _57256_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _28168_, clk);
  dff _57257_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _28180_[0], clk);
  dff _57258_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _28180_[1], clk);
  dff _57259_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _28180_[2], clk);
  dff _57260_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _28180_[3], clk);
  dff _57261_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _28180_[4], clk);
  dff _57262_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _28180_[5], clk);
  dff _57263_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _28180_[6], clk);
  dff _57264_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _28180_[7], clk);
  dff _57265_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _28170_[0], clk);
  dff _57266_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _28170_[1], clk);
  dff _57267_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _28170_[2], clk);
  dff _57268_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _28170_[3], clk);
  dff _57269_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _28170_[4], clk);
  dff _57270_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _28170_[5], clk);
  dff _57271_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _28170_[6], clk);
  dff _57272_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _28170_[7], clk);
  dff _57273_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _28136_, clk);
  dff _57274_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _28137_, clk);
  dff _57275_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _28138_, clk);
  dff _57276_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _28139_, clk);
  dff _57277_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _28140_, clk);
  dff _57278_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _28141_, clk);
  dff _57279_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _28142_, clk);
  dff _57280_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _28143_, clk);
  dff _57281_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _28171_[0], clk);
  dff _57282_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _28171_[1], clk);
  dff _57283_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _28171_[2], clk);
  dff _57284_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _28171_[3], clk);
  dff _57285_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _28171_[4], clk);
  dff _57286_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _28171_[5], clk);
  dff _57287_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _28171_[6], clk);
  dff _57288_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _28171_[7], clk);
  dff _57289_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _28172_[0], clk);
  dff _57290_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _28172_[1], clk);
  dff _57291_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _28172_[2], clk);
  dff _57292_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _28172_[3], clk);
  dff _57293_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _28172_[4], clk);
  dff _57294_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _28172_[5], clk);
  dff _57295_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _28172_[6], clk);
  dff _57296_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _28172_[7], clk);
  dff _57297_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _28144_, clk);
  dff _57298_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _28145_, clk);
  dff _57299_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _28146_, clk);
  dff _57300_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _28147_, clk);
  dff _57301_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _28148_, clk);
  dff _57302_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _28149_, clk);
  dff _57303_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _28150_, clk);
  dff _57304_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _28151_, clk);
  dff _57305_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _28173_[0], clk);
  dff _57306_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _28173_[1], clk);
  dff _57307_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _28173_[2], clk);
  dff _57308_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _28173_[3], clk);
  dff _57309_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _28173_[4], clk);
  dff _57310_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _28173_[5], clk);
  dff _57311_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _28173_[6], clk);
  dff _57312_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _28173_[7], clk);
  dff _57313_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _05317_, clk);
  dff _57314_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _05312_, clk);
  dff _57315_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _05315_, clk);
  dff _57316_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _05326_, clk);
  dff _57317_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _05324_, clk);
  dff _57318_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _04574_, clk);
  dff _57319_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _05360_, clk);
  dff _57320_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _04572_, clk);
  dff _57321_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _05381_, clk);
  dff _57322_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _05389_, clk);
  dff _57323_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _05387_, clk);
  dff _57324_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _05402_, clk);
  dff _57325_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _05395_, clk);
  dff _57326_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _05397_, clk);
  dff _57327_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _05412_, clk);
  dff _57328_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _04578_, clk);
  dff _57329_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11754_, clk);
  dff _57330_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _11888_, clk);
  dff _57331_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11806_, clk);
  dff _57332_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11893_, clk);
  dff _57333_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11733_, clk);
  dff _57334_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11735_, clk);
  dff _57335_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11737_, clk);
  dff _57336_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11803_, clk);
  dff _57337_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11752_, clk);
  dff _57338_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _11801_, clk);
  dff _57339_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11757_, clk);
  dff _57340_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11799_, clk);
  dff _57341_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11760_, clk);
  dff _57342_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11897_, clk);
  dff _57343_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11763_, clk);
  dff _57344_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11766_, clk);
  dff _57345_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _28182_[0], clk);
  dff _57346_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _28182_[1], clk);
  dff _57347_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _28182_[2], clk);
  dff _57348_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _28182_[3], clk);
  dff _57349_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _28182_[4], clk);
  dff _57350_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _28182_[5], clk);
  dff _57351_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _28182_[6], clk);
  dff _57352_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _28182_[7], clk);
  dff _57353_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _28218_[0], clk);
  dff _57354_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _28218_[1], clk);
  dff _57355_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _28218_[2], clk);
  dff _57356_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _28218_[3], clk);
  dff _57357_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _28218_[4], clk);
  dff _57358_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _28218_[5], clk);
  dff _57359_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _28218_[6], clk);
  dff _57360_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _28218_[7], clk);
  dff _57361_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _28219_[0], clk);
  dff _57362_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _28219_[1], clk);
  dff _57363_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _28219_[2], clk);
  dff _57364_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _28219_[3], clk);
  dff _57365_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _28219_[4], clk);
  dff _57366_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _28219_[5], clk);
  dff _57367_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _28219_[6], clk);
  dff _57368_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _28219_[7], clk);
  dff _57369_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _28183_[0], clk);
  dff _57370_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _28183_[1], clk);
  dff _57371_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _28183_[2], clk);
  dff _57372_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _28184_[0], clk);
  dff _57373_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _28184_[1], clk);
  dff _57374_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _28184_[2], clk);
  dff _57375_ (\oc8051_top_1.oc8051_decoder1.state [0], _28185_[0], clk);
  dff _57376_ (\oc8051_top_1.oc8051_decoder1.state [1], _28185_[1], clk);
  dff _57377_ (\oc8051_top_1.oc8051_decoder1.op [0], _28186_[0], clk);
  dff _57378_ (\oc8051_top_1.oc8051_decoder1.op [1], _28186_[1], clk);
  dff _57379_ (\oc8051_top_1.oc8051_decoder1.op [2], _28186_[2], clk);
  dff _57380_ (\oc8051_top_1.oc8051_decoder1.op [3], _28186_[3], clk);
  dff _57381_ (\oc8051_top_1.oc8051_decoder1.op [4], _28186_[4], clk);
  dff _57382_ (\oc8051_top_1.oc8051_decoder1.op [5], _28186_[5], clk);
  dff _57383_ (\oc8051_top_1.oc8051_decoder1.op [6], _28186_[6], clk);
  dff _57384_ (\oc8051_top_1.oc8051_decoder1.op [7], _28186_[7], clk);
  dff _57385_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _28187_, clk);
  dff _57386_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _28188_[0], clk);
  dff _57387_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _28188_[1], clk);
  dff _57388_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _28189_[0], clk);
  dff _57389_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _28189_[1], clk);
  dff _57390_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _28190_[0], clk);
  dff _57391_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _28190_[1], clk);
  dff _57392_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _28190_[2], clk);
  dff _57393_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _28191_[0], clk);
  dff _57394_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _28191_[1], clk);
  dff _57395_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _28191_[2], clk);
  dff _57396_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _28192_[0], clk);
  dff _57397_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _28192_[1], clk);
  dff _57398_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _28193_[0], clk);
  dff _57399_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _28193_[1], clk);
  dff _57400_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _28193_[2], clk);
  dff _57401_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _28193_[3], clk);
  dff _57402_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _28194_[0], clk);
  dff _57403_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _28194_[1], clk);
  dff _57404_ (\oc8051_top_1.oc8051_decoder1.wr , _28195_, clk);
  dff _57405_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _28234_, clk);
  dff _57406_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _28196_[0], clk);
  dff _57407_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _28196_[1], clk);
  dff _57408_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _28196_[2], clk);
  dff _57409_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _28196_[3], clk);
  dff _57410_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _28196_[4], clk);
  dff _57411_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _28196_[5], clk);
  dff _57412_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _28196_[6], clk);
  dff _57413_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _28196_[7], clk);
  dff _57414_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _28197_[0], clk);
  dff _57415_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _28197_[1], clk);
  dff _57416_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _28197_[2], clk);
  dff _57417_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _28197_[3], clk);
  dff _57418_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _28197_[4], clk);
  dff _57419_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _28197_[5], clk);
  dff _57420_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _28197_[6], clk);
  dff _57421_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _28197_[7], clk);
  dff _57422_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _28198_[0], clk);
  dff _57423_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _28198_[1], clk);
  dff _57424_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _28198_[2], clk);
  dff _57425_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _28198_[3], clk);
  dff _57426_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _28198_[4], clk);
  dff _57427_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _28198_[5], clk);
  dff _57428_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _28198_[6], clk);
  dff _57429_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _28198_[7], clk);
  dff _57430_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _28199_[0], clk);
  dff _57431_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _28199_[1], clk);
  dff _57432_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _28199_[2], clk);
  dff _57433_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _28199_[3], clk);
  dff _57434_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _28199_[4], clk);
  dff _57435_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _28199_[5], clk);
  dff _57436_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _28199_[6], clk);
  dff _57437_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _28199_[7], clk);
  dff _57438_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _28200_[0], clk);
  dff _57439_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _28200_[1], clk);
  dff _57440_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _28200_[2], clk);
  dff _57441_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _28200_[3], clk);
  dff _57442_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _28200_[4], clk);
  dff _57443_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _28200_[5], clk);
  dff _57444_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _28200_[6], clk);
  dff _57445_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _28200_[7], clk);
  dff _57446_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _28201_[0], clk);
  dff _57447_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _28201_[1], clk);
  dff _57448_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _28201_[2], clk);
  dff _57449_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _28201_[3], clk);
  dff _57450_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _28201_[4], clk);
  dff _57451_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _28201_[5], clk);
  dff _57452_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _28201_[6], clk);
  dff _57453_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _28201_[7], clk);
  dff _57454_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _28202_[0], clk);
  dff _57455_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _28202_[1], clk);
  dff _57456_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _28202_[2], clk);
  dff _57457_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _28202_[3], clk);
  dff _57458_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _28202_[4], clk);
  dff _57459_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _28202_[5], clk);
  dff _57460_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _28202_[6], clk);
  dff _57461_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _28202_[7], clk);
  dff _57462_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _28203_[0], clk);
  dff _57463_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _28203_[1], clk);
  dff _57464_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _28203_[2], clk);
  dff _57465_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _28203_[3], clk);
  dff _57466_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _28203_[4], clk);
  dff _57467_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _28203_[5], clk);
  dff _57468_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _28203_[6], clk);
  dff _57469_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _28203_[7], clk);
  dff _57470_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _28207_[0], clk);
  dff _57471_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _28207_[1], clk);
  dff _57472_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _28207_[2], clk);
  dff _57473_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _28207_[3], clk);
  dff _57474_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _28207_[4], clk);
  dff _57475_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _28204_[0], clk);
  dff _57476_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _28204_[1], clk);
  dff _57477_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _28204_[2], clk);
  dff _57478_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _28204_[3], clk);
  dff _57479_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _28204_[4], clk);
  dff _57480_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _28204_[5], clk);
  dff _57481_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _28204_[6], clk);
  dff _57482_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _28204_[7], clk);
  dff _57483_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _28204_[8], clk);
  dff _57484_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _28204_[9], clk);
  dff _57485_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _28204_[10], clk);
  dff _57486_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _28204_[11], clk);
  dff _57487_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _28204_[12], clk);
  dff _57488_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _28204_[13], clk);
  dff _57489_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _28204_[14], clk);
  dff _57490_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _28204_[15], clk);
  dff _57491_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _28205_[0], clk);
  dff _57492_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _28205_[1], clk);
  dff _57493_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _28205_[2], clk);
  dff _57494_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _28205_[3], clk);
  dff _57495_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _28205_[4], clk);
  dff _57496_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _28205_[5], clk);
  dff _57497_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _28205_[6], clk);
  dff _57498_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _28205_[7], clk);
  dff _57499_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _28205_[8], clk);
  dff _57500_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _28205_[9], clk);
  dff _57501_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _28205_[10], clk);
  dff _57502_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _28205_[11], clk);
  dff _57503_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _28205_[12], clk);
  dff _57504_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _28205_[13], clk);
  dff _57505_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _28205_[14], clk);
  dff _57506_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _28205_[15], clk);
  dff _57507_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _28225_[0], clk);
  dff _57508_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _28225_[1], clk);
  dff _57509_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _28225_[2], clk);
  dff _57510_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _28225_[3], clk);
  dff _57511_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _28225_[4], clk);
  dff _57512_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _28225_[5], clk);
  dff _57513_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _28225_[6], clk);
  dff _57514_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _28225_[7], clk);
  dff _57515_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _28225_[8], clk);
  dff _57516_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _28225_[9], clk);
  dff _57517_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _28225_[10], clk);
  dff _57518_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _28225_[11], clk);
  dff _57519_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _28225_[12], clk);
  dff _57520_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _28225_[13], clk);
  dff _57521_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _28225_[14], clk);
  dff _57522_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _28225_[15], clk);
  dff _57523_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _28225_[16], clk);
  dff _57524_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _28225_[17], clk);
  dff _57525_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _28225_[18], clk);
  dff _57526_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _28225_[19], clk);
  dff _57527_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _28225_[20], clk);
  dff _57528_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _28225_[21], clk);
  dff _57529_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _28225_[22], clk);
  dff _57530_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _28225_[23], clk);
  dff _57531_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _28225_[24], clk);
  dff _57532_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _28225_[25], clk);
  dff _57533_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _28225_[26], clk);
  dff _57534_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _28225_[27], clk);
  dff _57535_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _28225_[28], clk);
  dff _57536_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _28225_[29], clk);
  dff _57537_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _28225_[30], clk);
  dff _57538_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _28225_[31], clk);
  dff _57539_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _28206_, clk);
  dff _57540_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _28208_[0], clk);
  dff _57541_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _28208_[1], clk);
  dff _57542_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _28208_[2], clk);
  dff _57543_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _28208_[3], clk);
  dff _57544_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _28208_[4], clk);
  dff _57545_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _28208_[5], clk);
  dff _57546_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _28208_[6], clk);
  dff _57547_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _28208_[7], clk);
  dff _57548_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _28209_, clk);
  dff _57549_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _28210_, clk);
  dff _57550_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _28211_[0], clk);
  dff _57551_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _28211_[1], clk);
  dff _57552_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _28211_[2], clk);
  dff _57553_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _28211_[3], clk);
  dff _57554_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _28211_[4], clk);
  dff _57555_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _28211_[5], clk);
  dff _57556_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _28211_[6], clk);
  dff _57557_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _28211_[7], clk);
  dff _57558_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _28211_[8], clk);
  dff _57559_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _28211_[9], clk);
  dff _57560_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _28211_[10], clk);
  dff _57561_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _28211_[11], clk);
  dff _57562_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _28211_[12], clk);
  dff _57563_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _28211_[13], clk);
  dff _57564_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _28211_[14], clk);
  dff _57565_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _28211_[15], clk);
  dff _57566_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _28212_[0], clk);
  dff _57567_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _28212_[1], clk);
  dff _57568_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _28212_[2], clk);
  dff _57569_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _28212_[3], clk);
  dff _57570_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _28212_[4], clk);
  dff _57571_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _28212_[5], clk);
  dff _57572_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _28212_[6], clk);
  dff _57573_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _28212_[7], clk);
  dff _57574_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _28212_[8], clk);
  dff _57575_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _28212_[9], clk);
  dff _57576_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _28212_[10], clk);
  dff _57577_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _28212_[11], clk);
  dff _57578_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _28212_[12], clk);
  dff _57579_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _28212_[13], clk);
  dff _57580_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _28212_[14], clk);
  dff _57581_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _28212_[15], clk);
  dff _57582_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _28213_, clk);
  dff _57583_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _28215_, clk);
  dff _57584_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _28214_, clk);
  dff _57585_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _28216_[0], clk);
  dff _57586_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _28216_[1], clk);
  dff _57587_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _28216_[2], clk);
  dff _57588_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _28216_[3], clk);
  dff _57589_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _28216_[4], clk);
  dff _57590_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _28216_[5], clk);
  dff _57591_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _28216_[6], clk);
  dff _57592_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _28216_[7], clk);
  dff _57593_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _28217_[0], clk);
  dff _57594_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _28217_[1], clk);
  dff _57595_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _28217_[2], clk);
  dff _57596_ (\oc8051_top_1.oc8051_memory_interface1.reti , _28220_, clk);
  dff _57597_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _28221_[0], clk);
  dff _57598_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _28221_[1], clk);
  dff _57599_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _28221_[2], clk);
  dff _57600_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _28221_[3], clk);
  dff _57601_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _28221_[4], clk);
  dff _57602_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _28221_[5], clk);
  dff _57603_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _28221_[6], clk);
  dff _57604_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _28221_[7], clk);
  dff _57605_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _28222_, clk);
  dff _57606_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _28223_, clk);
  dff _57607_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _28224_[0], clk);
  dff _57608_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _28224_[1], clk);
  dff _57609_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _28224_[2], clk);
  dff _57610_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _28224_[3], clk);
  dff _57611_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _28226_[0], clk);
  dff _57612_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _28226_[1], clk);
  dff _57613_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _28226_[2], clk);
  dff _57614_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _28226_[3], clk);
  dff _57615_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _28226_[4], clk);
  dff _57616_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _28226_[5], clk);
  dff _57617_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _28226_[6], clk);
  dff _57618_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _28226_[7], clk);
  dff _57619_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _28226_[8], clk);
  dff _57620_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _28226_[9], clk);
  dff _57621_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _28226_[10], clk);
  dff _57622_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _28226_[11], clk);
  dff _57623_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _28226_[12], clk);
  dff _57624_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _28226_[13], clk);
  dff _57625_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _28226_[14], clk);
  dff _57626_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _28226_[15], clk);
  dff _57627_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _28226_[16], clk);
  dff _57628_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _28226_[17], clk);
  dff _57629_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _28226_[18], clk);
  dff _57630_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _28226_[19], clk);
  dff _57631_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _28226_[20], clk);
  dff _57632_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _28226_[21], clk);
  dff _57633_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _28226_[22], clk);
  dff _57634_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _28226_[23], clk);
  dff _57635_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _28226_[24], clk);
  dff _57636_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _28226_[25], clk);
  dff _57637_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _28226_[26], clk);
  dff _57638_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _28226_[27], clk);
  dff _57639_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _28226_[28], clk);
  dff _57640_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _28226_[29], clk);
  dff _57641_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _28226_[30], clk);
  dff _57642_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _28226_[31], clk);
  dff _57643_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _28227_, clk);
  dff _57644_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _28228_, clk);
  dff _57645_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _28229_, clk);
  dff _57646_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _28230_[0], clk);
  dff _57647_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _28230_[1], clk);
  dff _57648_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _28230_[2], clk);
  dff _57649_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _28230_[3], clk);
  dff _57650_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _28231_, clk);
  dff _57651_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _28232_, clk);
  dff _57652_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _28233_[0], clk);
  dff _57653_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _28233_[1], clk);
  dff _57654_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _28233_[2], clk);
  dff _57655_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _28233_[3], clk);
  dff _57656_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _28233_[4], clk);
  dff _57657_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _28233_[5], clk);
  dff _57658_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _28233_[6], clk);
  dff _57659_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _28233_[7], clk);
  dff _57660_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _28235_[0], clk);
  dff _57661_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _28235_[1], clk);
  dff _57662_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _28235_[2], clk);
  dff _57663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _05760_, clk);
  dff _57664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _05960_, clk);
  dff _57665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _28376_, clk);
  dff _57666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _05978_, clk);
  dff _57667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _05954_, clk);
  dff _57668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _05995_, clk);
  dff _57669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _08430_, clk);
  dff _57670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _06004_, clk);
  dff _57671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _06099_, clk);
  dff _57672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _06091_, clk);
  dff _57673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _06079_, clk);
  dff _57674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _08823_, clk);
  dff _57675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _09667_, clk);
  dff _57676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _08810_, clk);
  dff _57677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03245_, clk);
  dff _57678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _05758_, clk);
  dff _57679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _23830_, clk);
  dff _57680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _01451_, clk);
  dff _57681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _23831_, clk);
  dff _57682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _12130_, clk);
  dff _57683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _23832_, clk);
  dff _57684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _01449_, clk);
  dff _57685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _23833_, clk);
  dff _57686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _23848_, clk);
  dff _57687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _23826_, clk);
  dff _57688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _01458_, clk);
  dff _57689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _01805_, clk);
  dff _57690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _23827_, clk);
  dff _57691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _28281_, clk);
  dff _57692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _23828_, clk);
  dff _57693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _01455_, clk);
  dff _57694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _23829_, clk);
  dff _57695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _11651_, clk);
  dff _57696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _23819_, clk);
  dff _57697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _01469_, clk);
  dff _57698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _23821_, clk);
  dff _57699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _11103_, clk);
  dff _57700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _23822_, clk);
  dff _57701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _01466_, clk);
  dff _57702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _23824_, clk);
  dff _57703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _08743_, clk);
  dff _57704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _08268_, clk);
  dff _57705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _28325_, clk);
  dff _57706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _09898_, clk);
  dff _57707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _10730_, clk);
  dff _57708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _09900_, clk);
  dff _57709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _10065_, clk);
  dff _57710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _01755_, clk);
  dff _57711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _10079_, clk);
  dff _57712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _24596_, clk);
  dff _57713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _11369_, clk);
  dff _57714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _06729_, clk);
  dff _57715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _06008_, clk);
  dff _57716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _09060_, clk);
  dff _57717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _11365_, clk);
  dff _57718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _10210_, clk);
  dff _57719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _10080_, clk);
  dff _57720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _28324_, clk);
  dff _57721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _11645_, clk);
  dff _57722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _11292_, clk);
  dff _57723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _11362_, clk);
  dff _57724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _09009_, clk);
  dff _57725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _09014_, clk);
  dff _57726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _09011_, clk);
  dff _57727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _11332_, clk);
  dff _57728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _08675_, clk);
  dff _57729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _11330_, clk);
  dff _57730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _28321_, clk);
  dff _57731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _09050_, clk);
  dff _57732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _28322_, clk);
  dff _57733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _28323_, clk);
  dff _57734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _08826_, clk);
  dff _57735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _28318_, clk);
  dff _57736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _28319_, clk);
  dff _57737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _28320_, clk);
  dff _57738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _08621_, clk);
  dff _57739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _08628_, clk);
  dff _57740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _08701_, clk);
  dff _57741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _08703_, clk);
  dff _57742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _08706_, clk);
  dff _57743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _11302_, clk);
  dff _57744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _08589_, clk);
  dff _57745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _08591_, clk);
  dff _57746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _08601_, clk);
  dff _57747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _11313_, clk);
  dff _57748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _28317_, clk);
  dff _57749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _08578_, clk);
  dff _57750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _08646_, clk);
  dff _57751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _08446_, clk);
  dff _57752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _08303_, clk);
  dff _57753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _08322_, clk);
  dff _57754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _08350_, clk);
  dff _57755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _10083_, clk);
  dff _57756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _08514_, clk);
  dff _57757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _08535_, clk);
  dff _57758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _08484_, clk);
  dff _57759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _24341_, clk);
  dff _57760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _10086_, clk);
  dff _57761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _00673_, clk);
  dff _57762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _00700_, clk);
  dff _57763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _00560_, clk);
  dff _57764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _00569_, clk);
  dff _57765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _28316_, clk);
  dff _57766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _10221_, clk);
  dff _57767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _10153_, clk);
  dff _57768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _14775_, clk);
  dff _57769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _11077_, clk);
  dff _57770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _11074_, clk);
  dff _57771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _10261_, clk);
  dff _57772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _24662_, clk);
  dff _57773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _27162_, clk);
  dff _57774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _11272_, clk);
  dff _57775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _11043_, clk);
  dff _57776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _16923_, clk);
  dff _57777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _11041_, clk);
  dff _57778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _11053_, clk);
  dff _57779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _16163_, clk);
  dff _57780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _16092_, clk);
  dff _57781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _10155_, clk);
  dff _57782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _15340_, clk);
  dff _57783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _10164_, clk);
  dff _57784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _11036_, clk);
  dff _57785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _17272_, clk);
  dff _57786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _10159_, clk);
  dff _57787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _18400_, clk);
  dff _57788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _18361_, clk);
  dff _57789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _11013_, clk);
  dff _57790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _18635_, clk);
  dff _57791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _21036_, clk);
  dff _57792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _11707_, clk);
  dff _57793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _20873_, clk);
  dff _57794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _21572_, clk);
  dff _57795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _21268_, clk);
  dff _57796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _11768_, clk);
  dff _57797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _21283_, clk);
  dff _57798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _28367_, clk);
  dff _57799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _11740_, clk);
  dff _57800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _11723_, clk);
  dff _57801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _19311_, clk);
  dff _57802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _28366_, clk);
  dff _57803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _19422_, clk);
  dff _57804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _19021_, clk);
  dff _57805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _21623_, clk);
  dff _57806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _21000_, clk);
  dff _57807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _11817_, clk);
  dff _57808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _11819_, clk);
  dff _57809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _21130_, clk);
  dff _57810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _11656_, clk);
  dff _57811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _11689_, clk);
  dff _57812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _11655_, clk);
  dff _57813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _11725_, clk);
  dff _57814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _11727_, clk);
  dff _57815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _11563_, clk);
  dff _57816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _10924_, clk);
  dff _57817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _11567_, clk);
  dff _57818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _11580_, clk);
  dff _57819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _10792_, clk);
  dff _57820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _10972_, clk);
  dff _57821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _11833_, clk);
  dff _57822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _11860_, clk);
  dff _57823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _11525_, clk);
  dff _57824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _10807_, clk);
  dff _57825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _11529_, clk);
  dff _57826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _28365_, clk);
  dff _57827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _11539_, clk);
  dff _57828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _11553_, clk);
  dff _57829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _10799_, clk);
  dff _57830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _11559_, clk);
  dff _57831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _11478_, clk);
  dff _57832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _11495_, clk);
  dff _57833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _10930_, clk);
  dff _57834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _11499_, clk);
  dff _57835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _11507_, clk);
  dff _57836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _11514_, clk);
  dff _57837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _11521_, clk);
  dff _57838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _10810_, clk);
  dff _57839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _10938_, clk);
  dff _57840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _28363_, clk);
  dff _57841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _11453_, clk);
  dff _57842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _10832_, clk);
  dff _57843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _10981_, clk);
  dff _57844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _11463_, clk);
  dff _57845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _10829_, clk);
  dff _57846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _28364_, clk);
  dff _57847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _11364_, clk);
  dff _57848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _10941_, clk);
  dff _57849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _11371_, clk);
  dff _57850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _28362_, clk);
  dff _57851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _10842_, clk);
  dff _57852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _10982_, clk);
  dff _57853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _11399_, clk);
  dff _57854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _11425_, clk);
  dff _57855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _17928_, clk);
  dff _57856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _06394_, clk);
  dff _57857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _06549_, clk);
  dff _57858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _08941_, clk);
  dff _57859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _23803_, clk);
  dff _57860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _09759_, clk);
  dff _57861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _24503_, clk);
  dff _57862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _27341_, clk);
  dff _57863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _09948_, clk);
  dff _57864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _19717_, clk);
  dff _57865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _08952_, clk);
  dff _57866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _24857_, clk);
  dff _57867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _09781_, clk);
  dff _57868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _26446_, clk);
  dff _57869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _12364_, clk);
  dff _57870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _08948_, clk);
  dff _57871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _09805_, clk);
  dff _57872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _27368_, clk);
  dff _57873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _08957_, clk);
  dff _57874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _09026_, clk);
  dff _57875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _09801_, clk);
  dff _57876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _07024_, clk);
  dff _57877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _10987_, clk);
  dff _57878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _28375_, clk);
  dff _57879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _10614_, clk);
  dff _57880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _08963_, clk);
  dff _57881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _01784_, clk);
  dff _57882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _08962_, clk);
  dff _57883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _09252_, clk);
  dff _57884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _09806_, clk);
  dff _57885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _22413_, clk);
  dff _57886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _26327_, clk);
  dff _57887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _27156_, clk);
  dff _57888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _27562_, clk);
  dff _57889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _28237_, clk);
  dff _57890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _26617_, clk);
  dff _57891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _28238_, clk);
  dff _57892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _24967_, clk);
  dff _57893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _09062_, clk);
  dff _57894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _28239_, clk);
  dff _57895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _07458_, clk);
  dff _57896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _23654_, clk);
  dff _57897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _23868_, clk);
  dff _57898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _03196_, clk);
  dff _57899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _07615_, clk);
  dff _57900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _10732_, clk);
  dff _57901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _10670_, clk);
  dff _57902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _11193_, clk);
  dff _57903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _07360_, clk);
  dff _57904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _28242_, clk);
  dff _57905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _09024_, clk);
  dff _57906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _08626_, clk);
  dff _57907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _07358_, clk);
  dff _57908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _09887_, clk);
  dff _57909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _07613_, clk);
  dff _57910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _11262_, clk);
  dff _57911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _04284_, clk);
  dff _57912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _07604_, clk);
  dff _57913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _12111_, clk);
  dff _57914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _07430_, clk);
  dff _57915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _07380_, clk);
  dff _57916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _08497_, clk);
  dff _57917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _08507_, clk);
  dff _57918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _08377_, clk);
  dff _57919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _06085_, clk);
  dff _57920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _06071_, clk);
  dff _57921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _06151_, clk);
  dff _57922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _06174_, clk);
  dff _57923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _06158_, clk);
  dff _57924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _03212_, clk);
  dff _57925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _05755_, clk);
  dff _57926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _05804_, clk);
  dff _57927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _06326_, clk);
  dff _57928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _06298_, clk);
  dff _57929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _03202_, clk);
  dff _57930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _06444_, clk);
  dff _57931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _06423_, clk);
  dff _57932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _03161_, clk);
  dff _57933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _02340_, clk);
  dff _57934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _06069_, clk);
  dff _57935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _06933_, clk);
  dff _57936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _02157_, clk);
  dff _57937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _06531_, clk);
  dff _57938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _06508_, clk);
  dff _57939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _03144_, clk);
  dff _57940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _06595_, clk);
  dff _57941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _06591_, clk);
  dff _57942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _03143_, clk);
  dff _57943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _03133_, clk);
  dff _57944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _07125_, clk);
  dff _57945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _07094_, clk);
  dff _57946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _03129_, clk);
  dff _57947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _06884_, clk);
  dff _57948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _06866_, clk);
  dff _57949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _06831_, clk);
  dff _57950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _06942_, clk);
  dff _57951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _28311_, clk);
  dff _57952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _07272_, clk);
  dff _57953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _07278_, clk);
  dff _57954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _02171_, clk);
  dff _57955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _02440_, clk);
  dff _57956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _02496_, clk);
  dff _57957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _07026_, clk);
  dff _57958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _07018_, clk);
  dff _57959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _03102_, clk);
  dff _57960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _02345_, clk);
  dff _57961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _07397_, clk);
  dff _57962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _28310_, clk);
  dff _57963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _03118_, clk);
  dff _57964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _07479_, clk);
  dff _57965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _02175_, clk);
  dff _57966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _07187_, clk);
  dff _57967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _03096_, clk);
  dff _57968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _07737_, clk);
  dff _57969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _07786_, clk);
  dff _57970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _07759_, clk);
  dff _57971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _02180_, clk);
  dff _57972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _07532_, clk);
  dff _57973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _07523_, clk);
  dff _57974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _07611_, clk);
  dff _57975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _03087_, clk);
  dff _57976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _08098_, clk);
  dff _57977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _08093_, clk);
  dff _57978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _03084_, clk);
  dff _57979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _02349_, clk);
  dff _57980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _07697_, clk);
  dff _57981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _28309_, clk);
  dff _57982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _07678_, clk);
  dff _57983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _10757_, clk);
  dff _57984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _11154_, clk);
  dff _57985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _28335_, clk);
  dff _57986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _10727_, clk);
  dff _57987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _28336_, clk);
  dff _57988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _11208_, clk);
  dff _57989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _10536_, clk);
  dff _57990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _11221_, clk);
  dff _57991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _08897_, clk);
  dff _57992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _03078_, clk);
  dff _57993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _09081_, clk);
  dff _57994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _28307_, clk);
  dff _57995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _09089_, clk);
  dff _57996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _02193_, clk);
  dff _57997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _28308_, clk);
  dff _57998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _07847_, clk);
  dff _57999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _09114_, clk);
  dff _58000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _09742_, clk);
  dff _58001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _09980_, clk);
  dff _58002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _10151_, clk);
  dff _58003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _10088_, clk);
  dff _58004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _28306_, clk);
  dff _58005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _02198_, clk);
  dff _58006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _08895_, clk);
  dff _58007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _10401_, clk);
  dff _58008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _28303_, clk);
  dff _58009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _10367_, clk);
  dff _58010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _10344_, clk);
  dff _58011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _10914_, clk);
  dff _58012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _10825_, clk);
  dff _58013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _28304_, clk);
  dff _58014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _28305_, clk);
  dff _58015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _02209_, clk);
  dff _58016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _11024_, clk);
  dff _58017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _28302_, clk);
  dff _58018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _11183_, clk);
  dff _58019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _11181_, clk);
  dff _58020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _11169_, clk);
  dff _58021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _03046_, clk);
  dff _58022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _02359_, clk);
  dff _58023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _11714_, clk);
  dff _58024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _03030_, clk);
  dff _58025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _02363_, clk);
  dff _58026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _11240_, clk);
  dff _58027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _11270_, clk);
  dff _58028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _28301_, clk);
  dff _58029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _03042_, clk);
  dff _58030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _11335_, clk);
  dff _58031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _03027_, clk);
  dff _58032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _12007_, clk);
  dff _58033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _11970_, clk);
  dff _58034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _02223_, clk);
  dff _58035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _11550_, clk);
  dff _58036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _28300_, clk);
  dff _58037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _11487_, clk);
  dff _58038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _11715_, clk);
  dff _58039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _12065_, clk);
  dff _58040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _28298_, clk);
  dff _58041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _12121_, clk);
  dff _58042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _28299_, clk);
  dff _58043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _02227_, clk);
  dff _58044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _02449_, clk);
  dff _58045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _11779_, clk);
  dff _58046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _11804_, clk);
  dff _58047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _06408_, clk);
  dff _58048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _02998_, clk);
  dff _58049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _02368_, clk);
  dff _58050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _01629_, clk);
  dff _58051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _03010_, clk);
  dff _58052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _06666_, clk);
  dff _58053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _25117_, clk);
  dff _58054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _03007_, clk);
  dff _58055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _11823_, clk);
  dff _58056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _11600_, clk);
  dff _58057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _02989_, clk);
  dff _58058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _01387_, clk);
  dff _58059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _02983_, clk);
  dff _58060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _08559_, clk);
  dff _58061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _23855_, clk);
  dff _58062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _03002_, clk);
  dff _58063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _02310_, clk);
  dff _58064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _26116_, clk);
  dff _58065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _02801_, clk);
  dff _58066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _02306_, clk);
  dff _58067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _01744_, clk);
  dff _58068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _02812_, clk);
  dff _58069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _02805_, clk);
  dff _58070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _02418_, clk);
  dff _58071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _02744_, clk);
  dff _58072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _02466_, clk);
  dff _58073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _02780_, clk);
  dff _58074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _17283_, clk);
  dff _58075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _02774_, clk);
  dff _58076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _06391_, clk);
  dff _58077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _24932_, clk);
  dff _58078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _24812_, clk);
  dff _58079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _02751_, clk);
  dff _58080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _23690_, clk);
  dff _58081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _23751_, clk);
  dff _58082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _02763_, clk);
  dff _58083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _02423_, clk);
  dff _58084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _01390_, clk);
  dff _58085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _01365_, clk);
  dff _58086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _01679_, clk);
  dff _58087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _01583_, clk);
  dff _58088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _01311_, clk);
  dff _58089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _27985_, clk);
  dff _58090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _02970_, clk);
  dff _58091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _02371_, clk);
  dff _58092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _02483_, clk);
  dff _58093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _27128_, clk);
  dff _58094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _01092_, clk);
  dff _58095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _22334_, clk);
  dff _58096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _22307_, clk);
  dff _58097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _22242_, clk);
  dff _58098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _11710_, clk);
  dff _58099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _20898_, clk);
  dff _58100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _11080_, clk);
  dff _58101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _11095_, clk);
  dff _58102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _10610_, clk);
  dff _58103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _10601_, clk);
  dff _58104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _11112_, clk);
  dff _58105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _11120_, clk);
  dff _58106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _11128_, clk);
  dff _58107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _10562_, clk);
  dff _58108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _11136_, clk);
  dff _58109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _10556_, clk);
  dff _58110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _11146_, clk);
  dff _58111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _08162_, clk);
  dff _58112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _07516_, clk);
  dff _58113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _09277_, clk);
  dff _58114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _28297_, clk);
  dff _58115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _09305_, clk);
  dff _58116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _02237_, clk);
  dff _58117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _11704_, clk);
  dff _58118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _06250_, clk);
  dff _58119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _08928_, clk);
  dff _58120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _02250_, clk);
  dff _58121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _25124_, clk);
  dff _58122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _08657_, clk);
  dff _58123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _02958_, clk);
  dff _58124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _02978_, clk);
  dff _58125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _02391_, clk);
  dff _58126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _02247_, clk);
  dff _58127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _24608_, clk);
  dff _58128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _25184_, clk);
  dff _58129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _11287_, clk);
  dff _58130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _02253_, clk);
  dff _58131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _07617_, clk);
  dff _58132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _06699_, clk);
  dff _58133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _06643_, clk);
  dff _58134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _09159_, clk);
  dff _58135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _02260_, clk);
  dff _58136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _26631_, clk);
  dff _58137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _01727_, clk);
  dff _58138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _09913_, clk);
  dff _58139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _02925_, clk);
  dff _58140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _28296_, clk);
  dff _58141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _10342_, clk);
  dff _58142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _09972_, clk);
  dff _58143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _02489_, clk);
  dff _58144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _28295_, clk);
  dff _58145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _08582_, clk);
  dff _58146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _08432_, clk);
  dff _58147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _02903_, clk);
  dff _58148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _10637_, clk);
  dff _58149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _11664_, clk);
  dff _58150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _08850_, clk);
  dff _58151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _02874_, clk);
  dff _58152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _02395_, clk);
  dff _58153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _27585_, clk);
  dff _58154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _02890_, clk);
  dff _58155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _02885_, clk);
  dff _58156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _02571_, clk);
  dff _58157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _02898_, clk);
  dff _58158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _23684_, clk);
  dff _58159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _22695_, clk);
  dff _58160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _22593_, clk);
  dff _58161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _11732_, clk);
  dff _58162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _23037_, clk);
  dff _58163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _23199_, clk);
  dff _58164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _23058_, clk);
  dff _58165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _11712_, clk);
  dff _58166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _21845_, clk);
  dff _58167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _11691_, clk);
  dff _58168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _19656_, clk);
  dff _58169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _19605_, clk);
  dff _58170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _19503_, clk);
  dff _58171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _11641_, clk);
  dff _58172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _23682_, clk);
  dff _58173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _23680_, clk);
  dff _58174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _22786_, clk);
  dff _58175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _11777_, clk);
  dff _58176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _23734_, clk);
  dff _58177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _23733_, clk);
  dff _58178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _11830_, clk);
  dff _58179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _23746_, clk);
  dff _58180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _23744_, clk);
  dff _58181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _11775_, clk);
  dff _58182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _23755_, clk);
  dff _58183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _23715_, clk);
  dff _58184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _11773_, clk);
  dff _58185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _23689_, clk);
  dff _58186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _23687_, clk);
  dff _58187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _11881_, clk);
  dff _58188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _23695_, clk);
  dff _58189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _23693_, clk);
  dff _58190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _23692_, clk);
  dff _58191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _24901_, clk);
  dff _58192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _24847_, clk);
  dff _58193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _11578_, clk);
  dff _58194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _28333_, clk);
  dff _58195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _10349_, clk);
  dff _58196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _23696_, clk);
  dff _58197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _28334_, clk);
  dff _58198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _23716_, clk);
  dff _58199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _24615_, clk);
  dff _58200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _24854_, clk);
  dff _58201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _24851_, clk);
  dff _58202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _24834_, clk);
  dff _58203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _24219_, clk);
  dff _58204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _24168_, clk);
  dff _58205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _24141_, clk);
  dff _58206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _24134_, clk);
  dff _58207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _10558_, clk);
  dff _58208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _01411_, clk);
  dff _58209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _11574_, clk);
  dff _58210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _23688_, clk);
  dff _58211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _23683_, clk);
  dff _58212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _09992_, clk);
  dff _58213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _11610_, clk);
  dff _58214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _10823_, clk);
  dff _58215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _25211_, clk);
  dff _58216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _01891_, clk);
  dff _58217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _28236_, clk);
  dff _58218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _24937_, clk);
  dff _58219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _24952_, clk);
  dff _58220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _24943_, clk);
  dff _58221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _25077_, clk);
  dff _58222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _25060_, clk);
  dff _58223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _06471_, clk);
  dff _58224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _06467_, clk);
  dff _58225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _08316_, clk);
  dff _58226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _06288_, clk);
  dff _58227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _06278_, clk);
  dff _58228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _06270_, clk);
  dff _58229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _06363_, clk);
  dff _58230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _06354_, clk);
  dff _58231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _28315_, clk);
  dff _58232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _23763_, clk);
  dff _58233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _23760_, clk);
  dff _58234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _23758_, clk);
  dff _58235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _24022_, clk);
  dff _58236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _24008_, clk);
  dff _58237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _11608_, clk);
  dff _58238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _06413_, clk);
  dff _58239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _09474_, clk);
  dff _58240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _05782_, clk);
  dff _58241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _05778_, clk);
  dff _58242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _05773_, clk);
  dff _58243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _06638_, clk);
  dff _58244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _09546_, clk);
  dff _58245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _06240_, clk);
  dff _58246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _06232_, clk);
  dff _58247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _05823_, clk);
  dff _58248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _05835_, clk);
  dff _58249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _08798_, clk);
  dff _58250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _05893_, clk);
  dff _58251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _05905_, clk);
  dff _58252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _05897_, clk);
  dff _58253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _06655_, clk);
  dff _58254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _05720_, clk);
  dff _58255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _08372_, clk);
  dff _58256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _06527_, clk);
  dff _58257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _06510_, clk);
  dff _58258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _08318_, clk);
  dff _58259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _06572_, clk);
  dff _58260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _06563_, clk);
  dff _58261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _08388_, clk);
  dff _58262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _03342_, clk);
  dff _58263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _06137_, clk);
  dff _58264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _06129_, clk);
  dff _58265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _06123_, clk);
  dff _58266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _06198_, clk);
  dff _58267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _06181_, clk);
  dff _58268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _06170_, clk);
  dff _58269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _09016_, clk);
  dff _58270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _06034_, clk);
  dff _58271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _07333_, clk);
  dff _58272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _07180_, clk);
  dff _58273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _02869_, clk);
  dff _58274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _07842_, clk);
  dff _58275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _28294_, clk);
  dff _58276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _04504_, clk);
  dff _58277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _04489_, clk);
  dff _58278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _02877_, clk);
  dff _58279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _11618_, clk);
  dff _58280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _11605_, clk);
  dff _58281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _02834_, clk);
  dff _58282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _28293_, clk);
  dff _58283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _02855_, clk);
  dff _58284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _10945_, clk);
  dff _58285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _02848_, clk);
  dff _58286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _02400_, clk);
  dff _58287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _01817_, clk);
  dff _58288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _01596_, clk);
  dff _58289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _02298_, clk);
  dff _58290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _11721_, clk);
  dff _58291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _12091_, clk);
  dff _58292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _02827_, clk);
  dff _58293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _02405_, clk);
  dff _58294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _11149_, clk);
  dff _58295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _10141_, clk);
  dff _58296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _04147_, clk);
  dff _58297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _10340_, clk);
  dff _58298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _10484_, clk);
  dff _58299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _03941_, clk);
  dff _58300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _04278_, clk);
  dff _58301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _04355_, clk);
  dff _58302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _01442_, clk);
  dff _58303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _03965_, clk);
  dff _58304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _09809_, clk);
  dff _58305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _04161_, clk);
  dff _58306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _09855_, clk);
  dff _58307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _28292_, clk);
  dff _58308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _03950_, clk);
  dff _58309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _04281_, clk);
  dff _58310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _10005_, clk);
  dff _58311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _28291_, clk);
  dff _58312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _09638_, clk);
  dff _58313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _03972_, clk);
  dff _58314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _09693_, clk);
  dff _58315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _03970_, clk);
  dff _58316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _09695_, clk);
  dff _58317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _04179_, clk);
  dff _58318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _04334_, clk);
  dff _58319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _04357_, clk);
  dff _58320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _09183_, clk);
  dff _58321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _09471_, clk);
  dff _58322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _03984_, clk);
  dff _58323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _28289_, clk);
  dff _58324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _03982_, clk);
  dff _58325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _28290_, clk);
  dff _58326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _04184_, clk);
  dff _58327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _04295_, clk);
  dff _58328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _09068_, clk);
  dff _58329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _09141_, clk);
  dff _58330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _03997_, clk);
  dff _58331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _09155_, clk);
  dff _58332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _03996_, clk);
  dff _58333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _28288_, clk);
  dff _58334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _04197_, clk);
  dff _58335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _04211_, clk);
  dff _58336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _04343_, clk);
  dff _58337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _08926_, clk);
  dff _58338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _08932_, clk);
  dff _58339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _04004_, clk);
  dff _58340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _08939_, clk);
  dff _58341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _04002_, clk);
  dff _58342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _08944_, clk);
  dff _58343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _28286_, clk);
  dff _58344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _04216_, clk);
  dff _58345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _28287_, clk);
  dff _58346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _04029_, clk);
  dff _58347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _08867_, clk);
  dff _58348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _04213_, clk);
  dff _58349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _08871_, clk);
  dff _58350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _08923_, clk);
  dff _58351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _03754_, clk);
  dff _58352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _04268_, clk);
  dff _58353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _04353_, clk);
  dff _58354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _08722_, clk);
  dff _58355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _04039_, clk);
  dff _58356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _08724_, clk);
  dff _58357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _04218_, clk);
  dff _58358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _08755_, clk);
  dff _58359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _04128_, clk);
  dff _58360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _03606_, clk);
  dff _58361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _04143_, clk);
  dff _58362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _03721_, clk);
  dff _58363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _04124_, clk);
  dff _58364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _03733_, clk);
  dff _58365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _04272_, clk);
  dff _58366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _03747_, clk);
  dff _58367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _04051_, clk);
  dff _58368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _08523_, clk);
  dff _58369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _04049_, clk);
  dff _58370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _08718_, clk);
  dff _58371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _04227_, clk);
  dff _58372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _04345_, clk);
  dff _58373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _03648_, clk);
  dff _58374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _04137_, clk);
  dff _58375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _06940_, clk);
  dff _58376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _04075_, clk);
  dff _58377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _07158_, clk);
  dff _58378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _04073_, clk);
  dff _58379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _07161_, clk);
  dff _58380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _04229_, clk);
  dff _58381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _08155_, clk);
  dff _58382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _04064_, clk);
  dff _58383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _06669_, clk);
  dff _58384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _06710_, clk);
  dff _58385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _04102_, clk);
  dff _58386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _06725_, clk);
  dff _58387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _04100_, clk);
  dff _58388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _06785_, clk);
  dff _58389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _04241_, clk);
  dff _58390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _04349_, clk);
  dff _58391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _04263_, clk);
  dff _58392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _04359_, clk);
  dff _58393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _06094_, clk);
  dff _58394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _04115_, clk);
  dff _58395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _06650_, clk);
  dff _58396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _04108_, clk);
  dff _58397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _06652_, clk);
  dff _58398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _04260_, clk);
  dff _58399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _04330_, clk);
  dff _58400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _04202_, clk);
  dff _58401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _04239_, clk);
  dff _58402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _06789_, clk);
  dff _58403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _04200_, clk);
  dff _58404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _04287_, clk);
  dff _58405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _04297_, clk);
  dff _58406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _06832_, clk);
  dff _58407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _03863_, clk);
  dff _58408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _06812_, clk);
  dff _58409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _06799_, clk);
  dff _58410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _06817_, clk);
  dff _58411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _04190_, clk);
  dff _58412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _03864_, clk);
  dff _58413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _03875_, clk);
  dff _58414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _06742_, clk);
  dff _58415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _06421_, clk);
  dff _58416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _06448_, clk);
  dff _58417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _04816_, clk);
  dff _58418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _06901_, clk);
  dff _58419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _06911_, clk);
  dff _58420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _06887_, clk);
  dff _58421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _06752_, clk);
  dff _58422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _06746_, clk);
  dff _58423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _06302_, clk);
  dff _58424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _06343_, clk);
  dff _58425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _06365_, clk);
  dff _58426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _04840_, clk);
  dff _58427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _06374_, clk);
  dff _58428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _05078_, clk);
  dff _58429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _06396_, clk);
  dff _58430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _06415_, clk);
  dff _58431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _05096_, clk);
  dff _58432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _06219_, clk);
  dff _58433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _06244_, clk);
  dff _58434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _04869_, clk);
  dff _58435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _06265_, clk);
  dff _58436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _04863_, clk);
  dff _58437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _06284_, clk);
  dff _58438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _05086_, clk);
  dff _58439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _04896_, clk);
  dff _58440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _06118_, clk);
  dff _58441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _05110_, clk);
  dff _58442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _06140_, clk);
  dff _58443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _06156_, clk);
  dff _58444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _05107_, clk);
  dff _58445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _06200_, clk);
  dff _58446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _06214_, clk);
  dff _58447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _05142_, clk);
  dff _58448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _06021_, clk);
  dff _58449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _06041_, clk);
  dff _58450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _04935_, clk);
  dff _58451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _05256_, clk);
  dff _58452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _06063_, clk);
  dff _58453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _06083_, clk);
  dff _58454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _04925_, clk);
  dff _58455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _05890_, clk);
  dff _58456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _05913_, clk);
  dff _58457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _05945_, clk);
  dff _58458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _04951_, clk);
  dff _58459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _05951_, clk);
  dff _58460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _05150_, clk);
  dff _58461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _05993_, clk);
  dff _58462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _06014_, clk);
  dff _58463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _05485_, clk);
  dff _58464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _05045_, clk);
  dff _58465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _05809_, clk);
  dff _58466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _05839_, clk);
  dff _58467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _04966_, clk);
  dff _58468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _05860_, clk);
  dff _58469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _05882_, clk);
  dff _58470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _04963_, clk);
  dff _58471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _05385_, clk);
  dff _58472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _05409_, clk);
  dff _58473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _05377_, clk);
  dff _58474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _05068_, clk);
  dff _58475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _05422_, clk);
  dff _58476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _05451_, clk);
  dff _58477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _05054_, clk);
  dff _58478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _05471_, clk);
  dff _58479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _05689_, clk);
  dff _58480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _05707_, clk);
  dff _58481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _05168_, clk);
  dff _58482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _05714_, clk);
  dff _58483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _05728_, clk);
  dff _58484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _05765_, clk);
  dff _58485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _05789_, clk);
  dff _58486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _04975_, clk);
  dff _58487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _05024_, clk);
  dff _58488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _05608_, clk);
  dff _58489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _05018_, clk);
  dff _58490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _05615_, clk);
  dff _58491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _05283_, clk);
  dff _58492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _05631_, clk);
  dff _58493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _05681_, clk);
  dff _58494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _04993_, clk);
  dff _58495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _05504_, clk);
  dff _58496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _05042_, clk);
  dff _58497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _05519_, clk);
  dff _58498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _05200_, clk);
  dff _58499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _05525_, clk);
  dff _58500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _05543_, clk);
  dff _58501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _05583_, clk);
  dff _58502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _05033_, clk);
  dff _58503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _06811_, clk);
  dff _58504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _04361_, clk);
  dff _58505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _04351_, clk);
  dff _58506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _04339_, clk);
  dff _58507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _04438_, clk);
  dff _58508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _04432_, clk);
  dff _58509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _04414_, clk);
  dff _58510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _06824_, clk);
  dff _58511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _03860_, clk);
  dff _58512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _04645_, clk);
  dff _58513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _06805_, clk);
  dff _58514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _04469_, clk);
  dff _58515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _04483_, clk);
  dff _58516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _04474_, clk);
  dff _58517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _06813_, clk);
  dff _58518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _04565_, clk);
  dff _58519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _04092_, clk);
  dff _58520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _06750_, clk);
  dff _58521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _03823_, clk);
  dff _58522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _03799_, clk);
  dff _58523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _03784_, clk);
  dff _58524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _03927_, clk);
  dff _58525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _03901_, clk);
  dff _58526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _03887_, clk);
  dff _58527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _06890_, clk);
  dff _58528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _05057_, clk);
  dff _58529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _05040_, clk);
  dff _58530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _05099_, clk);
  dff _58531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _03993_, clk);
  dff _58532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _04010_, clk);
  dff _58533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _06754_, clk);
  dff _58534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _04077_, clk);
  dff _58535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _04709_, clk);
  dff _58536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _04691_, clk);
  dff _58537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _06918_, clk);
  dff _58538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _04798_, clk);
  dff _58539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _04765_, clk);
  dff _58540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _04758_, clk);
  dff _58541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _04987_, clk);
  dff _58542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _04981_, clk);
  dff _58543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _10744_, clk);
  dff _58544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _10521_, clk);
  dff _58545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _04368_, clk);
  dff _58546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _04857_, clk);
  dff _58547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _04846_, clk);
  dff _58548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _04943_, clk);
  dff _58549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _04938_, clk);
  dff _58550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _04918_, clk);
  dff _58551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _03963_, clk);
  dff _58552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _03435_, clk);
  dff _58553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _03622_, clk);
  dff _58554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _03610_, clk);
  dff _58555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _03452_, clk);
  dff _58556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _03723_, clk);
  dff _58557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _03683_, clk);
  dff _58558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _03448_, clk);
  dff _58559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _11620_, clk);
  dff _58560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _11613_, clk);
  dff _58561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _28285_, clk);
  dff _58562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _11115_, clk);
  dff _58563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _06424_, clk);
  dff _58564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _02275_, clk);
  dff _58565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _02634_, clk);
  dff _58566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _06455_, clk);
  dff _58567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _11866_, clk);
  dff _58568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _06399_, clk);
  dff _58569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _25221_, clk);
  dff _58570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _24526_, clk);
  dff _58571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _03802_, clk);
  dff _58572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _03745_, clk);
  dff _58573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _02315_, clk);
  dff _58574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _04374_, clk);
  dff _58575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _24880_, clk);
  dff _58576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _28284_, clk);
  dff _58577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _09066_, clk);
  dff _58578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _06380_, clk);
  dff _58579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _04582_, clk);
  dff _58580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _08330_, clk);
  dff _58581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _07425_, clk);
  dff _58582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _06410_, clk);
  dff _58583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _09039_, clk);
  dff _58584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _09020_, clk);
  dff _58585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _08832_, clk);
  dff _58586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _08846_, clk);
  dff _58587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _08855_, clk);
  dff _58588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _04381_, clk);
  dff _58589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _10898_, clk);
  dff _58590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _09683_, clk);
  dff _58591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _08586_, clk);
  dff _58592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _08598_, clk);
  dff _58593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _04388_, clk);
  dff _58594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _28282_, clk);
  dff _58595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _08689_, clk);
  dff _58596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _08704_, clk);
  dff _58597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _28283_, clk);
  dff _58598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _08662_, clk);
  dff _58599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _08488_, clk);
  dff _58600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _08493_, clk);
  dff _58601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _08495_, clk);
  dff _58602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _04404_, clk);
  dff _58603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _04688_, clk);
  dff _58604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _08634_, clk);
  dff _58605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _08632_, clk);
  dff _58606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _06330_, clk);
  dff _58607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _06275_, clk);
  dff _58608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _00907_, clk);
  dff _58609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _08288_, clk);
  dff _58610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _08292_, clk);
  dff _58611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _04406_, clk);
  dff _58612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _08555_, clk);
  dff _58613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _08539_, clk);
  dff _58614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _08553_, clk);
  dff _58615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _00574_, clk);
  dff _58616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _00605_, clk);
  dff _58617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _27170_, clk);
  dff _58618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _24660_, clk);
  dff _58619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _24800_, clk);
  dff _58620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _04408_, clk);
  dff _58621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _08364_, clk);
  dff _58622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _28280_, clk);
  dff _58623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _03425_, clk);
  dff _58624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _03885_, clk);
  dff _58625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _07384_, clk);
  dff _58626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _23707_, clk);
  dff _58627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _27821_, clk);
  dff _58628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _27588_, clk);
  dff _58629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _07382_, clk);
  dff _58630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _07845_, clk);
  dff _58631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _28374_, clk);
  dff _58632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _09926_, clk);
  dff _58633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _03594_, clk);
  dff _58634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _08969_, clk);
  dff _58635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _09902_, clk);
  dff _58636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _04674_, clk);
  dff _58637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _10112_, clk);
  dff _58638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _08965_, clk);
  dff _58639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _10861_, clk);
  dff _58640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _11315_, clk);
  dff _58641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _10943_, clk);
  dff _58642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _11324_, clk);
  dff _58643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _11340_, clk);
  dff _58644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _10854_, clk);
  dff _58645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _11001_, clk);
  dff _58646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _11355_, clk);
  dff _58647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _11266_, clk);
  dff _58648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _10885_, clk);
  dff _58649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _11274_, clk);
  dff _58650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _10947_, clk);
  dff _58651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _11294_, clk);
  dff _58652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _28361_, clk);
  dff _58653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _10869_, clk);
  dff _58654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _10985_, clk);
  dff _58655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _10993_, clk);
  dff _58656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _28359_, clk);
  dff _58657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _11052_, clk);
  dff _58658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _10919_, clk);
  dff _58659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _28360_, clk);
  dff _58660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _10917_, clk);
  dff _58661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _11070_, clk);
  dff _58662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _10968_, clk);
  dff _58663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _28356_, clk);
  dff _58664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _11212_, clk);
  dff _58665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _11223_, clk);
  dff _58666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _28357_, clk);
  dff _58667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _28358_, clk);
  dff _58668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _11022_, clk);
  dff _58669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _11032_, clk);
  dff _58670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _10921_, clk);
  dff _58671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _10900_, clk);
  dff _58672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _11142_, clk);
  dff _58673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _10963_, clk);
  dff _58674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _28353_, clk);
  dff _58675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _28354_, clk);
  dff _58676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _11173_, clk);
  dff _58677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _28355_, clk);
  dff _58678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _11189_, clk);
  dff _58679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _28350_, clk);
  dff _58680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _10908_, clk);
  dff _58681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _11099_, clk);
  dff _58682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _11110_, clk);
  dff _58683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _28351_, clk);
  dff _58684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _10904_, clk);
  dff _58685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _11123_, clk);
  dff _58686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _28352_, clk);
  dff _58687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _11653_, clk);
  dff _58688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _28348_, clk);
  dff _58689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _19097_, clk);
  dff _58690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _11730_, clk);
  dff _58691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _11717_, clk);
  dff _58692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _11743_, clk);
  dff _58693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _11719_, clk);
  dff _58694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _28349_, clk);
  dff _58695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _11576_, clk);
  dff _58696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _10660_, clk);
  dff _58697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _11847_, clk);
  dff _58698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _28346_, clk);
  dff _58699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _28347_, clk);
  dff _58700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _11808_, clk);
  dff _58701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _11821_, clk);
  dff _58702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _21091_, clk);
  dff _58703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _10361_, clk);
  dff _58704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _11546_, clk);
  dff _58705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _11555_, clk);
  dff _58706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _10358_, clk);
  dff _58707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _28344_, clk);
  dff _58708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _28345_, clk);
  dff _58709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _11561_, clk);
  dff _58710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _11569_, clk);
  dff _58711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _11509_, clk);
  dff _58712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _10373_, clk);
  dff _58713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _11515_, clk);
  dff _58714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _10371_, clk);
  dff _58715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _11519_, clk);
  dff _58716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _10678_, clk);
  dff _58717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _11527_, clk);
  dff _58718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _10364_, clk);
  dff _58719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _11459_, clk);
  dff _58720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _11472_, clk);
  dff _58721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _10385_, clk);
  dff _58722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _11481_, clk);
  dff _58723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _28343_, clk);
  dff _58724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _11489_, clk);
  dff _58725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _10685_, clk);
  dff _58726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _11504_, clk);
  dff _58727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _11403_, clk);
  dff _58728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _11428_, clk);
  dff _58729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _10393_, clk);
  dff _58730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _11442_, clk);
  dff _58731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _28342_, clk);
  dff _58732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _11451_, clk);
  dff _58733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _10691_, clk);
  dff _58734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _10773_, clk);
  dff _58735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _10413_, clk);
  dff _58736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _28341_, clk);
  dff _58737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _11367_, clk);
  dff _58738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _10407_, clk);
  dff _58739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _11377_, clk);
  dff _58740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _10405_, clk);
  dff _58741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _11380_, clk);
  dff _58742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _10695_, clk);
  dff _58743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _11277_, clk);
  dff _58744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _11298_, clk);
  dff _58745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _10513_, clk);
  dff _58746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _11300_, clk);
  dff _58747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _11308_, clk);
  dff _58748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _11321_, clk);
  dff _58749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _28340_, clk);
  dff _58750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _11328_, clk);
  dff _58751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _10766_, clk);
  dff _58752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _11039_, clk);
  dff _58753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _11047_, clk);
  dff _58754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _11066_, clk);
  dff _58755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _10634_, clk);
  dff _58756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _11072_, clk);
  dff _58757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _10739_, clk);
  dff _58758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _11268_, clk);
  dff _58759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _28337_, clk);
  dff _58760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _10724_, clk);
  dff _58761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _11231_, clk);
  dff _58762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _11252_, clk);
  dff _58763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _11026_, clk);
  dff _58764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _28338_, clk);
  dff _58765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _11030_, clk);
  dff _58766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _28339_, clk);
  dff _58767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _23854_, clk);
  dff _58768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _11257_, clk);
  dff _58769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _28058_, clk);
  dff _58770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _06262_, clk);
  dff _58771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _25328_, clk);
  dff _58772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _17786_, clk);
  dff _58773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _11028_, clk);
  dff _58774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _18055_, clk);
  dff _58775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _11838_, clk);
  dff _58776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _11422_, clk);
  dff _58777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _10199_, clk);
  dff _58778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _10143_, clk);
  dff _58779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _10128_, clk);
  dff _58780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _11444_, clk);
  dff _58781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _10587_, clk);
  dff _58782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _10056_, clk);
  dff _58783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _27475_, clk);
  dff _58784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _28314_, clk);
  dff _58785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _15309_, clk);
  dff _58786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _10954_, clk);
  dff _58787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _18261_, clk);
  dff _58788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _01289_, clk);
  dff _58789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _25041_, clk);
  dff _58790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _25429_, clk);
  dff _58791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _24487_, clk);
  dff _58792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _11417_, clk);
  dff _58793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _24233_, clk);
  dff _58794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _24875_, clk);
  dff _58795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _24238_, clk);
  dff _58796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _10061_, clk);
  dff _58797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _11592_, clk);
  dff _58798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _11420_, clk);
  dff _58799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _25142_, clk);
  dff _58800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _11890_, clk);
  dff _58801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _23823_, clk);
  dff _58802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _11218_, clk);
  dff _58803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _23863_, clk);
  dff _58804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _03574_, clk);
  dff _58805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _13886_, clk);
  dff _58806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _06965_, clk);
  dff _58807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _01736_, clk);
  dff _58808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _11396_, clk);
  dff _58809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _06722_, clk);
  dff _58810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _04921_, clk);
  dff _58811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _11384_, clk);
  dff _58812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _10208_, clk);
  dff _58813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _08550_, clk);
  dff _58814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _26316_, clk);
  dff _58815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _08762_, clk);
  dff _58816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _11617_, clk);
  dff _58817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _11210_, clk);
  dff _58818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _26479_, clk);
  dff _58819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _24781_, clk);
  dff _58820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _11203_, clk);
  dff _58821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _28313_, clk);
  dff _58822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _25105_, clk);
  dff _58823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _11187_, clk);
  dff _58824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _27422_, clk);
  dff _58825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _11171_, clk);
  dff _58826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _10227_, clk);
  dff _58827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _26321_, clk);
  dff _58828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _11196_, clk);
  dff _58829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _08600_, clk);
  dff _58830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _10094_, clk);
  dff _58831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _23481_, clk);
  dff _58832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _10118_, clk);
  dff _58833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _10301_, clk);
  dff _58834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _11244_, clk);
  dff _58835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _04164_, clk);
  dff _58836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _01876_, clk);
  dff _58837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _11157_, clk);
  dff _58838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _24101_, clk);
  dff _58839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _07035_, clk);
  dff _58840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _28312_, clk);
  dff _58841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _10229_, clk);
  dff _58842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _01627_, clk);
  dff _58843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _11140_, clk);
  dff _58844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _11133_, clk);
  dff _58845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _11709_, clk);
  dff _58846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _11832_, clk);
  dff _58847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _10239_, clk);
  dff _58848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _09544_, clk);
  dff _58849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _09479_, clk);
  dff _58850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _11121_, clk);
  dff _58851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _10448_, clk);
  dff _58852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _10271_, clk);
  dff _58853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _05983_, clk);
  dff _58854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _05881_, clk);
  dff _58855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _12491_, clk);
  dff _58856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _11108_, clk);
  dff _58857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _12718_, clk);
  dff _58858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _12867_, clk);
  dff _58859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _10136_, clk);
  dff _58860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _11178_, clk);
  dff _58861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _12057_, clk);
  dff _58862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _11868_, clk);
  dff _58863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _14118_, clk);
  dff _58864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _11090_, clk);
  dff _58865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _14393_, clk);
  dff _58866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _11082_, clk);
  dff _58867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _13278_, clk);
  dff _58868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _11097_, clk);
  dff _58869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _13632_, clk);
  dff _58870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _10139_, clk);
  dff _58871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _01586_, clk);
  dff _58872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _23867_, clk);
  dff _58873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _23869_, clk);
  dff _58874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _12087_, clk);
  dff _58875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _23930_, clk);
  dff _58876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _12082_, clk);
  dff _58877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _23947_, clk);
  dff _58878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _01581_, clk);
  dff _58879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _01446_, clk);
  dff _58880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _01802_, clk);
  dff _58881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _23849_, clk);
  dff _58882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _23857_, clk);
  dff _58883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _12113_, clk);
  dff _58884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _23860_, clk);
  dff _58885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _12106_, clk);
  dff _58886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _23866_, clk);
  dff _58887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _23552_, clk);
  dff _58888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _23815_, clk);
  dff _58889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _04983_, clk);
  dff _58890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _23816_, clk);
  dff _58891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _01472_, clk);
  dff _58892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _01807_, clk);
  dff _58893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _23817_, clk);
  dff _58894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _23818_, clk);
  dff _58895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _15959_, clk);
  dff _58896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _09829_, clk);
  dff _58897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _01439_, clk);
  dff _58898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _04506_, clk);
  dff _58899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _09072_, clk);
  dff _58900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _28370_, clk);
  dff _58901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _10845_, clk);
  dff _58902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _24720_, clk);
  dff _58903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _22462_, clk);
  dff _58904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _20174_, clk);
  dff _58905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _20109_, clk);
  dff _58906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _19987_, clk);
  dff _58907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _05923_, clk);
  dff _58908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _20458_, clk);
  dff _58909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _20605_, clk);
  dff _58910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _05916_, clk);
  dff _58911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _26128_, clk);
  dff _58912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _05687_, clk);
  dff _58913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _26219_, clk);
  dff _58914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _05677_, clk);
  dff _58915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _04641_, clk);
  dff _58916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _25878_, clk);
  dff _58917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _05694_, clk);
  dff _58918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _26022_, clk);
  dff _58919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _05626_, clk);
  dff _58920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _26516_, clk);
  dff _58921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _04501_, clk);
  dff _58922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _04741_, clk);
  dff _58923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _26280_, clk);
  dff _58924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _26297_, clk);
  dff _58925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _26336_, clk);
  dff _58926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _05647_, clk);
  dff _58927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _28268_, clk);
  dff _58928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _07319_, clk);
  dff _58929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _28269_, clk);
  dff _58930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _09077_, clk);
  dff _58931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _09110_, clk);
  dff _58932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _09106_, clk);
  dff _58933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _07317_, clk);
  dff _58934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _28270_, clk);
  dff _58935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _28271_, clk);
  dff _58936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _07311_, clk);
  dff _58937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _07705_, clk);
  dff _58938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _07687_, clk);
  dff _58939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _07684_, clk);
  dff _58940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _28272_, clk);
  dff _58941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _07784_, clk);
  dff _58942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _07770_, clk);
  dff _58943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _08752_, clk);
  dff _58944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _08748_, clk);
  dff _58945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _07772_, clk);
  dff _58946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _08899_, clk);
  dff _58947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _07314_, clk);
  dff _58948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _07820_, clk);
  dff _58949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _07815_, clk);
  dff _58950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _07792_, clk);
  dff _58951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _11159_, clk);
  dff _58952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _07681_, clk);
  dff _58953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _01227_, clk);
  dff _58954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _07680_, clk);
  dff _58955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _02944_, clk);
  dff _58956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _23796_, clk);
  dff _58957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _07688_, clk);
  dff _58958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _06956_, clk);
  dff _58959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _07343_, clk);
  dff _58960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _11161_, clk);
  dff _58961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _04519_, clk);
  dff _58962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _07676_, clk);
  dff _58963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _24879_, clk);
  dff _58964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _23753_, clk);
  dff _58965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _11326_, clk);
  dff _58966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _28253_, clk);
  dff _58967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _28368_, clk);
  dff _58968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _10976_, clk);
  dff _58969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _11106_, clk);
  dff _58970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _11238_, clk);
  dff _58971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _09095_, clk);
  dff _58972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _28369_, clk);
  dff _58973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _09831_, clk);
  dff _58974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _11532_, clk);
  dff _58975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _11117_, clk);
  dff _58976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _06757_, clk);
  dff _58977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _08978_, clk);
  dff _58978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _25302_, clk);
  dff _58979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _08976_, clk);
  dff _58980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _24841_, clk);
  dff _58981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _09820_, clk);
  dff _58982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _28371_, clk);
  dff _58983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _19973_, clk);
  dff _58984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _19921_, clk);
  dff _58985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _20409_, clk);
  dff _58986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _20330_, clk);
  dff _58987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _20263_, clk);
  dff _58988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _11667_, clk);
  dff _58989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _18879_, clk);
  dff _58990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _18851_, clk);
  dff _58991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _27440_, clk);
  dff _58992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _27343_, clk);
  dff _58993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _01189_, clk);
  dff _58994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _01417_, clk);
  dff _58995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _01244_, clk);
  dff _58996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _11501_, clk);
  dff _58997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _25064_, clk);
  dff _58998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _24291_, clk);
  dff _58999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _01623_, clk);
  dff _59000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _09997_, clk);
  dff _59001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _23740_, clk);
  dff _59002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _23713_, clk);
  dff _59003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _27428_, clk);
  dff _59004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _27364_, clk);
  dff _59005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _27165_, clk);
  dff _59006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _09995_, clk);
  dff _59007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _11557_, clk);
  dff _59008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _01897_, clk);
  dff _59009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _01886_, clk);
  dff _59010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _09999_, clk);
  dff _59011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _01273_, clk);
  dff _59012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _01139_, clk);
  dff _59013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _01122_, clk);
  dff _59014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _01656_, clk);
  dff _59015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _07690_, clk);
  dff _59016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _11552_, clk);
  dff _59017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _08335_, clk);
  dff _59018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _08530_, clk);
  dff _59019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _11548_, clk);
  dff _59020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _01798_, clk);
  dff _59021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _01721_, clk);
  dff _59022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _01708_, clk);
  dff _59023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _11523_, clk);
  dff _59024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _09263_, clk);
  dff _59025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _09261_, clk);
  dff _59026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _09239_, clk);
  dff _59027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _11536_, clk);
  dff _59028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _09350_, clk);
  dff _59029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _09360_, clk);
  dff _59030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _28332_, clk);
  dff _59031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _11780_, clk);
  dff _59032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _28331_, clk);
  dff _59033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _10269_, clk);
  dff _59034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _09428_, clk);
  dff _59035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _09419_, clk);
  dff _59036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _09413_, clk);
  dff _59037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _09691_, clk);
  dff _59038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _09578_, clk);
  dff _59039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _07701_, clk);
  dff _59040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _11317_, clk);
  dff _59041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _10018_, clk);
  dff _59042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _10618_, clk);
  dff _59043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _11614_, clk);
  dff _59044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _10647_, clk);
  dff _59045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _11885_, clk);
  dff _59046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _11851_, clk);
  dff _59047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _23793_, clk);
  dff _59048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _24974_, clk);
  dff _59049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _24107_, clk);
  dff _59050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _10020_, clk);
  dff _59051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _18983_, clk);
  dff _59052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _11164_, clk);
  dff _59053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _23752_, clk);
  dff _59054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _07788_, clk);
  dff _59055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _03167_, clk);
  dff _59056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _03159_, clk);
  dff _59057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _11497_, clk);
  dff _59058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _03663_, clk);
  dff _59059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _03608_, clk);
  dff _59060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _11493_, clk);
  dff _59061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _10194_, clk);
  dff _59062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _27257_, clk);
  dff _59063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _08726_, clk);
  dff _59064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _28330_, clk);
  dff _59065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _10039_, clk);
  dff _59066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _04032_, clk);
  dff _59067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _03922_, clk);
  dff _59068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _11483_, clk);
  dff _59069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _06707_, clk);
  dff _59070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _06702_, clk);
  dff _59071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _08869_, clk);
  dff _59072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _11466_, clk);
  dff _59073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _28329_, clk);
  dff _59074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _08980_, clk);
  dff _59075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _11461_, clk);
  dff _59076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _07520_, clk);
  dff _59077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _07267_, clk);
  dff _59078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _07199_, clk);
  dff _59079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _09457_, clk);
  dff _59080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _09266_, clk);
  dff _59081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _09636_, clk);
  dff _59082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _28326_, clk);
  dff _59083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _10052_, clk);
  dff _59084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _28327_, clk);
  dff _59085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _28328_, clk);
  dff _59086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _08893_, clk);
  dff _59087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _04838_, clk);
  dff _59088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _23810_, clk);
  dff _59089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _01478_, clk);
  dff _59090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _23811_, clk);
  dff _59091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _23813_, clk);
  dff _59092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _23812_, clk);
  dff _59093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _01610_, clk);
  dff _59094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _23814_, clk);
  dff _59095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _23804_, clk);
  dff _59096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _23769_, clk);
  dff _59097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _01359_, clk);
  dff _59098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _23770_, clk);
  dff _59099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _23771_, clk);
  dff _59100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _01235_, clk);
  dff _59101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _23772_, clk);
  dff _59102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _01579_, clk);
  dff _59103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _23797_, clk);
  dff _59104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03681_, clk);
  dff _59105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _23799_, clk);
  dff _59106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _01505_, clk);
  dff _59107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _23800_, clk);
  dff _59108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _11353_, clk);
  dff _59109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _23801_, clk);
  dff _59110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _01487_, clk);
  dff _59111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _23681_, clk);
  dff _59112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _23783_, clk);
  dff _59113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _23785_, clk);
  dff _59114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _25917_, clk);
  dff _59115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _23786_, clk);
  dff _59116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _01510_, clk);
  dff _59117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _23795_, clk);
  dff _59118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _25419_, clk);
  dff _59119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _28246_, clk);
  dff _59120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _23774_, clk);
  dff _59121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _23775_, clk);
  dff _59122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _01225_, clk);
  dff _59123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _23776_, clk);
  dff _59124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _01223_, clk);
  dff _59125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _23778_, clk);
  dff _59126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _01576_, clk);
  dff _59127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _04593_, clk);
  dff _59128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _23864_, clk);
  dff _59129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _23865_, clk);
  dff _59130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _24307_, clk);
  dff _59131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _01184_, clk);
  dff _59132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _25521_, clk);
  dff _59133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _26181_, clk);
  dff _59134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _06227_, clk);
  dff _59135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _18710_, clk);
  dff _59136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _06206_, clk);
  dff _59137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _09112_, clk);
  dff _59138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _06963_, clk);
  dff _59139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _11603_, clk);
  dff _59140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _03776_, clk);
  dff _59141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _28279_, clk);
  dff _59142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _23853_, clk);
  dff _59143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _24652_, clk);
  dff _59144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _06168_, clk);
  dff _59145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _25016_, clk);
  dff _59146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _26497_, clk);
  dff _59147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _04417_, clk);
  dff _59148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _10612_, clk);
  dff _59149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _04561_, clk);
  dff _59150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _04866_, clk);
  dff _59151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _03430_, clk);
  dff _59152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _04294_, clk);
  dff _59153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _04224_, clk);
  dff _59154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _02121_, clk);
  dff _59155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _02427_, clk);
  dff _59156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _03833_, clk);
  dff _59157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _03821_, clk);
  dff _59158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _03441_, clk);
  dff _59159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _04699_, clk);
  dff _59160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _26308_, clk);
  dff _59161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _08648_, clk);
  dff _59162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _08664_, clk);
  dff _59163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _28079_, clk);
  dff _59164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _23710_, clk);
  dff _59165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _23737_, clk);
  dff _59166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _04422_, clk);
  dff _59167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _16578_, clk);
  dff _59168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _01168_, clk);
  dff _59169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _06105_, clk);
  dff _59170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _11233_, clk);
  dff _59171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _03403_, clk);
  dff _59172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _27085_, clk);
  dff _59173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _11056_, clk);
  dff _59174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _04832_, clk);
  dff _59175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _04433_, clk);
  dff _59176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _03419_, clk);
  dff _59177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _04512_, clk);
  dff _59178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _04551_, clk);
  dff _59179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _03406_, clk);
  dff _59180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _04135_, clk);
  dff _59181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _04126_, clk);
  dff _59182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _04112_, clk);
  dff _59183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _06066_, clk);
  dff _59184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _04256_, clk);
  dff _59185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _04364_, clk);
  dff _59186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _06097_, clk);
  dff _59187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _06507_, clk);
  dff _59188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _06081_, clk);
  dff _59189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _04595_, clk);
  dff _59190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _09169_, clk);
  dff _59191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _04436_, clk);
  dff _59192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _04705_, clk);
  dff _59193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _08986_, clk);
  dff _59194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _09650_, clk);
  dff _59195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _09316_, clk);
  dff _59196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _06075_, clk);
  dff _59197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _10502_, clk);
  dff _59198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _10719_, clk);
  dff _59199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _13987_, clk);
  dff _59200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _06023_, clk);
  dff _59201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _11748_, clk);
  dff _59202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _12042_, clk);
  dff _59203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _11816_, clk);
  dff _59204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _06043_, clk);
  dff _59205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _12675_, clk);
  dff _59206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _12659_, clk);
  dff _59207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _05888_, clk);
  dff _59208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _23685_, clk);
  dff _59209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _05878_, clk);
  dff _59210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _04612_, clk);
  dff _59211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _21304_, clk);
  dff _59212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _22016_, clk);
  dff _59213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _21654_, clk);
  dff _59214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _22674_, clk);
  dff _59215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _15454_, clk);
  dff _59216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _15403_, clk);
  dff _59217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _04439_, clk);
  dff _59218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _13083_, clk);
  dff _59219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _13359_, clk);
  dff _59220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _13257_, clk);
  dff _59221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _06028_, clk);
  dff _59222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _13906_, clk);
  dff _59223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _03379_, clk);
  dff _59224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _04661_, clk);
  dff _59225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _04658_, clk);
  dff _59226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _04649_, clk);
  dff _59227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _03401_, clk);
  dff _59228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _04735_, clk);
  dff _59229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _04743_, clk);
  dff _59230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _02126_, clk);
  dff _59231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _16902_, clk);
  dff _59232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _16841_, clk);
  dff _59233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _16780_, clk);
  dff _59234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _16699_, clk);
  dff _59235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _04441_, clk);
  dff _59236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _14926_, clk);
  dff _59237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _06019_, clk);
  dff _59238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _15566_, clk);
  dff _59239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _18585_, clk);
  dff _59240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _18742_, clk);
  dff _59241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _18653_, clk);
  dff _59242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _05948_, clk);
  dff _59243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _19554_, clk);
  dff _59244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _05936_, clk);
  dff _59245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _17475_, clk);
  dff _59246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _17344_, clk);
  dff _59247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _18241_, clk);
  dff _59248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _18222_, clk);
  dff _59249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _18111_, clk);
  dff _59250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _05976_, clk);
  dff _59251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _04605_, clk);
  dff _59252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _15938_, clk);
  dff _59253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _16061_, clk);
  dff _59254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _15990_, clk);
  dff _59255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _05833_, clk);
  dff _59256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _23694_, clk);
  dff _59257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _23691_, clk);
  dff _59258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _23708_, clk);
  dff _59259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _23706_, clk);
  dff _59260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _23697_, clk);
  dff _59261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _04448_, clk);
  dff _59262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _23350_, clk);
  dff _59263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _23764_, clk);
  dff _59264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _23759_, clk);
  dff _59265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _23802_, clk);
  dff _59266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _23784_, clk);
  dff _59267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _23732_, clk);
  dff _59268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _23730_, clk);
  dff _59269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _05846_, clk);
  dff _59270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _23745_, clk);
  dff _59271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _05373_, clk);
  dff _59272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _04748_, clk);
  dff _59273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _05432_, clk);
  dff _59274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _03438_, clk);
  dff _59275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _05429_, clk);
  dff _59276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _00886_, clk);
  dff _59277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _03247_, clk);
  dff _59278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _03219_, clk);
  dff _59279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _04540_, clk);
  dff _59280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _00748_, clk);
  dff _59281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _05474_, clk);
  dff _59282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _04535_, clk);
  dff _59283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _00020_, clk);
  dff _59284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _05494_, clk);
  dff _59285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _05483_, clk);
  dff _59286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _04663_, clk);
  dff _59287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _03661_, clk);
  dff _59288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _05391_, clk);
  dff _59289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _05420_, clk);
  dff _59290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _03544_, clk);
  dff _59291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _04568_, clk);
  dff _59292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _03712_, clk);
  dff _59293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _03677_, clk);
  dff _59294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _03758_, clk);
  dff _59295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _23825_, clk);
  dff _59296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _23820_, clk);
  dff _59297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _05796_, clk);
  dff _59298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _24011_, clk);
  dff _59299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _23983_, clk);
  dff _59300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _23949_, clk);
  dff _59301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _04463_, clk);
  dff _59302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _03625_, clk);
  dff _59303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _25035_, clk);
  dff _59304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _24980_, clk);
  dff _59305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _04472_, clk);
  dff _59306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _24399_, clk);
  dff _59307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _24246_, clk);
  dff _59308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _24572_, clk);
  dff _59309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _24598_, clk);
  dff _59310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _24587_, clk);
  dff _59311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _25120_, clk);
  dff _59312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _25100_, clk);
  dff _59313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _25257_, clk);
  dff _59314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _25247_, clk);
  dff _59315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _05717_, clk);
  dff _59316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _24825_, clk);
  dff _59317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _24844_, clk);
  dff _59318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _24828_, clk);
  dff _59319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _25543_, clk);
  dff _59320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _25536_, clk);
  dff _59321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _25525_, clk);
  dff _59322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _05713_, clk);
  dff _59323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _25667_, clk);
  dff _59324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _25763_, clk);
  dff _59325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _05703_, clk);
  dff _59326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _04636_, clk);
  dff _59327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _27419_, clk);
  dff _59328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _27490_, clk);
  dff _59329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _05591_, clk);
  dff _59330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _04651_, clk);
  dff _59331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _27337_, clk);
  dff _59332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _05613_, clk);
  dff _59333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _05603_, clk);
  dff _59334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _26462_, clk);
  dff _59335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _05549_, clk);
  dff _59336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _27518_, clk);
  dff _59337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _27501_, clk);
  dff _59338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _27513_, clk);
  dff _59339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _27593_, clk);
  dff _59340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _27559_, clk);
  dff _59341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _05580_, clk);
  dff _59342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _27435_, clk);
  dff _59343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _07140_, clk);
  dff _59344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _04665_, clk);
  dff _59345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _28090_, clk);
  dff _59346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _00003_, clk);
  dff _59347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _28112_, clk);
  dff _59348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _04527_, clk);
  dff _59349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _28018_, clk);
  dff _59350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _28067_, clk);
  dff _59351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _04516_, clk);
  dff _59352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _27842_, clk);
  dff _59353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _27810_, clk);
  dff _59354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _27913_, clk);
  dff _59355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _27906_, clk);
  dff _59356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _05532_, clk);
  dff _59357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _27627_, clk);
  dff _59358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _27706_, clk);
  dff _59359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _05105_, clk);
  dff _59360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _02140_, clk);
  dff _59361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _02430_, clk);
  dff _59362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _04890_, clk);
  dff _59363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _04859_, clk);
  dff _59364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _04843_, clk);
  dff _59365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _04970_, clk);
  dff _59366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _04956_, clk);
  dff _59367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _07002_, clk);
  dff _59368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _05732_, clk);
  dff _59369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _07147_, clk);
  dff _59370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _07270_, clk);
  dff _59371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _05752_, clk);
  dff _59372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _05768_, clk);
  dff _59373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _06996_, clk);
  dff _59374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _05776_, clk);
  dff _59375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _05787_, clk);
  dff _59376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _06991_, clk);
  dff _59377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _07207_, clk);
  dff _59378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _05793_, clk);
  dff _59379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _05811_, clk);
  dff _59380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _06961_, clk);
  dff _59381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _05814_, clk);
  dff _59382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _05827_, clk);
  dff _59383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _05529_, clk);
  dff _59384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _05496_, clk);
  dff _59385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _02144_, clk);
  dff _59386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _04997_, clk);
  dff _59387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _05028_, clk);
  dff _59388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _05016_, clk);
  dff _59389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _05165_, clk);
  dff _59390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _05144_, clk);
  dff _59391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _05692_, clk);
  dff _59392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _07016_, clk);
  dff _59393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _05696_, clk);
  dff _59394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _07154_, clk);
  dff _59395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _05710_, clk);
  dff _59396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _07008_, clk);
  dff _59397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _05723_, clk);
  dff _59398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _07151_, clk);
  dff _59399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _07165_, clk);
  dff _59400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _05623_, clk);
  dff _59401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _05635_, clk);
  dff _59402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _07031_, clk);
  dff _59403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _07222_, clk);
  dff _59404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _05673_, clk);
  dff _59405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _07021_, clk);
  dff _59406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _05674_, clk);
  dff _59407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _05573_, clk);
  dff _59408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _07047_, clk);
  dff _59409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _05576_, clk);
  dff _59410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _05594_, clk);
  dff _59411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _07041_, clk);
  dff _59412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _07224_, clk);
  dff _59413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _05596_, clk);
  dff _59414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _05610_, clk);
  dff _59415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _05224_, clk);
  dff _59416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _07276_, clk);
  dff _59417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _05458_, clk);
  dff _59418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _05477_, clk);
  dff _59419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _07070_, clk);
  dff _59420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _05490_, clk);
  dff _59421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _07067_, clk);
  dff _59422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _05491_, clk);
  dff _59423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _05510_, clk);
  dff _59424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _07061_, clk);
  dff _59425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _05514_, clk);
  dff _59426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _07176_, clk);
  dff _59427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _05527_, clk);
  dff _59428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _05545_, clk);
  dff _59429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _07052_, clk);
  dff _59430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _05569_, clk);
  dff _59431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _07253_, clk);
  dff _59432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _05265_, clk);
  dff _59433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _07137_, clk);
  dff _59434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _05268_, clk);
  dff _59435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _28278_, clk);
  dff _59436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _05272_, clk);
  dff _59437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _05280_, clk);
  dff _59438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _07195_, clk);
  dff _59439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _07085_, clk);
  dff _59440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _07256_, clk);
  dff _59441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _05400_, clk);
  dff _59442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _05424_, clk);
  dff _59443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _07081_, clk);
  dff _59444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _05434_, clk);
  dff _59445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _07074_, clk);
  dff _59446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _05449_, clk);
  dff _59447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _05358_, clk);
  dff _59448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _07099_, clk);
  dff _59449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _07261_, clk);
  dff _59450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _05363_, clk);
  dff _59451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _05369_, clk);
  dff _59452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _07089_, clk);
  dff _59453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _05375_, clk);
  dff _59454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _07087_, clk);
  dff _59455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _01821_, clk);
  dff _59456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _08890_, clk);
  dff _59457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _08888_, clk);
  dff _59458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _01600_, clk);
  dff _59459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _08886_, clk);
  dff _59460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _05294_, clk);
  dff _59461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _05303_, clk);
  dff _59462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _07131_, clk);
  dff _59463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _05310_, clk);
  dff _59464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _05330_, clk);
  dff _59465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _07128_, clk);
  dff _59466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _28277_, clk);
  dff _59467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _05332_, clk);
  dff _59468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _05335_, clk);
  dff _59469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07120_, clk);
  dff _59470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _05353_, clk);
  dff _59471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _06073_, clk);
  dff _59472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _06046_, clk);
  dff _59473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _08145_, clk);
  dff _59474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _05163_, clk);
  dff _59475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _05154_, clk);
  dff _59476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _05869_, clk);
  dff _59477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _05866_, clk);
  dff _59478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _05843_, clk);
  dff _59479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _06120_, clk);
  dff _59480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _06112_, clk);
  dff _59481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _08143_, clk);
  dff _59482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _06211_, clk);
  dff _59483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _06165_, clk);
  dff _59484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _07295_, clk);
  dff _59485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _05940_, clk);
  dff _59486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _05930_, clk);
  dff _59487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _06529_, clk);
  dff _59488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _07297_, clk);
  dff _59489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _06286_, clk);
  dff _59490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _06267_, clk);
  dff _59491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _06403_, clk);
  dff _59492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _06401_, clk);
  dff _59493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _06389_, clk);
  dff _59494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _06134_, clk);
  dff _59495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _06841_, clk);
  dff _59496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _06927_, clk);
  dff _59497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _06908_, clk);
  dff _59498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _06903_, clk);
  dff _59499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _08074_, clk);
  dff _59500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _28275_, clk);
  dff _59501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06578_, clk);
  dff _59502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _06583_, clk);
  dff _59503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _06815_, clk);
  dff _59504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _06803_, clk);
  dff _59505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _06602_, clk);
  dff _59506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _28276_, clk);
  dff _59507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _06453_, clk);
  dff _59508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _06474_, clk);
  dff _59509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _06469_, clk);
  dff _59510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _06552_, clk);
  dff _59511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _06954_, clk);
  dff _59512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _06949_, clk);
  dff _59513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _07049_, clk);
  dff _59514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _07043_, clk);
  dff _59515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _07028_, clk);
  dff _59516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _08060_, clk);
  dff _59517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _06874_, clk);
  dff _59518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _06870_, clk);
  dff _59519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _28274_, clk);
  dff _59520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _07092_, clk);
  dff _59521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _07078_, clk);
  dff _59522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _07133_, clk);
  dff _59523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _07149_, clk);
  dff _59524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _07143_, clk);
  dff _59525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _07300_, clk);
  dff _59526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _07495_, clk);
  dff _59527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _07837_, clk);
  dff _59528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _28273_, clk);
  dff _59529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _07233_, clk);
  dff _59530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _07231_, clk);
  dff _59531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _07203_, clk);
  dff _59532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _07280_, clk);
  dff _59533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _07289_, clk);
  dff _59534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _07285_, clk);
  dff _59535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _07527_, clk);
  dff _59536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _07524_, clk);
  dff _59537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _07822_, clk);
  dff _59538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _07338_, clk);
  dff _59539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _07356_, clk);
  dff _59540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _07347_, clk);
  dff _59541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _07438_, clk);
  dff _59542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _07427_, clk);
  dff _59543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _07599_, clk);
  dff _59544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _07817_, clk);
  dff _59545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _07647_, clk);
  dff _59546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _07628_, clk);
  dff _59547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _07307_, clk);
  dff _59548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _07497_, clk);
  dff _59549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _07492_, clk);
  dff _59550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _07484_, clk);
  dff _59551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _10999_, clk);
  dff _59552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _10997_, clk);
  dff _59553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _07729_, clk);
  dff _59554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _28265_, clk);
  dff _59555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _10310_, clk);
  dff _59556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _10219_, clk);
  dff _59557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _07745_, clk);
  dff _59558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _10403_, clk);
  dff _59559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _10399_, clk);
  dff _59560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _07322_, clk);
  dff _59561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _28266_, clk);
  dff _59562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _09864_, clk);
  dff _59563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _09838_, clk);
  dff _59564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _09791_, clk);
  dff _59565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _10116_, clk);
  dff _59566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _28267_, clk);
  dff _59567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _11179_, clk);
  dff _59568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _28264_, clk);
  dff _59569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _07723_, clk);
  dff _59570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _07436_, clk);
  dff _59571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _10709_, clk);
  dff _59572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _10802_, clk);
  dff _59573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _10779_, clk);
  dff _59574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _07731_, clk);
  dff _59575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _07720_, clk);
  dff _59576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _11282_, clk);
  dff _59577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _11310_, clk);
  dff _59578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _11305_, clk);
  dff _59579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _07715_, clk);
  dff _59580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _11034_, clk);
  dff _59581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _28263_, clk);
  dff _59582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _11151_, clk);
  dff _59583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _11348_, clk);
  dff _59584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _11544_, clk);
  dff _59585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _28261_, clk);
  dff _59586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _11538_, clk);
  dff _59587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _28262_, clk);
  dff _59588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _11249_, clk);
  dff _59589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _11247_, clk);
  dff _59590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _11228_, clk);
  dff _59591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _12075_, clk);
  dff _59592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _12071_, clk);
  dff _59593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _11825_, clk);
  dff _59594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _11814_, clk);
  dff _59595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _11810_, clk);
  dff _59596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _07703_, clk);
  dff _59597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _11878_, clk);
  dff _59598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _11965_, clk);
  dff _59599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _07329_, clk);
  dff _59600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _11587_, clk);
  dff _59601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _11593_, clk);
  dff _59602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _28258_, clk);
  dff _59603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _07707_, clk);
  dff _59604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _28259_, clk);
  dff _59605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _28260_, clk);
  dff _59606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _11415_, clk);
  dff _59607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _05918_, clk);
  dff _59608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _05957_, clk);
  dff _59609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _05938_, clk);
  dff _59610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _02148_, clk);
  dff _59611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _05366_, clk);
  dff _59612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _05321_, clk);
  dff _59613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _05289_, clk);
  dff _59614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _05598_, clk);
  dff _59615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _12119_, clk);
  dff _59616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _07695_, clk);
  dff _59617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _03386_, clk);
  dff _59618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _07694_, clk);
  dff _59619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _07442_, clk);
  dff _59620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _28257_, clk);
  dff _59621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _12033_, clk);
  dff _59622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _12026_, clk);
  dff _59623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _28254_, clk);
  dff _59624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _07446_, clk);
  dff _59625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _10203_, clk);
  dff _59626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _28255_, clk);
  dff _59627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _08830_, clk);
  dff _59628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _28256_, clk);
  dff _59629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _25090_, clk);
  dff _59630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _07335_, clk);
  dff _59631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _07623_, clk);
  dff _59632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _28243_, clk);
  dff _59633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _08930_, clk);
  dff _59634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _07640_, clk);
  dff _59635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _09621_, clk);
  dff _59636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _07353_, clk);
  dff _59637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _03071_, clk);
  dff _59638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _03696_, clk);
  dff _59639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _01220_, clk);
  dff _59640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _23756_, clk);
  dff _59641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _07407_, clk);
  dff _59642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _23714_, clk);
  dff _59643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _27374_, clk);
  dff _59644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _07673_, clk);
  dff _59645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _03636_, clk);
  dff _59646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _03121_, clk);
  dff _59647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _11280_, clk);
  dff _59648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _07569_, clk);
  dff _59649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _28251_, clk);
  dff _59650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _11045_, clk);
  dff _59651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _11005_, clk);
  dff _59652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _28252_, clk);
  dff _59653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _12126_, clk);
  dff _59654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _12115_, clk);
  dff _59655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _11728_, clk);
  dff _59656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _07545_, clk);
  dff _59657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _11812_, clk);
  dff _59658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _07543_, clk);
  dff _59659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _11602_, clk);
  dff _59660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _11650_, clk);
  dff _59661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _28250_, clk);
  dff _59662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _07489_, clk);
  dff _59663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _28244_, clk);
  dff _59664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _06646_, clk);
  dff _59665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _06727_, clk);
  dff _59666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _07642_, clk);
  dff _59667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _07455_, clk);
  dff _59668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _11635_, clk);
  dff _59669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _11883_, clk);
  dff _59670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _28245_, clk);
  dff _59671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _27630_, clk);
  dff _59672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _28247_, clk);
  dff _59673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _08734_, clk);
  dff _59674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _28248_, clk);
  dff _59675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _07667_, clk);
  dff _59676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _09529_, clk);
  dff _59677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _09346_, clk);
  dff _59678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _28249_, clk);
  dff _59679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _09728_, clk);
  dff _59680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _07579_, clk);
  dff _59681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _07390_, clk);
  dff _59682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _07429_, clk);
  dff _59683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _07588_, clk);
  dff _59684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _07586_, clk);
  dff _59685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _28240_, clk);
  dff _59686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _05807_, clk);
  dff _59687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _06987_, clk);
  dff _59688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _07592_, clk);
  dff _59689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _04507_, clk);
  dff _59690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _07594_, clk);
  dff _59691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _04946_, clk);
  dff _59692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _28241_, clk);
  dff _59693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _02284_, clk);
  dff _59694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _02256_, clk);
  dff _59695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _01148_, clk);
  dff _59696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _09707_, clk);
  dff _59697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _27110_, clk);
  dff _59698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _10949_, clk);
  dff _59699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _09108_, clk);
  dff _59700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _28373_, clk);
  dff _59701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _25875_, clk);
  dff _59702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _08971_, clk);
  dff _59703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _07401_, clk);
  dff _59704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _09817_, clk);
  dff _59705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _03339_, clk);
  dff _59706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _09725_, clk);
  dff _59707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _03241_, clk);
  dff _59708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _09849_, clk);
  dff _59709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _08392_, clk);
  dff _59710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _28372_, clk);
  dff _59711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _06674_, clk);
  dff _59712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _06676_, clk);
  dff _59713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _06696_, clk);
  dff _59714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _06670_, clk);
  dff _59715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _09502_, clk);
  dff _59716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _11433_, clk);
  dff _59717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _06736_, clk);
  dff _59718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _07173_, clk);
  dff _59719_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _59720_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _59721_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _59722_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _59723_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _59724_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _59725_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _59726_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _59727_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _59728_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _59729_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _59730_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _59731_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _59732_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _59733_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _59734_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _59735_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _59736_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _59737_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _59738_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _59739_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _59740_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _59741_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _59742_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _59743_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _59744_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _59745_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _59746_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _59747_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _59748_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _59749_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _59750_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _59751_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _28377_, clk);
  dff _59752_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _28378_[0], clk);
  dff _59753_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _28378_[1], clk);
  dff _59754_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _28378_[2], clk);
  dff _59755_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _28378_[3], clk);
  dff _59756_ (\oc8051_top_1.oc8051_sfr1.bit_out , _28379_, clk);
  dff _59757_ (\oc8051_top_1.oc8051_sfr1.wait_data , _28380_, clk);
  dff _59758_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _28381_[0], clk);
  dff _59759_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _28381_[1], clk);
  dff _59760_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _28381_[2], clk);
  dff _59761_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _28381_[3], clk);
  dff _59762_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _28381_[4], clk);
  dff _59763_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _28381_[5], clk);
  dff _59764_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _28381_[6], clk);
  dff _59765_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _28381_[7], clk);
  dff _59766_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10496_, clk);
  dff _59767_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10525_, clk);
  dff _59768_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10523_, clk);
  dff _59769_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10419_, clk);
  dff _59770_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10656_, clk);
  dff _59771_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10640_, clk);
  dff _59772_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10463_, clk);
  dff _59773_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10236_, clk);
  dff _59774_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _07405_, clk);
  dff _59775_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _07403_, clk);
  dff _59776_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _07413_, clk);
  dff _59777_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _07411_, clk);
  dff _59778_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _07410_, clk);
  dff _59779_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _07416_, clk);
  dff _59780_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _07419_, clk);
  dff _59781_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06574_, clk);
  dff _59782_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _09965_, clk);
  dff _59783_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _10109_, clk);
  dff _59784_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _10106_, clk);
  dff _59785_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _10072_, clk);
  dff _59786_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _10048_, clk);
  dff _59787_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _09911_, clk);
  dff _59788_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _10146_, clk);
  dff _59789_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _09770_, clk);
  dff _59790_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09935_, clk);
  dff _59791_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _10099_, clk);
  dff _59792_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _10010_, clk);
  dff _59793_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _09967_, clk);
  dff _59794_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _10103_, clk);
  dff _59795_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _10101_, clk);
  dff _59796_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _10007_, clk);
  dff _59797_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _09814_, clk);
  dff _59798_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _06634_, clk);
  dff _59799_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _06561_, clk);
  dff _59800_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _16327_, clk);
  dff _59801_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _16306_, clk);
  dff _59802_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _16265_, clk);
  dff _59803_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _23805_, clk);
  dff _59804_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _23794_, clk);
  dff _59805_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _15545_, clk);
  dff _59806_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _15524_, clk);
  dff _59807_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _06819_, clk);
  dff _59808_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _15857_, clk);
  dff _59809_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _17867_, clk);
  dff _59810_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _06627_, clk);
  dff _59811_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _14987_, clk);
  dff _59812_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _15098_, clk);
  dff _59813_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _06631_, clk);
  dff _59814_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _15382_, clk);
  dff _59815_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _15361_, clk);
  dff _59816_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _06487_, clk);
  dff _59817_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _23806_, clk);
  dff _59818_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _14554_, clk);
  dff _59819_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _23789_, clk);
  dff _59820_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _27260_, clk);
  dff _59821_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _24915_, clk);
  dff _59822_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _25019_, clk);
  dff _59823_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _14744_, clk);
  dff _59824_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _23807_, clk);
  dff _59825_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _23792_, clk);
  dff _59826_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _01698_, clk);
  dff _59827_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _14262_, clk);
  dff _59828_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _14241_, clk);
  dff _59829_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _14220_, clk);
  dff _59830_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _14199_, clk);
  dff _59831_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _23808_, clk);
  dff _59832_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _23791_, clk);
  dff _59833_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _23798_, clk);
  dff _59834_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _01703_, clk);
  dff _59835_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _13695_, clk);
  dff _59836_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _13674_, clk);
  dff _59837_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _13653_, clk);
  dff _59838_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _13611_, clk);
  dff _59839_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _13590_, clk);
  dff _59840_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _23809_, clk);
  dff _59841_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _23790_, clk);
  dff _59842_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _00821_, clk);
  dff _59843_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _23773_, clk);
  dff _59844_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _07608_, clk);
  dff _59845_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _23782_, clk);
  dff _59846_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _23777_, clk);
  dff _59847_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _23781_, clk);
  dff _59848_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _23780_, clk);
  dff _59849_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _23779_, clk);
  dff _59850_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _10960_, clk);
  dff _59851_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _23762_, clk);
  dff _59852_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _23761_, clk);
  dff _59853_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _07621_, clk);
  dff _59854_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _23768_, clk);
  dff _59855_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _23765_, clk);
  dff _59856_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _23767_, clk);
  dff _59857_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _23766_, clk);
  dff _59858_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _10878_, clk);
  dff _59859_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _23750_, clk);
  dff _59860_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _23749_, clk);
  dff _59861_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _23748_, clk);
  dff _59862_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _23747_, clk);
  dff _59863_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _07631_, clk);
  dff _59864_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _23754_, clk);
  dff _59865_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _23757_, clk);
  dff _59866_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _11084_, clk);
  dff _59867_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _23736_, clk);
  dff _59868_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _23735_, clk);
  dff _59869_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _07671_, clk);
  dff _59870_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _23743_, clk);
  dff _59871_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _23739_, clk);
  dff _59872_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _23742_, clk);
  dff _59873_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _23741_, clk);
  dff _59874_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _11060_, clk);
  dff _59875_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10321_, clk);
  dff _59876_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10304_, clk);
  dff _59877_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10295_, clk);
  dff _59878_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10307_, clk);
  dff _59879_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10323_, clk);
  dff _59880_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10231_, clk);
  dff _59881_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _10002_, clk);
  dff _59882_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _07583_, clk);
  dff _59883_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _09777_, clk);
  dff _59884_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _09774_, clk);
  dff _59885_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _09702_, clk);
  dff _59886_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _09889_, clk);
  dff _59887_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _09876_, clk);
  dff _59888_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _09732_, clk);
  dff _59889_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _09861_, clk);
  dff _59890_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _07590_, clk);
  dff _59891_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _05147_, clk);
  dff _59892_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _04677_, clk);
  dff _59893_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _11019_, clk);
  dff _59894_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _10891_, clk);
  dff _59895_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _06762_, clk);
  dff _59896_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _11598_, clk);
  dff _59897_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _11226_, clk);
  dff _59898_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _11295_, clk);
  dff _59899_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _11285_, clk);
  dff _59900_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _01847_, clk);
  dff _59901_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _09714_, clk);
  dff _59902_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _07482_, clk);
  dff _59903_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _08950_, clk);
  dff _59904_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _08904_, clk);
  dff _59905_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _08169_, clk);
  dff _59906_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _08057_, clk);
  dff _59907_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _07735_, clk);
  dff _59908_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _10027_, clk);
  dff _59909_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _08140_, clk);
  dff _59910_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _10145_, clk);
  dff _59911_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _04825_, clk);
  dff _59912_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _04619_, clk);
  dff _59913_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _04481_, clk);
  dff _59914_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _06782_, clk);
  dff _59915_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _01270_, clk);
  dff _59916_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _01356_, clk);
  dff _59917_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _08542_, clk);
  dff _59918_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _10279_, clk);
  dff _59919_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _23738_, clk);
  dff _59920_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _06791_, clk);
  dff _59921_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _01268_, clk);
  dff _59922_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _03700_, clk);
  dff _59923_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _02759_, clk);
  dff _59924_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _01495_, clk);
  dff _59925_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _25539_, clk);
  dff _59926_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _04365_, clk);
  dff _59927_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _01872_, clk);
  dff _59928_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _01353_, clk);
  dff _59929_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _03730_, clk);
  dff _59930_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _03590_, clk);
  dff _59931_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _03580_, clk);
  dff _59932_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _01412_, clk);
  dff _59933_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _27718_, clk);
  dff _59934_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _06806_, clk);
  dff _59935_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _08328_, clk);
  dff _59936_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _05204_, clk);
  dff _59937_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _05182_, clk);
  dff _59938_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _06839_, clk);
  dff _59939_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _06792_, clk);
  dff _59940_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _11622_, clk);
  dff _59941_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _11626_, clk);
  dff _59942_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _11624_, clk);
  dff _59943_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _24948_, clk);
  dff _59944_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _11632_, clk);
  dff _59945_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _11630_, clk);
  dff _59946_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _06661_, clk);
  dff _59947_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _06973_, clk);
  dff _59948_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _11351_, clk);
  dff _59949_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _11343_, clk);
  dff _59950_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _11346_, clk);
  dff _59951_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _11214_, clk);
  dff _59952_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _11138_, clk);
  dff _59953_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _11185_, clk);
  dff _59954_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _11068_, clk);
  dff _59955_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _06946_, clk);
  dff _59956_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _06921_, clk);
  dff _59957_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _05262_, clk);
  dff _59958_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _05251_, clk);
  dff _59959_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _05254_, clk);
  dff _59960_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _10713_, clk);
  dff _59961_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _10701_, clk);
  dff _59962_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _10705_, clk);
  dff _59963_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _10676_, clk);
  dff _59964_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _07103_, clk);
  dff _59965_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _10488_, clk);
  dff _59966_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _10347_, clk);
  dff _59967_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _10379_, clk);
  dff _59968_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _10172_, clk);
  dff _59969_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _10134_, clk);
  dff _59970_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _10132_, clk);
  dff _59971_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _10130_, clk);
  dff _59972_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _06567_, clk);
  dff _59973_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _06708_, clk);
  dff _59974_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _09641_, clk);
  dff _59975_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _23686_, clk);
  dff _59976_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _09646_, clk);
  dff _59977_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _09643_, clk);
  dff _59978_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _12253_, clk);
  dff _59979_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _09651_, clk);
  dff _59980_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _09648_, clk);
  dff _59981_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _06684_, clk);
  dff _59982_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _23731_, clk);
  dff _59983_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _23729_, clk);
  dff _59984_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _23728_, clk);
  dff _59985_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _23727_, clk);
  dff _59986_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _23726_, clk);
  dff _59987_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _23722_, clk);
  dff _59988_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _23862_, clk);
  dff _59989_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _23858_, clk);
  dff _59990_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _23851_, clk);
  dff _59991_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _23723_, clk);
  dff _59992_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _23861_, clk);
  dff _59993_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _06514_, clk);
  dff _59994_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _06502_, clk);
  dff _59995_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _03909_, clk);
  dff _59996_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _04300_, clk);
  dff _59997_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _27655_, clk);
  dff _59998_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _27668_, clk);
  dff _59999_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _23856_, clk);
  dff _60000_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _27665_, clk);
  dff _60001_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _23852_, clk);
  dff _60002_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _23724_, clk);
  dff _60003_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _23859_, clk);
  dff _60004_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _27661_, clk);
  dff _60005_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _23725_, clk);
  dff _60006_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _23850_, clk);
  dff _60007_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _23721_, clk);
  dff _60008_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _23720_, clk);
  dff _60009_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _23719_, clk);
  dff _60010_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _23718_, clk);
  dff _60011_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _23717_, clk);
  dff _60012_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _27658_, clk);
  dff _60013_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _27690_, clk);
  dff _60014_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _27702_, clk);
  dff _60015_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _27697_, clk);
  dff _60016_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _27693_, clk);
  dff _60017_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _23712_, clk);
  dff _60018_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _23711_, clk);
  dff _60019_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _23709_, clk);
  dff _60020_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _06512_, clk);
  dff _60021_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _23705_, clk);
  dff _60022_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _23704_, clk);
  dff _60023_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _23703_, clk);
  dff _60024_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _23702_, clk);
  dff _60025_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _23701_, clk);
  dff _60026_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _23698_, clk);
  dff _60027_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _23844_, clk);
  dff _60028_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _23837_, clk);
  dff _60029_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _23847_, clk);
  dff _60030_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _23836_, clk);
  dff _60031_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _03899_, clk);
  dff _60032_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _23843_, clk);
  dff _60033_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _23839_, clk);
  dff _60034_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _23846_, clk);
  dff _60035_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _23838_, clk);
  dff _60036_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _23842_, clk);
  dff _60037_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _23840_, clk);
  dff _60038_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _23845_, clk);
  dff _60039_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _27623_, clk);
  dff _60040_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _23841_, clk);
  dff _60041_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _23699_, clk);
  dff _60042_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _23835_, clk);
  dff _60043_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _23700_, clk);
  dff _60044_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _23834_, clk);
  dff _60045_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _23788_, clk);
  dff _60046_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _23787_, clk);
  dff _60047_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _27621_, clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
